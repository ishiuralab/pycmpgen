module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [12:0] src14;
    reg [11:0] src15;
    reg [10:0] src16;
    reg [9:0] src17;
    reg [8:0] src18;
    reg [7:0] src19;
    reg [6:0] src20;
    reg [5:0] src21;
    reg [4:0] src22;
    reg [3:0] src23;
    reg [2:0] src24;
    reg [1:0] src25;
    reg [0:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3])<<23) + ((src24[0] + src24[1] + src24[2])<<24) + ((src25[0] + src25[1])<<25) + ((src26[0])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2024af672fcab06c2bda2fd528a57ddb5beddc38bfabc3c82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a710456c16f0ab43834a34f113238d81f5dc60665427129b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b905e94f26644cd6040593697e61c96fa0e066729f8d6c79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8a916c092d0095bae8ed0577f00b438f171b72320ad1c8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfea2cc5f5188fcba2c231dc6b6b815212a94c198eea0414c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ffb278156543615e6a30105140a711b842746238ad0df510;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a085b7cf174d49db0a19d9128517bcfe916bb563bc848103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d27e1d73ee937e64f4a6946b411f6586bd9a11110370cf06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb60b004325d38a9cdd2b9240442cb911aeabc2a5480678af0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc5e2d7e26fa6dd34f57a53d225b692b728d45ed99e197c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19557352d3808220ab1ab147a75f5548df148410747bb8877;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d92dff0d289452f40af47c91e98e0d46e25da881eab00fce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he12cbd5c1255503b932839534503a03f4d08b3af8931c860;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fb47fbf9bc255b421b0687c89e9ddf0bc866935f02cf2e1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h648f0e6af155df479eab2892b40e12a30d96b3840fe05ee7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c155dba0b87b57a4c536dee63892e9337890b50e912191a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8abf918fb5faed83413c9d11ea53fd311f4dcf24bc37f4f7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9753bf012014bab1b97bd7fdcabd84e3c3fc7adfb65efa234;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8322389a53ad5aef7938786ed51fd8855fc1efa6b5e50f043;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0af7f08aab65097b98751ad9b2455b030c477a8f8c1c3aea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5dd747f97c4d2ac4f09dcf27bd4445419acd07df4a6d0379;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9445c004416cfac803bde03b9fddd121dc4fe39309cbc0bc0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7f66aae139c639b6ec8be1f6a6488e7008a8b67b1cab5ada;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc1a274d4ff04f901b857a251bd53500c4373ee1d63507c7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64538a809e83dd6803fec9b486b4919ef1e575f0d9e8c1a9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19a1116a293fed9713104457fdd38780787fcbebd01285d26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a020f2ad4962278b37e7418df34f655213b40753ad82372e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1048c77802da32cdc5ea4c8e04691854f964822748477ac90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8dd08e50baee8d2b8382ce5bd4f85f2514ca077e0787f77d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h436faca4e2dd3bdd6d9fec8ffcebb86715b18360a64108b3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20d37b13b71cc4e7d334fc80f2886d0de5c14972cb145ca2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbd14eaf97994cb24414ddf875e911f23df2c66cf5fbdd2a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf544c56ebbca1aad062e823172d1a1fc96e77c51e948be741;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha80bcbe404e40a452eb0af9746291651ab6aa2738d1d01bb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f4f3e00c0261acea2682422086ed12b351e14715af940150;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88522a37918051a0a1a85b6864dfa44c9c5ed6b3c501f2cd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13f062e98a26752abe1b09bcafc370d19693c17b8efc5b81c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e6e8ae4f12ec1bd4b0db01d3252cbf2c9171866d421c3b10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12cfa2ff217ec93182dc67e582ca1358b5e6126403165e73a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70cfeed044be41a2a597f03495f00b44fc496b045c5c5752d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9b20e6cb8b64100b3ef4b92e1fa3befaa32cd993b80c55de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab28224626736ac77e75a3e25d86ce570c1be2a44a98f9ac2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bc70de43d77adc588a5b1af551c640a0e6db1249d48ea6ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5227eb6d879f0f90af0a60dbf7baf9cc0f1677cdc122c4a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h685db21c369eb4d48ae3c93545e2c38df452af4a60440395f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3baeb8bf9246e34b560ed3b22f7b78315f46e1fb0e1335507;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc49aca98bca2dfc87866c327b9a9f632b1bcf2d361d88f71a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h436d544a8b307c6ac9d0f0a224803cae8e7bd479f303f2730;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h636b7e17f207d8f20ef7ecdaefa59db5d0a07e8e71599bbb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb286ceca566d608fbf82f68b225b62efd8087a1cf1c34e6b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0d5ed55a739a53b68e753e1ce5b0cf4c9aa89ee39652ebac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d4eafbf4e0c2ada4ff77c1f4c549a3078dc5c4ca70ba0bb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h116ed1e76780978043728da604f6163333017e3312a37a752;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2b16c530afa4aa1c6794e3e139aa7265f16ad6adf2774d60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f128c4d6749e89cf32b0c669daa11534b043af21feff2739;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0b113c0b045ee1807c6f2a2dfe21c99f3a3c91878264bb9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c699d827ebf1ad3b79e7d0c1afe584bdd952b02143b8e9a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2266ae8ba2fed7310536808250c6f08995dfc66c0dd9dd70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf17867a66a2d288305d85b695bc131d984ee8e3818c49aede;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fc4bb3b95be0f8b6a75ee4ed0189611975a6917e8c3f13c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ddc61bbf4b5e97c1698c3d941d6366d677ab4f88d6a2fca9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5eaca0858f75122b4dbc0c9d02434d4133f1817a05d85dc22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe517bf1c1e5ab33964423102a7b421c8a05379748bd5f34a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h430279f8ebc60a6883e8d717b3b8c9b7ef27b40346c8fb29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57e817052ba0f2b1b0bfd03291040902ed2a785a5f4f2027;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21a14f60718b37ec013fddbd023c9f650e0232c9b2c44a4bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2867d54a32a1d962e0828e1c781c3af174061f3d8d08e82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9df8e806b8c0ead4e390d19bd692d026554fd31b8fbc3e53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d61c7ba6469bcaadcdf75683b809deac3c2f1d241767932;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b6159105d83e3463a58fa7ee7a1c43de98880af1c281ddb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14a2a84417a4d041d4b5048579c668b777b02a2e62a15bb84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f850660ef66fc0382d7292d156c194736448cf0af24a62fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41f64d81925d8464ab8b902b8372a9bc077b7a950037a12cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bc60f18c21b354aa334ab880039ba35acf83f06858c91c88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55392bb550a45bda14ca613f44aec6b7172f90466daaea6f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16bb1c3879fd757c30ded7234b87823a4eaea2005fff91368;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e786ae1768c60feb0b799aad620194a1f48b32b5228bbe50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8505c4830f87e77d3f833de3eceaba330e5a961b7e4d646cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8918fe264b0125066633a6d7cd36849e6c537f8aa66071a79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbfefdd43c481dce018efabe609d8c28e8d5fa65f2d2da154;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a1dcb8731ebe3d2dfaa2f6a45d231016e7974f011384363c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d33d626befe0d6d329318f352fa0e5843a426c498222f67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8867c1e3f63844585d6d955ef9de16cbcb8c9c6d7febec9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h909f619c222f0c4485ae7062f259251d9ac86443d024b4082;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h380e988b5e0aec83629c21dfb9b3aa0e045c5b188d51e216b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3552f40736cb87561a8a8c7f2d2c99b13f706d46fd7f82146;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c5957d4b0205bae7e09dba68d8b0fe281ddef45a5381e99f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd31888096435c716e80e046e46b0d04a61fb0c7ff64e88065;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0e243392f2603ecc23453e1a1eea05a9c7c1bf8ba82552e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc50f34844c745f0d4e12fb517dd893afd35faa2957ddb273;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34c2bf8366034f55ab26efc603a3501e9979821930c02a468;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3f2183785e0bd2e4d069bc1f00e0b3e903660821264f42a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0774fee537e9bfd9b9a5fffd3907c27e8a13d10be64d1f2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc06af5442005428fa8136913f1db9a0d26a196b8824a94eb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff35a7c6fc9940bf677230983255660afd5c33a98805fbf88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c632c5adc2ec7036b7bae91d4985fdfdee1fcd84695262d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ed14031906666d5429851e13a988b4b72923ce7834f16358;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb7e5e250e632cdd8e9bcac7c374a06b4a2b65db6b6590dc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff38f44e72c89709c64574c17800727a5c12ed65b732bfe53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h223192bbc07cb3d552aa4324816928a516ea7bc177fd01093;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc4455cf438ef1cfce63e2c68e536f24ea508f342156463ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11f0f11e6d22aeae8bf7237c9803d5cffc4a1e1f353fceaf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h176393f0e79a8472ced4688caf58083394d87d78a2f3190cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd2997f0ccd2aefad1f07f8a330588f0b13d7c68b1a32c5c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55127551838ad3202e1dc8a561a3b29ef76f5ea04feba95b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdf5c891acbf6b443403e1ca62e490693fd9a4e7101dd519a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2d294eacb4a1036b026e62d9196629d509e67b47153bde01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43cbfd19aa594159d6a66b46ceacb520b8422e8f03d882c8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fe5b5cbcb988ad26c0bb3ee1bc9a2ffd254651f18779137d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb11c0ccbd8b8832974b9fea969841473845ae2e14c7eeed4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7738305367b1664b28bc4b46b3add36caf6dda438bde0097;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcc6dff1e881516554e7fe05aad88faa0cadfe17ef3fbd62e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1221555e31074166a21cc1a93f1e5e38435ba74c740559c05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24bcebf05af35972835a735c238760b9e2e04933c34a5d5fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h169f13f00f832840c5ef341050af85ae7e17f522a707640bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fba1a019b6c16f09bf8eee7139044232a3376d5d9c176348;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79f1d98e72b811960742b44fe2346b21c09dc2996b7e44ccf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h690ca82816566a507fe23e8275c354ab5ae407ff3a6f7f625;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40e6a449ef28f25c51d729cd40f6097385d202660d5c49552;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6afaacec5c152e260ea7a08e326140c3b860e6eef1ecde582;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2060da73ac1f3942f15630a6de4eb31dacb052b47f715d21f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dc482ccec5a5c0c4aa96c917238d189c91d06a486ae302fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42060bf6dc2c837ec5543900f82cf89ba26cb9da491dcf3c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9514c08d020e9da4fb99273bfb8cd8b6f3c7a04560c41c16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heecce8bbcd2dcd26a24ed49943801578d6382f2a01b7bfcf4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcdd3c2e38e1bacaa53d94e529259fff6e07034fe4bd8875f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c21ebed252962f2235912cd06508111ff78e33ec9e7bf8f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8012c1cfeb7f2a209e98b3db237d97d95c42906c4e7bebe58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38839e446399b2e57d4155cc5751d4fe2db4bb69717238547;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc953207e9f474d12cbb66fae7efd7d451b9387866009d3cf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7f05cf1ea946340c995d7d2b1773d057a88d2088cf9dd15f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33d1bfbf299edcef1a2445cbb3d7993f51b2af72f9606134d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13a09fb4192715505df08bc4b2b378573ed5dfe3b83e29ff7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ebe07f7f927040ae8573fc9cd2484c8a28929d5fe7147cff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc066de27e2d61867d16cb1d6d0c8ce640ed0a1e187845b13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc65cf67b7a70bcf7b0998e6399da8556a2d41ddd48013d544;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he67bc5d225ede5067bb77a0706e574e5723338cb944b16b30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4888fa68fabb70958825ac4077f391e95ea1c9dfdecd7ccd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fee3fce435fc614b74eab11ca09b38549ce2a637010416d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h760fadce020b69f502ea07deb53bad6eea30ed92ce40cc31a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5fbe99749272f7f2f26c653b164aa394cf7b317eb28cb6f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8368fbe7670764d6e5eebdd9b5e18339cd38f0f07517edc8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h157a312a6be7d749da6bbe85d85dd3445ca4345c2db381e4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e35fb1e16212a20aed60d343f1f95e021ef2b7661d1b2e6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b72d53b5886a80d32e8c0224ccd1102afd1b5f5a4ac8d949;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h380780c3c9c39513cca5251f692a5de24eb0f8ea5d7b06e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h603a65f4e1172757783258528dd399b45af6eb0c8d2a10d36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h692266a965b2fb4d34ab99bc8aa0e2c56a5d7fec39e4c951e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a37cf859e63a75afcc2efd32b3c8641fb290029586f64bcc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h407bd3e2909327de96ef4fc84d0dc7018cc0aaca0a7c16a40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f8ecea410e0105780f2f0af2c8dad0fc15050c2f8c73d90b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd29e99e679ca88b67d6961f75e3406b36fbf70d9386f84e93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f1fea4b5d0e0f2d336c48654114a62426a5704ac11238bae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadbe3d27d6f441a69ed1f086e2af8aa013ad524ebadb95cb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0284fabbe0d4f53efc5bfe1e9d757647b97920eaaf38fac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76535f8d80e55269706b3d8746e9d7c5fa2d19a2739b3dc95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78d6475a3b52f7400e5a475f1d5e885df059331d4065f54a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h293b5592832f33a8c19e7665057135ade771fafcb2d97ae75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b0592a55810e4ded2dc24fc883195fb2d1efeb43e29a7df4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h923f95cc84386057c526cc9c0e51ac2ebb2437cb9567d1d10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97abf116ac367cfc2d96a6c8ec471aa86c12b56b8a40405c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87a85b1855009330d9521b6f48b97c30a0479cbca7b1970e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79f88c95216eea55db032987bf5f8e321cce4a6549103dea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a0c062f3befb4572f19917e8764f77bc05345efb7965f784;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5110d2e1923a014373afdf15b3e12f6179046424cc5b0d0ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0fe7f01da111b79cb57d9662f80b2feaae9348ea74322d76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a7f789e8b21b122c1817aba27e144e23c7bea5d68d7081a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3854f69143e5f7bf21de103ffedf9d55def521698b8b41c37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbecd9a6f04f7c956a5430b265a1eb57dc5e1ebc0a45520e6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e47b68c3a37bfeb95ce7e6ba314498bc94e6f5d3186e041;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h891bbc873309d6785a1b4e54b39f9cb0f9706e3d99c349ac8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1c358b5df9218861a8baab9cad4ce87460a9948de8a3cd9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b12acff5fec8e08ab3ac96b2b61c35c07bd53ba25736d28a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h133b24036f23dfe3ce781face0963594298422afa10db19be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h968add3127fbe5c6d587d314030b7ad225432613f92c70259;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h714100bef421c96a4376c199d68c03955a73ed0521c3d5e06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdad3398f3f73bdcf98c64815e3438670428c2f1511de601c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h820024ee719f58510bddf7774819c98829bfd56a79e47a3e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbaa7b018c7fc8cb5e6cb38142b48b5ac565eab18dfd2d3b9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h855c77e06d80c71a4c012d6b1804a424640505e24e60c24a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0fccaf2a7db58182cdf2ceeef64b1f1740449a37f6cb6e5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9313ac830274f50f62fbee49dec66d36dfeffd603e23a1b57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49cac79d1ade8a2b46303e99310bb7a9477c885b9cdfcc4a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb78beced5608505d117e729bbcaa98df7e32a14e5993ee4cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe0ca8b9045a702a229b6ca37e3ef41a8144cd41c66c4e406;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2412a39ad9f8d98f64fb9f65e2affcf5ddac7255dcf13e114;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3275338294e29aa07bb46d1686ccbcab3de0b6f4e46c4aa24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b7e849ea492f02cdf8d58319bec44ae1a398043331c2f6a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h800e09888ce93e278d061c5fce1b87f9c37172743c3ffb7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a45bccfaf0ef000684227be3a802881b13b7e9f952bd68de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa99d1ea136b82a78cdbc424345a49b7872a875f524406085;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8c61e0cd97eedb913b0ee61e7d06158a512e3e2deb8f6f73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84e91fe3a2b26dc7a45e86e3fb0f1ad033dc54b5f7d782e69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecbbad38845533b32be8fa3165122b58a01cf29c9e1d0738f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5613995bdedffe07bb468bf8c11e136d4a84d960696071726;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47ea5d657c869a34e3de7e11f1c67275969b513db7d702702;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e766ab109ccef6587d2a7c2f814b39ab476f0622562d7e36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30c84ea0cf64e244e49b4e783c06f03785b6e2292fc1dd035;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h532e1e1c67d73292f2e166d0ce1f0923bf1779ff3aad7259;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51ff17008f5444f355d553e72293f049df6cb129e4b8687bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe0efde666f8be90bdcc317a7bc6d80dc7ffaae57627c2495;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29edd70f09f7f2b769a78cd9b26a50a62d4da5ae5a9814d05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac8b23d32bb318b9f789bf3934a67947215513e9939bb4e38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddce5c6917090041ff2cb5477fdb33d9c6a5ab160d0928a45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7d880347f3de38cefaf5537166a68c2fa75c8a4b357e5846;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b02da23cb5f7a2d5e9d59186c1a00b168f13fbf2c05f3b42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc23fa7e6db0e9c6a004c568f2b1c3f775636366c7bb7c3d7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3931745f4d23d05be66ad30980a60635d2a6ca55ea48b5e3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb832585e4c228ad9f8d1c0ce52a94c6ef86a9b7b69a8e98e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2191cdf9884b9bc56e7b870d3fd511e9beeec1194ae2bd72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he756e03834b1a51b929870ceb079a82f4cfa4ec70ea3a06e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ceacaa56d68691f413e749709357206eaca768914a2f9179;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e6226ac2eb04d2bf3e684b4f68e37943e6e812211c290374;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3aeec9ce89b6d9c1375c3bfb5bab867bba2006e2421a2942;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha82c3c98832cd3f920717f71ecbb80c4fb1f6e67bb700a81e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1160cdb86807899b8065215d9bdc9275d1855585d427152d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30f5596073169004488d17a203e58c872fc6fe286deb46dfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cb18e97ffca069fea833b34055488c5c52c2851c75f9b2e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51415e5286b42f3c8202b1d623bb2020f2d11afa5a5c0ab2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8901a28386954cff705358862dc7194dbfb0073cc871fb08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9e2f9d9be10f3c835db6431b6b1aceba9b73f55747ca5113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93e65fbce7b5798d37da2372db951d20826e7f8be2ea3d311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h882bffb7a4b5f645a5c6667d4022dd324718e6923181fd38b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf1922d426a9098eee938f53c9a1a1dbe1cab0acbf9c3f714;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4c5b4c6c79bd036b491e89b4ee7fb7c2de7a2af10b84d61e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae92bcf1927bd3a0c100b55cf8b27dd58f17829e59e06924c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc240283209ef0f9a90b478acac42815b7e1395d74ded07300;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h990987f50d8a7211ac0391e9b4a4812c7528f1b5567760d3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd46670cda2e4cded95aaba914a6525164e62d11013187ab78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb299eabb95fc7b78af034706e730ab632fe6808c15f92b41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eb832624a9531154039ffae906c7c642b4c3f85ad23fd576;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c5b48e783f82371e683119739390216143a8e8487c3771aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h791d2a8956612c8fe0266759fbf94c2767e540e3ba1f16e1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a4eddf8e245c0daf509b3adb9a873d24fb27fe6ea53a89cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fea13edcb33307aac2bed4a4b184b93d8e874685a4fb2d01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57bfd8305866134da4cadb9dd23bff1e4d2910e7e1bc16c4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3e02e711c39a85e78215692bf701d51a8745cf64162691a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73b7d28704081aa333f52c2c09b1ec660052593632727cf9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h556f8c69bd225341a45447d1fad04450c2a613cd618f27384;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b3cb31edeb68bb39117b771af0be67632cbf386bd02222fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25ef56017799089741ed73ff086dbccb7458883d8edb86150;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b90d83466030de6e84d0852e2eeb7feb777ea8e79248d31e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha98a87cf1d4ae5f7fdb4c4bd0ee0cd1975de65d5b4c5c9aa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59e78d62395fe5d39ecf0638ba15e9f444dfe4e8b1f9b42c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef6b70fae8d50921921969a30e57906545433f94d45a0c951;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7815e6a40a9b1b640cde2489597527a4f0570f88dfae64740;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d05caaa79792d9a8356ca14622d0a72a504cb34192519c92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd0770406fabb8a2c1f201d0f402010612a4320993bc71bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h546413af97b70fa098b9f4c9c2768ccf8c25a511572e43be9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2f7c8e8d127ecf4472674a6c54a46280c021d042d4e10d3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b7c66c1ba285d450e7ea277e37f4dfc40de192ca6e5a1f7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fcc3d3a75786e40bd3ca9d822c254c9d0e01974ebee917f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4b2ba6e4a4749147c47a852d92e74ae560ee5dbd9cdf829f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha10ba9d397d890713e294873e51ba559d73414b5946d90e8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f0f45975ad1340389e6134a8930eabfb1b49138f10a6fba6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c7430c6719fe25bb84a1d0b6209c4b2d5e0f818a627391d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd68b253f2a14de5aeb60b5724de76dd7d3007345f2dc87e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25fadf6942b83716cbecb45bdce2af7e71dc907b57a2659b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf45b7ea90c25a6ef4b9e910c7daaeda0f544cf1f6cd3cb65c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fe6cbb5461aeb49b4c3139c0a5290e6b6dad786588090cf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffe85d8a6e30e30c27db9893a5b251076b1c971d7e339b8b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d8b35e41827f60e65f7c9b49e0e8528fdab1e001bdfe0e27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ae0cf21b3709eb24546d66c44a6fca4ce3066e6813cf64e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6b129308f2620a9635a352e2e61efa0ab4490513c90a6a43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h562aba7708a68dc67e84fc290b507e2179205e4676f348b93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb21d73ca9b812b25beaf1e20bcdd5bcea9c2991ec8fd8b31f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cae71df69cc63312a9a261b0de55ba0ea6a404992222c624;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1277138c63134aac694c715bfb5281b156525eb322455ddd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd577b53ba73e87be1d03fa6afe936586cb2179458c787cdf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee64105fa6a322996b185273e7db6319949b57bcb9936426b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2b8c7af36dccebed3a0612efdc4699fcdc436e17d779829e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ae5f73364ba67e36bfcbe3b1059fc7cdc4bf9e9df82ad16b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b6fae59592002a7395c4a78351d9bbd373d9a701f376898e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2324c43897128ff32e350115cceb5373f2f2f82b995166404;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1b2d325395e8b69a718f2fae6bbadbbe019e96a75257ef36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ae9762d7a37471dfe5442f6f171a2678c20459ebc9944e55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h114fd6e74d5340b4a5038c203abb1d1292ac73c93a279c02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18b5bba95c28e8e2deeaa3c963d1530448cb1bfadcdd9c1a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h515c8390778f7626784e3887723a9176bb2653e6a3c14d85b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h608b8ccd1b80302e0ee611354cf035de8e0e3ca9e77f63c9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadd5a5ba558100d83a0c1a0cf5dece7bc27ea7a2637e544df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbc2d021c06dabca81747da537a1efc6dc54845f23749807;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb50c3d9b6cad3ca2aa6d0ab109d6a199670b70ce2f1d18f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h787b259787c6da44c0caf10b1accf1122569e5fbe024f2c5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacc087da7222b9e61988a9b6df78b2abe0496659600d28bdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cf1c8bb2807fa0d5d719e780d8329940966d6c0f93b85ce1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd736a040e549465ca6448afb396991d800086c1bfe7d5a36b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha071ed046505f198a516b6bc42f41c2f4dbf4c565cfc89780;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3c836b8a024120ec991d615a7d182d68c6242f849619fcb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e5fc2c521643c408ccd1f95b006aa62e65ae6731b44ced35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dcdd0349f4ec0908ebff2273e216fa2cb482b41dcc1eddbc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf176df5735e35c55af392d7506b6647ff4efbe44809ecfd69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e89afd8056128b70b73d08c840c947f838ddf2038b20d665;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb314126dba8f0fefb2b7a1146c44e2599fe73f3d00125012c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb66d9b59a1040f1b04a72700b3827f9f20ac588db90c582b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66b522c7f602866cc039548de3a8bcc0eb98b83c72a4d6747;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6aa3ad88b8d3678fb1418363eca826bb3fad898cf35b8cda1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c95089935961de1cbb9949e6df0d74840cf84b57a63eebc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h470d4c5ac42c4e349c5bbe7a5f82a77d037bd4bb6d5c0b833;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc78eaaecbf9b2334f17e88dc9a94e929f8dd1f4112d66842;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbcf8a02230610b5c228b4b68378c5d75d92046e06bb018a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13f1ef8bd29079f13f88107a14fd502bc8f1aa90fca16191c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9d7ab3261314c78977cf3ccb6d953c1ea41710cd3b0c262c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8e1aa1856d005f63948e14df66633dacd7137311a90ff12b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he43c2afa88d97a114836f4f6e5132409896129d02fe42ae9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3e01175214d89cf8bcbc1aa3551fc82c36902e417b0a4727;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6464d130c26dc326aa8f1397dc0dd10caa176e3cbaff9507;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb55c6abd7df92f0cc94f798e0d9954827c777ce4aaadfbf9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda7388419a933d0a42b555318c1eeb72ce5fe7436363ae71f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ade8f4dca205d3f5c2250029da3104eea5ebc282b762688d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9b7d3a7eb0e8a7cff50b13fd17a42af741cb5e23821117c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha70281d6e3161972fd82f959a3f1955249e1e7761c91af826;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d13366663d52a68bdd22f19d6f6db3055834f0d276768b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349596a0bc4cff2740d9e3134492578fe6d31dbe59617d090;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff750adcb7f66fb437421d87d7d70890a407d7a6c881ac700;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74f20191f516488e7d875629b1fffb920f7b6cae175bafad2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4627ff91b8f22804452ae5791b52011fd026d686fb7bc5be5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8826e213305e30b2bbd4287fe38c59672a2a27a781baddeb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98a3704923ac8363aadbe1d772778033075cff2b6b90413d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5867ad402a86e600f1f15c66e2cfc6dbc98dce289cd36d66e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he93f397c79c10955720e367be0d5a6166944a9c84e57c3c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6f49423e864c5986cc3068c4bae2b6cd61ae25a7272484f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc750020a16e316df08b8a472808316d0459f922c252a8d5bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90cac9942afa077a6ec240ba2a8d91a3fda62cfa000653767;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd0848834f2963d47513099a78b2ce17e86c203d65193dc39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd112c542fdb24fe626152d3f09e6c1e3ea5fb581bca207f0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h292a50ed488e7b31e40f40557c6232e0a5923e8c770fb1f27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9471474c8d87fe1d16e4e6d22d737b1569cf3b7c4fffbb3fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe61b1cad8383b83e540bf3903901fa65b0b3c96152a8e2ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27d97eae538d8e089da8eda1b3846185b92cfa20ae10747dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd71947226e547677cfd67315c4f07e58333d627fcc62203e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12f5e96f1455c0933ad7addb9077ae71fe0343987605e62ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d32e05177291e4aaeefe38b171a6ec4b7e0302fb8dc61220;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fb1c60d5c09e8a5cc311c47993fe4590cde2adffe3a4e523;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7d36a4708baf40cc323582a4c75213971d6a9db2f9838013;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5a6d81da7a942c337037c8d0f83490eb649283341750122d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26e22bbd7a9a3e03519ba6b90d0d6bbc17395a1ec08faae32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8849d3de6e33c075d8805518b3b6227afac2ab1ea7deb24c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e744ccea8470fd377de6a0eed5a53385e3308655905a7566;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66881c49e07a8d38592698cc0ee4d43aed8832d616455258b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e940ed2efa0948a1206ee6447d2c97ac154b82131cbe391d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h801e45bc18f087b5e10eed114348ccf02e5f6856cca70152a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84fd6bc445fd84337f33bca8ecfd859d18772f7eea36a1db1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bff9bcec4830e9625c24cd6460c2dfc28baf57bc82690040;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h318410ed25ea5532dedf27780347bdf6dcf6a9a2d5ac10a81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ac89578807c9d61295565c8793d1cc8f3b0a4973bd540622;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa44d5bf0f526807eaf8bdfb1ca78a4485b4271078ea6966e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75879ee6c6e5ee4c7e4fbe027f4564e5606999e66b8efb2a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4201b7b646bbfd1b5948f6992882ec63d6ca7b795fcea1a35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e442c37d3580e2733b5e507dbf6de7cd70c6e0dbdc9faa90;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60c6dfc359c42f4e7e3acdf659340bff2f7d650b50df8d8a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ed31ea190c1be1758d2d88f1a7e0b0e812f01eb840006a16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4460a46cc889eea5b589127585e702d89a6c52f5b520e483;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73f35c5021983a27aca7e5c960acbbdeba0da0bb8a3607d3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7a2fa0125b13d6e4d81482cfbb6ba471290a0a1d7cd942d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h957637aba50de0c6aaf46ba9cd67d661540fe08db97d4bdbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92227b17a97a2e3e3aaad8b5156c47f9b3e5e483297e13bba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44903de3a29885a66d214d4f344000cfd8cbc63fac0e6a7a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12a3bdf2b95c9326d8f273735bdcb8ad30b28fc5c66eec1e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6c266be11cd6b938d83adbe3ac165569e005f35af91114ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h264181e2618295ca331e48d8da2949ec6f07deee96388b49d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fc5978075c04656716182ffd4fa97b1a9ddb1b8a92609dd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h508c3cf8ddbcabf0ff71389e09c5d1a7fed9f19cece8b736b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14a4684c77ce88ade5c1009c783232a9d6bdb7d90c26ee294;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe67b7c2ebbb2553ba7961d94bf1b8813584bf2a8c033d67b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdd827c334e686e88d25e81704b79afe4027cbab9a56fbc8e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h552ddf336f3def619392f021fd0c52986e7b455eb0ba47bdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha09ed3ed235dc1cc465ab6f74c58467d4930a4929ff15b36f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ce720993ed4190ca5c7c4f0d21c2218543656d382f3a674a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h380d7e01aa8e402834094db26bd42eced0e4920648095b0af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25da403ae225d6323c854a65509ede82ccd01a388aeeed290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h396dd2f5eb2f590871cb2ea1683983450a55ec93c3c3dd38c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf392ccb1392858c85b2fbac565fc135ab4f4918ef9df0c425;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha40efbc78ab4fb3c99d3a42913a7972ff9454d2cbb6349154;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a196972e237fc40fd92bf74db064cdb41353a772b009c5ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bccdcd5430c8c8cd812a8b1621563fd97e14569d3cfeec6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf33db445551c4a77a8d1d782698fe7cfdcd1c0d2c0646a1f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cc465d05a92df679d80b4988aea76c5050e2f6ee66636243;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c366fa9fc17df0561143fda9f3994cfc7c0520b79e7dcaac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd626b847e7e1cb3f60b1139a403f1803aea9d27f86da04d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e3d079c8203b14211293daa73e33d714854c999e08d15ad0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd48cfd01392a1400d158b8a9f98bd238bc60f79033a9bba13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4da1325f25ee2e2f0510f957d3385d206d2b678ed95714eb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16ecff9b435d8c50646542a22b8b7e0bc1d036369dc5298dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3729f3b79ca0c2264be95947c1b83016dbe29bd92673056f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5384ddfd71e2fff9637a1505d30ae9c2af2a16d408117ad1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84338945e2c855bd626b5794f138293883aa231ca081c13dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25835e8a09b6aac97442fffc73d7e26b88326679aeb150f20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37753e7b546ae977d6ecbd234788beed024f329d0aedae8c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e2a417e138d0a24862805be4b5e19ae9190e57464452dec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5b487161c8512e2680ae7ef5a3b9924f7fd44d46210319c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b2a6c9adceb1e1b980dd05f58dfa9e67effc3a788c2e60ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf439951a108e5fa92a403cc3585defdb0674eacfcd076bfc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bf86d46debe236b3ccee7c740af0ea5fa25730640f28d74e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c894b70c3a590d661c826b41633f49d4735baeb141f6d3a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha377c67789ce08a340e89cf341e576aea5b9b483fae8fa7bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5f6f7e07d9d4c0247fe9c8db51ff38549f5ea719187aa65c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h699856f1c6206ebc8fde1260b2f82164f53d504c9991a5910;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h621d960e1a571860d4339f8a45cfe6d2598fc96ca38af9e88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h149de5548bc1216beae4c49c3a436186b817969506a9c822f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e1f9b530aede916f689101b3b1f90b3fc2a8be46cc67fb9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a0e11390c3d34aadcd37c92ac4a1926c85e6eebdd61998e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4af7a49a937973aeb5ef21fa33c324b425ced52c65ba1ff64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67fb3ce28621e785906faa42b3a67d8c7bd892fec075709ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48c757871e39901b4ddf22718001d2a59cb2c0b442d42dfd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc27f8badf33dbf22ea81ab7789177a125dcf8f225a370e6cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h307875571bbfea882a9a364bd0e620e38a915d204d9bd23c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ebd481ac10684a4f087f4613039eb151dcd03a7a6283b7cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6022e2b866ee18b6f612ee5208100d16365789e130af9d408;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha77404b4d5e70ad25041a93801cc6dfbc080988d6b676932b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7cf9667e1ba0006e3945a1ac5ee3aa40937f8103886fb413;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b699201ca9dd031b6cfd41d0967407a86635e7921dba3984;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c8b447faa04be27e83181b16ce4cae4827b03970e4a5f253;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5b17d45e45641cac4dbccf749a3c1bbf44ec86e2cb529e2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dde528faf91f3684f312fba9b08f27854d1b778e6c6b2973;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcef9ee532523dc27111778a046dd5f2052e093d21c9d4238b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72148d75d7a261227f8d66a0a9611ea7577ad47390d9e7e00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b91999600c9dfa59bf73750a7af7575e0bb228f5086674e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17425f5d64e776f25672525b58b403a3b1c01a95429b901b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he52dd098e14120161a86d16c0ef54864ff167917e6f64e4fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94f98bff8670f1454adb0dc410ecef2d6071ecf667d2dded9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71117ad70e65e74cb5d6aa6b3a99eecb523b90aacd4b453e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c2ec97b40beb4297bf228654010b2f2d36c7d1a2d2608e39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1361354e8a7f9055c89346345adbdf8432b1305f900d2fab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc8fa7cbb244f51095eb975587c60e93f7c16aaf11c74a41b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcba1ed33d88812251135ba666a4de33a4c19d7ca6f1916e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18e2a93892aa3a7019342ec5d8e27063df26f601794c1b196;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0654d400dd138c0557e96d9da1ecc4a8a74a0d4bab06fbfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92c2f7348248c640d654fcb76ca5d47ee9016b9447b947526;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he725c43fd375e446c6fcf31de15f29d84155451212b3ab66d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc01cb7c893c5a9fa168086567f4eea591e28964f86b7550d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa6c273c1b336afd5a1716c1a541586dd6961c35bdae3e535;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e6d7e414a2469fd87bdf90f62304996d1ca966941ecbd0c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4790156671a5362964d5de627eb810af0e3ef7e828d43a483;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88b10891b6ad32ad9744b78d965dc80e5e8d124640f9a13ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha489466fa55e0147a74d8ca8b61128873af6137968c88e26c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf6e444afed2b4f3f01b8f9487d9fcb63fa5a009a7edc9f36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84b6689aa9517ec1e5d1adce90e644749de28d0e29a7f29af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10a4ebb23ac4772a37f5faa634658092bda71a736d9a3e608;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72df7e8b6cd2233713e46c1f1266f53bec77abe543fb49f7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha02ed7ee98930aa865750b36f24da25031040f7d3c2ab76b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3958792500c24e786024aafbe6318c8d9969116d72e9c2dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ae3d2cc8656247fad68499986fb290f0bf154fed8900bd4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5f6eb3163c0d8b0d4e8118abe7add288098c3d014005ddf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc97613bbc1df56f9c59c08b92020a7662271d34ab8368425c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc11b4c5554e8a9c294563d488b53d894f35b5fa6561b09f4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd1006b15d6e1ff608801ccbf30b4b93eec9df898a0f0ca79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf3285a349c00ef328da76c749ab02db47f7df5a1f05be282;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha23c71d9fe1d3c61662cbf9811dd9b01e4d8a79069493e5ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c04e4ca8ac9abdf95824531932010083e73660e7bb1e5a45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cafd5f9bc0cc3303877df5a85877d7d89f63e7b15a7a38dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b30a837b4557bf3072add9ceec4246a27088188940a1f9a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haebe6853994de9d13f5df9bedac12d0d1ec140cee6c95d227;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h949e0d410b5ad131e6ba6e841690e1cb2878218e49505028d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a71ef3ed85ffea7e805b97985be637e5b297baf07883fa9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h910e02acc7f8169d3f350aba1a75bf3aadcd0fa96ba83ceb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56e598c234cd7c707443642fd86c85e142fbd4c9f4e66549c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h800657acdbf3bf2ffab1017ba13c2f8938a1d422bdaafdbc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h536f206df2a71fe22cc2a9209333b9f8d9a05ab7493623946;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71994d9b68e2d1ed57d682ff7eba1dc6ae8eb983c7de67012;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf94664ea1920ef7e763c743ff79ef4e5a07473e3d41068153;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2c163e8bba3386e3de7afbb8fbbac02e9aae3ed2f8de6c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57812d5123bca9290a1cff7c9d26e10ad07f361277b6e76a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha45c581ce1c5c355e9605d963e730f05a122aaf932e7622bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d0d232235f2d6f76528746255ea4520d2ac2a97879730cd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1de26592924c9ea0f5ffd859223199f9e0cd1200b20cb3e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23061739ae8c08a362c9416dc671f9aa9417474118115c6f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84c7194d100f69f3b031eaf73e0b735ad255b181f7283195c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee87f473d8765945b6ff60d8e8c95b54b08dcb3e12dee98be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6abf30a4351e3743a2ca3bb861838a383d46cb75bb63d1c63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2041df240be37c2a33f68888d0aa4b3f632591c8258aed070;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f3063997cc4ec697bf0b45db50983a119571509a381759ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5498dfc27081211a4132d00936158ebb05c282aca251a30d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d5436222a13aa037351c7633e9c9434aed2818969b44862f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44a01a896f02a0f41db5a86bd0bf67352fe6b16d0b293b70b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fe16c934a0d43c3d50ccb7283d58970e5653fcaec118f325;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90a19781915bb705fa6f103baf77640f3f05dca8ae8a1c7fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb76e2361e7e56a69a0b9c678218e707fb29a7af49f959dfe7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1fac60e1f9feb34d964120f99fb2c023e1e5925007069889;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ca038dc8c8f862003686177c240c9f93ab4958344743e816;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd2e6b6deaa33f1e57cf823b8eefb5c49c3568614c71569a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf97fc35bce5e1d76f5024f03d3d2f69dbbf95dcc5ca44ec48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86bbec3360ef241946b7f398a57e85433bee8a351dab47759;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21cfac37d8b080f8a361b433a92ba29da1e24b500c9a410a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h880bcdfab9d6615b368e16e8a17ef413c6b5ae699652d7ed8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69966e383298603d8159a74f5ac1ac477edcf3149fc707422;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8796dd6488bfed69e10994abc83726073546200adc8ba3751;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h893a32451a7ffa510b184d13a512e8ace7f23670fdff8c85d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h360abcecbc1da2390c911e368a242efbbe8274d8f32e8f393;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5057f041863c3cdab9d0f27a9f39d289de764398b6ba7a1ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c90203ce2dd1343d1f82f0f65736584e98a85aff407aa7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ade8ba91546233eecdb9d7a2e263b636cab171db88276106;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c11cfafdfcad0e24a868cc2ecddcac7a20c5ac821b4f1979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h320873394bc6ce98ee8ebb9a72e926a71edb82281b6050bf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75a4580ac95e76ec51b1be0b34c42704449fb507343ef2e9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77e72a739c1a0d6c1f07ec277f42e34793e61dec1bc1d87f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebc90ebd7573445baf224c85a18cc4e349db507cf9fe92b3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7f81b762deee9bf584ffad0c8d15ac62ea1886aab7ee714f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb20bba06bb11ae45df0a4ac4b2f9dfab06777a347d5d5a8db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee90acb57e022e46a7340e763b32e371a922c84d99a07399e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdde90734da888c8a38d5836ba75c9f4118edda7bbedc4b46c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63ca1fbb882e831c3e7ae63723515b62355b45bc2c3c59311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcc3c622ee5ae72e8dfca81f009a7e34bb9f65631c342e6ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1c2c151b8d9d6b124dc800d64b81cbdf59cdf0072163c83a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e3b44d7522082a6fdfd7d969e3e580b81f2935126d4afea5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba1f8920a788ef3864561c58e66246661312295d0a7b2d6d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37c27957ed21db28fff56cd332ab1fd1013d9910cc642e75d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he003c8a600b81a3ddc10d915a01a75f5d34e057e5ffd98c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h397ecaa203afb8369100fdd58c15d8d5d456b1bee96b010e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8ec74b2893bbc534bc6477de6bb5f10ba66f6ab86576ef46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h790d8a119ba861e47a41df246aa584b9226ac3b371eeba956;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6af336856797cf768b16984fc55d519438380a5ce34f308cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h849be80de720976e03c1549463b62f15d1581e6d77e6523e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5956c9f2ddddeb6aaf5af30d4d6db7bffb975599cf8b301fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8521fe29d7e90bfff9017701f7390e0df81a8884cf76d6f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92aee4b510bb9a4b387a58d4c9855ebd25487dd712822ad6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h964f57b58500474fea0d22d537dcffa15c1c3a574f2bb2673;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bb1680e2653020757179e971f3feb7b32092b6d41beb07c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h871610368db0b6699c68d14446d58e9d87547440515d8fa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0831d4fe4b65634fe9e25bfe9bb7985ed8cfd93bde2f7cb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf42db7a64b0608b4a3aa38bf6dfd67262e65bdbc2c2997a91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2251ce5d62ffb573d46796668bf694d67bcb741e23a3981eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b222dbaa9451bd788462947a8148147ac73265d507425088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77ad5b982668458e1ad86e1480be98448e578a64d7e54f507;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9b78672fa6c5a0903de3e78224c40c0332d4fa3b49ba14fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d389438da47ea0a00319789fe51aa3ff8b31e688846fe8d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8634a1452af8b68e68d680d62d24fdc171b0919436564deb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed456a9874ffd9cfbd14bcf5fb8dd8eb75f963bd6a074e97f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d1a73b1434127f2a4e013aafc40adf4b9d4fa666e6481aed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b64f348bf5f9cf2332b0792b470e13b4b17dc9b77d6ae828;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d6e899ca78ef447ce4ae526b573d8eb573d8f4e82ac7c71b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fe3516bd13627c4d8b487663acb6f145d850e8dd52858b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h231f7b5e4fb52fedd7c903e4c706c847b8a5944444622cbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e81e877eb3612b6a6d028500b78f217528d3978ffbc0960f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39794ef1506013192c4017f0658767796e7d8445c5c878075;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ea091de3e9a556bacbbe458e49b33f04bed80e774b04b0ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha20c9abfb2390f727272e58cf42f86e847c4b1bed903bc8d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e17f57cc34f1264cf731cd7d0e314a755d089d684856eacc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h949d325db537f010401b4e83c8a3cd32e2f32903efa26e300;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8175c4f46497286f77f0c203226c2e1578e21a281af24e028;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1087103dd826980ea730d062c2dc8152ff79248996596571a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ebaac43a8b2dcf5a4e208a348d148ccf7ea52ff6f691951e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75cdd349f48b6ec5b8c0c8fd335cdc537c50da8ffafab8e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b2c764cf256adc7413a346ba7261b246902b39cbf3b9e13e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2451df45fd982269b58fc806108afb99996bf28db4e68b60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bcbc21cc1d6a5f0c27554ab76dea852095a1b46a4228f837;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97913cf3f25afc3a48e81bb71ee59b473af862f1ff74b37d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61399577beddcb5caf6d975496ffd9e4ed066b3fded5ee52c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c439c741ec150dd98213b3cc83c225ba0809b5e1ea1841b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6ecd7bceab7c0f9dc08dcaeb0dea0a17adc93900dc540bd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67e17476e18a7d6042b65fc9b1f8fd8107b2ce0352928405c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haab52fc1160cf98c5c9765af07ffa16b71c7444dd75a21ae0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac87b50822927ee1ecf3e7ac59f9e8a2a5c5e65a741460344;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1d51636c69622d1c61309ced6d86d2b2fa94e3630c2d4c84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5d993d58ba28ec78d3bc3bf015c8eb51052f071f3919e7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf30b948cdfe6cc9faa6708ad2101a4afd06b643240070530;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb23ec22b7e43fcc8b86cd89a30bc6472090b9fa79e3bba52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6157180f74b53585da2b803f76e5514cd125aae23b199df71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56445c254bf45f94f85f7bc5459ccea4242378de7ec033226;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4bfa300e5e692edf7a0f06831e6be5dd067c5b382db986e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5662b2fd1da0a54572256a4d812c154df5b1b9e5e7d763805;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62dff969f356a1468e96fc507bdbe6b3c96ec0a7837c36349;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1ed250875f8655c64c15fd47250526cb92405f8f24b6e5a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf34b8a11b40315996fe49a0ff781f1f37b293e2a88a12d70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4d419623978ce7260f8b818cda848e885b7ab19951dd26b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb57ec985cd4acf52a93d04b879dbaf9a67d5ea6f4b2425ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c99e48b4ed445e602b0c2b3de61c88dabf5c2acc81813099;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h347181774643dfa51bed1c84bbb3ec760a980beb0e0ea109;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f424b123543915d3f54d0365b6f5311b3e2f91505a53a0a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40eb3ff389b815423cb2b2469a5894af03b4ce827446dc9cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f53d25239540f47803c280ca6ae180e7001a2b54180063cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8702846e3fd1b4de6d150e90dadf032b5889e99196ae2b3ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d4379dd1ca3a558c0e0563255acf779f5a26d9d407c88917;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86ad1a5b0a79d97df0703871e3ad66b40f43c7e960ef8bd0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h869fcff667bb04f2f7f4dd2365079db08d35a84510de168ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c781b3c3500b773cb00ff669e2f499c3fefb11f0e843b7b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63ce6df8a946036856e169b43981a4f3a11aea574a39c2e0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b13be9e08cfa6f5ed155141d1b559d97e28ff0a363b07322;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1dfaaff6635a114eda00a53964a0336783dfcfe97cfe7f4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91d573268e7637459d6976c2b2a477b20c2f0c68cc45fb2cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d40a5b9fb70a763868623df5a2c50b9bbf09a0b44b11cc20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22d02f6acd937efd020ced323a702c00f2a831787c38a0083;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70ef395785992b44f8c72431ac687f4327fdefcb4a7b8009f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcda1bcb30b0dee362621fede235377192532783e381bdbd95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64bc06349d781bec993ef40c0c52eba547112ed27b83b243f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e05d3bde876277a8d6df3607ea7f0da0c32f02700ec90ab3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d03e91d1aeaf63f6081ce443ead4813ef59f0dd73571d08a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha001876d775fb7c327913c23788cca51f8911e4221a57f2e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a48b356faad9702cd7c56d4820396a5a2886f3b8015fcf1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81bb1b263f1207f2ab123c31c1eb1e555912583af40e4b438;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29b5cc3a6a144661989c1dddf8dfc771b09bffe5a1f5fdce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h262cd17bf9f6efd798d62f9daf537da708f65e632c15e4f00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4633bb594a39f019ba78a79e97f76b10942182766f14e731;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf6d204a8f7b9c997d04ca10f4c7695665a7f9fd5cb753296;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef54c57d84e22db5df9acac0d6380d87da18296fec534c854;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdea2bd2c8d42caf38262e832b81866630ea2cd5941168f618;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3da12b7eae2a62e32ff11636b70223986cb57ed846f583777;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb19bc7f53d782abd01f5972124133f094edaf43267c8942dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa27c162d94917b4871929fd85782e17af71d3a4be31095b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c2a6aaa76358baf9e1285e0bba72621c4e5120d6a20b1845;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59f61c52ba9efd0eb2d2ffd901cb75cea82b2788264ffc45e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha175e1fadb9a91090d5fee980264aacc5169cf863f2993df9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0c5c2763cdb29960113a3058bdcec57f17ed78eb806d077a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5af8581b529a9f4a799458b6f04eb56f20b647475578110ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f4ef373939ee7d10a10d22ef85c044aa25c909330a1305d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c6090f4087d860f0875c4dbae90e660573f5269cc07e51b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd794a1a0c889632d80f4f02483c7237849c27ca8c48b99cfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea9c1abbe3a002f12a2c9baadee25ae05591f65cebcf4282;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h164b16aad2cee9192edbdc63d593571ca027fe0762963d2a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h896a21daa1ea0fec04151c8a8ffae0c161d7f8fe927e7420e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h980303e0f5eb8bcf128f4331842c22f347d74bb0c8ded6038;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2884d34f50f995b7b234b81a80558bd181d9ae798fc02dff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21d5c28877cadb106146d2bf71bb05ead87cd902f154fcf61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce9f2031d6c1723673ab1779d2e4f16f01b1fa68517ac6c85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9bb6cc5577c95bec549d85c3eb9c3ddfc1c4b3d078202ac4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4aefb6e941c26bed48c80edda96ca1fdb2a4aff5e8490f5db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d839770adccc39bed4348fb299f414fd29d4d69e12ffae48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb68c2f4d457a596116e8b3ceee2f48a80e2a7f205197ef76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20980feadb4181819fa225f9df539f3721d66984b3acf9eaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h944aa28b30b804b4f7534ee7d6f07652a3a938968efb217ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8f01bd158c60ddd8380966a91655bd4ac6951b08dc90f3b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef2a9ff070c2140bc7862004f4ff0d70baf299b276f39cb58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef65c9ce00a1d54cb09ba4379c65be6c5b99c8261d059f81a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5bd5314592c7bed2bc845092aeea9bfa6768e2c1ed9e6670;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d452bad5adb888b60480228989a5c3207a5d48a766b744c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0e1917a01376ddf319e96be4872908de77a23d0594c4511c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7144e5d46f2d1740c3a6f1d05e8a024b4985faf0ac1fab43c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92ef2a9ff875b5df5467df9c6bdd14362c96cf13dcc3535a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b1ea4b0d7c7f4b0f4f92d030a2cb5d55adb183830db5f91f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b872d69cccf2e6277af502dc875c343d910f6dd1c2342183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h856ed1e0f7dac09b7612a98ac68525f4d3b4a1662669050e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6588e6c13ee9166f931ee7aae01374532752111b75779f66b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec5ffa045df882b106b6c1d37de8867a45ab3ff7bc5cf2610;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35ec21a62fc89a031bd8fb28a817b69cd194b84b85a802a24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc36df9a058909ae65de5b7d48c40bdb02a039ebfd255577e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7600514e5a1b79351ce370c25827b0d10426e553a7408948c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e8a6841280fea80662f5e8bfae7a48afd744c380de5f49d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h312f9ae357caa849206cdaaf503517be02e00b588061139ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h916b67e6875da25dad554e7d7262c24a433f27ed4fae79027;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd457125253c3adb8651183e2f62cbf9c67e35c2b563e1696b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e8934f71add56528bb71fbb80cc08ab016406f2d6e9b1b56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15aed1c645b9ab2acc607efeffb0917c536b689d4aa0fde6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8fafe01c564662bdb00ff09829bed924473939a214c8e155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2369dd28309b042f106587a9033c5e5c7a5a3ceb3d89933b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcca6fea0c48ab0a50a5ab7c9279557d70c32dc273257cbefa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b32bdefc7a0f3b4871adf05f811bb9ffea8d117bfecad90e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a5b25b97044757d93ecfcde9ae6318d6348cf8e603eda61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51ac081292fcf12328eadd15ad010590c2fa27f68bb44b1a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab9f2a46dc3250d7c6b8337c25e6c69ccc40a68b20bf2349;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heeaca28b71c07004d517400e9d0db8e8e0d3eb301377fc7fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h799b91d6e6b23ba58dc4e11deabed5f3477095e880cb84e79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bf4ebe32e16385d8d8e74d30d61e5dd1e365bb0e857b0605;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb951ecec95c0a81866e56a8bad2c178de9f51d60ea0b7756b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0dc459871c944c647f2b3873bb8f345580c22cd76b8a9e8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b2e03ce8604983685932a01afa2b853321e76feee1541901;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66ba7bc68337e1995fba390618d9df1a6ee36c5334b5042e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25191778d7ab772aee0fb42608ed542b1e3e97b74d033c676;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9476792d649b1da87bb020c7957b32bfcfffa8e12ec6680cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c001e28bb3ad53e51f1519f861801a4eccd5fbd5f350b62b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d9208a0dfb33c0bcf8dba6984757edc94752442aa6c930b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he93b22a2da77e77e822960489e6a59b4156e27d3d97065207;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74f4971442fa4166e06cdd8577fea098d65231aa862659e7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc38dc24786997731a4eeee2e6483ab9bf91c69697fd1e1a55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b960c7ed15059fe14a7ae6cee1c5f11d26376a0aa9ad29cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42a66ca99bbdfbec876abafc7d0b53151dc83d83f9117624e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62fdeacddaf4d16958137686295242d80dff6d65ce82fb53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5e17191132b5efaf8d5244c837199a14a2b690c9aa08b6a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2700ce1241f31dc12693081b1b02c28eb60b8db3b35582db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h862aab5f1e886477b593554a09b60ec4f8976db6235dcc4f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he01672b66951049e5b70c95dfa994962bbcef165eb199c926;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8143256cb05f218393247bf0ac634ab9e0eccfe45ab41605c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c4a1d45112ae772167e121768002ee53f573d005382d3dd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41248df06f10fd01581a975d86b0ab4213db8d7d08936f8c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2afec7adf5e0ddbab0000857f5c6c3dbe4f6e67ffba7ce79b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20e5aac0506ff06d9568cf82ba3520e8c211db087d8694234;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h279c0a7f095d64b404f8588c48055b11f4b95f2e8afda1f1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37a42daea20ac7cb2f059cff127c51adf9ebdeb7cfb017dee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h216eb0abc8b499581caf31e441413694462b820a3662e96a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a984d852ec23d7f157ac4271ce8508ba6aedfcb819e5a3fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fd678d3ec46e1fa4d512ede5d1d6c048ba0de4f619964d9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde12bfd57cea009c625c84438fd934660581f95e3f17fa763;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf8396a26aa39f7680c983fdb4637f1b2c971af8b4c3a7adf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c7d4e86d0c1f438ad9bc109e31152259061be0369bf724bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d4174d7df900c91b3287e3d292e023db670b4571a7bb266b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15fb5d6b6826738c568c1da13842374f2387a60f09c74ebd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba8050f608f2f9bea71e0a120a10dfcfc2b779e3b194f4fb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5997f89f2dcf4176f799cdd69c24a9b19dcf796deb7be2be6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfeea30e4ff07c2f710ce9680e3d7d0a4363062d7d8f12681e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f72f227ecd3d4e3cd8a3d841fced2cf898633a5db51b89bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17c7d0817b779157ff0dcaf7c3f58f8561e8c066df67a2191;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h770fb32e51e9daf9bb7cf3f04fda8cf0cce9d4be6efea83d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffe0eb42aece79c13a0c47a23cfbfb969194591dc91914a33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h725e9856683781a0bde461d9b733bf374ff9a4be63d1816a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc25c9606128d1053fcef9342f5d12e09a2bbfa64e40b5da2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2149e251f6c50439fe63b5076744f17c2f1747fe8e61b48b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ae9c801380c084969d8aa11b0141e4283f93abd7a25988f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c634b66b3de0e00377e92a078ae5c10e570cd121a6446563;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9bd402c46332a6e8ac9222c74cd08ce3c88419d596578486;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62efa59a48726cf9b04350a2a644e776231a6a2d34df3812d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e52a7f93c58a43f25a10514b073db48494f68f4ba70e18a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d5dc54bea6f677654c135cd9b987d5d885c2ae1c203acc92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e9ddbef96300674a58cb99e5d885d4ebe84acf55e68f7b89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfee5c1d429389e453c9eee756f4028443fad115c637b60c2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5858d48cc2b70797dadd31bf4b4fd8e623b490173f7ea83f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b65034466f04f541dd4827d009343af15a7bb3ce73c196fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34cdd4040e7f4f72bc0dc5a666e8ae2f87cd6a8a672c2925b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4954ad77830e2608e31b12faebcad4362a7fd800d458dbf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e55b71b9f4a27d373dc6bb7993f22f91e43c8c2952e2ac5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56f8b0f8a3be0d400edbf7a8f20e2289a160c5dcedd9d4750;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86c4b3dfa848cdce5961b2473e38798436f5c9990b9e38175;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb843aea87f9e0df35fd9d6fffd81ae598fc895d832dd24786;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f16e8524736a6591219322c03a580ee437543bb94cc58147;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f58471bc40f3e0b260e844ce89c2c7a8aa428901c682b2c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a2dd80c1fd29ba6fba1db3a576371c261a0eed3a1efdb314;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f4a774e352fe3004ef844b4131add38ed65b458545813785;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5eac0d720845b5a3362e570c2be802ca7bfdfc074710116e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61e89fa55a6399295873bc59150f7cc354265224235cf839;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbc2f85003d40149e6677d57d53c55be08452de56593be973;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6437e8397c011ab584323efb849a9ca478cb592f98758f8fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25f667c760ff57b46bdd22f8ef214e10120bee63f4a58433c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2163c3ad64f060b3b699aebb86ec8544fe9e58856349188c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5ef379e8a26fc57167756d39d70d4de576cb9d0478d096a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0ef123a87b9d99718ced1fe69b4f08c3c1c8052a2f8b7f98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha958f36f7be2f19c9a160d249a39575c5a862228273e9ad99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6adcb900563c85a41d3cfbc4ddba823c73f4e4ed47c574fa1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53bdde5b312ea1326f9700a8096eb3c9fc08249f332f056da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5877bd058eb33af3284d537bf326ba1613eb6e39ab6258549;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h459e69f289e196bbd3f3acebb538aad9363837fb263125867;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7d384c604381c7e40a56e14f9b2fd2ff3d80452df247b5af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73de8cc3b0fbcb0fde5ae53875c2cbf39651f4997b0411e2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h181c76b414139b98910503f17b06148ce672fb2b1db6b3e64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc504f48ba125d13c245f052e6bd2b37601c998a7d43c7af01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80a6d98346400aa2d6e1d6d9600500c543cf2efbe9456c137;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8acfb638e5a1a9d1fdd20de588acc30eb5ecd6dd1ad871eb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb60a947efca5bbfb79d0649def760b3ffa17cb7bb4423c54d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cf997c938322bb6acd6f76347a0f3427dd2bd6387cb9c8dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he332b844c658f206ead819600c0eba0595d05e87a1d98f989;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d82e04087aa2677c557ffb39bf8c64a7ae01a18a94da7823;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9971bc0ab8aa8918906ce1959349d2bd3c8dfec449293b91b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47cd5fed4eb70f5efd2b18299395807d6eea5e2713c8466f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41e69e1dd7598b332bc7f95eaad62ecf2b82b6de8bdf9a648;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6720ff11edcd962aca85e689de7884d470f204f56ef620757;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44d45f09255cba25378f370824383fb1564bd82318e036f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b1e7cd5a85ba15ce1447b24f2f63e4e4b552a6a37cf3da4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h206c65cbdaf5114910a8b533b023e16f0836757908c73356e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8996f30d19f1ed49e7f9823d33d996253d0c2f959ce4692b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he141899d3a13ab137bbfb457dea4d2ea696ae606506a8c311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc66a3cef17bd0d7444f99fc913bc4975ad2a275f45173dce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb26c8fafe812af7d31c664bda6044f42554b2e6e5aea66d23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ad0c1b89613110c11abfff8edc97f537bb078d4662d7e230;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed79353e43d4898af7df6672d326d87830f7ae2acb73ee489;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ccc3f1d03b530ea52ff66d98039f8ba6e290d6995539b606;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdcdecdcf9c7a11b3d443128ce70d1d0b281a8dd87302cf98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90491c86d76198cc945d2e7bc09a183f8b18c77c0b2a8e280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b2b53c3424c92bd5d3d2d6ee2483c27d0dab832ea8b134d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2d1ed8dc1d2cd625c3d08c2cce74cd197f001ac73ac8a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfda7d15976f400221c33b0dc457ba82223d5d186bea3bd2ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfadc878fe9faf6e90fa8324156e0a38706f34ce45d18cbe93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda0060cab4ad8de47bee8b67a2d352991bfcfe9a3b5a5454;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c93f2be35a917b028e31a2161c61ccf1144f7b7d2470d7e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha12ecee2d95654ff14f0673be903c64240aa15a595ae0163b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d7e7f770f5ab69f7539a987b0a014620433b2a2c9b4972ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67e4c6d94d1b7c4b24f16094953b753027f971efe81179daa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb2fba7eceb722e725d82707561257cd987fcbc321c77d460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha944f7df329c37f28353b1370d352aeb0169fa0524b7fda8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1800db9fcf026fbc8016ae9c8bf4e496f71f11c6091db373d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73cf3a2277036433a9741b76977bca9811dd5ac6b4152f66a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14d72248bf54b37fb35f1fcc04a89ae9e4cc028dd645582b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d1ed738e39c2a2e5db8e8954b98a03a5a0d4605c80a70c30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62f97eb489eedf97bb8a655471649192d04a8e2b7a69505f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h544ef75b05e1ee35b765b45e0752964f7b1e7accd258c5cf9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82ede1755e242234039109d5a2de440525d8fb75aa601ff80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b90e902c10a47cbdf8161c6878b0fcf6f8f7b6371b9f12f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea9b8f09b9d4ac6c81fca71ce97ce0c626a0cec24f3b3141d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb12d3c7ff53112aee2695d29c405240608bb3284ce081c76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c8b0e5835e87e02421eda5e5be6a79b125c1995cb2083afb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef2cf443e59a97622dabbe9429d412ccb35dd0badd419b78b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdea8f9803f1981f6697d117bc45a078240a22fc0d29e04f4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h672d451461158cb31a40f52a3e3f9a0caec8318291d71705e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h252f3d96c8d2b9878c0a5e022c3c4b05df9ca9255beb51e16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb816d939397052cd75c9ee4225536189a2e82e18b5b13f517;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46169aaa90926a1b76789d33cac117a3337756d8206e6181d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3ed55af5ab810d0ba83d721159294c63031da0e9571288ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8682afbf189a4dd98908bdc80de52d587b681431bdb0ec6e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f0a7ae72254f8bd3cabf54304b6c1015c112401c2570833;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3851cbdccdab080c7339d5b2d458609822a93f21cc9ac3598;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h326dc08086e9025d44d9f6b1b57578ba6ac125b944488fa6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc73cf3bf0e3158bd0fac690ba5f75c7ba91c72cdb9310b4d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8158ce64923eda0f2688a4c0b7e8ab65cef0c9350b950a6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h251f3205157ac8f51f2fb014f8d2acc8b1a47634dbe6efb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97701a57ecc1b23fe76ff2693dc8940f0472b1de4b137a91e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf111f5b2e7120b525083e5eb525935a798866fe3d9f539613;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f66faa589e4458f295cc2902b076b6b933e44ee0256fa9aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73746608dacdde3a012d687fdb644c5474d47c73127d5e1f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a73cc6e5e7e6ae759c4cfa2485abe30e95e7a36eb732a05b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefaaabd1ed2a9ee7d7d14099748244724dfc7c160ef7f67fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9f5a6418bfb61715ebac0183727c701489a863e02345c2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7e75ed5952fd5b97c320f827415b73f791a0b6613a8baa5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb857efd34c13b34e5d100901b3ec2d85baf8a6ebc2876c88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53601ea1b7c262a83e14dafa890dd3a22eee3758d4b763388;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2aaca8a78f5b08c5042602dcdc25815d33593effd2ea50875;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7aa8c41b431cb3bab745b3c47613e07149e1ada28b3d7ebd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8a8a8bfb39bb95948484d7a0e32f12710e250fcc5863b3e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe1e60913b993280e4d66f2216dc481c221e3b16879f66f38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50a716cffa99e784847af3565da2edb626928dbe40ac625b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6c7f668e6bdfd78da4b7ab6fc7411e59452f5487b3d4b202;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbbfaf930d31449deabf2001d8451b3490529c9e714f6aad7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9dd0ef3a4d83e39fca6baa583476ac32bb6f086a03eb6bac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha955aaa75e496a75e388917781e3c79dec119a9c3b0de5306;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63514dcf747ecb2d9151f8a9d37d04685afc0f80363943b57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b38ca2c28266bd8613cafe205476dfcfd1575edcd75e1b0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf05473c4e6e050f448257f4ded6e6b053b056f572adb07c88;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h986f970b03267f075c7a1a7c5120da2686fb6d36759dad16b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd4f133f9db4102fb0066a6460e550e9daa3d89c3183a2061;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a90ec83cc590fd98401396b5b7483f8e5716e08d984e2537;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h944405399a28e501d985f94704227e1712b670018361ba308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha28a73247bffee14da139602e6dce55ae0f69eeb35c21cdae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fa27792c55312ebce742436ea9f6d12f201b621fef49644b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f906284556aecf08cff8399a6245023ad68470c472e231c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac2af6f412a87819c23d0e90a5b234d0fe317aec8fcf17738;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1f4a8b2bab30785cf86f225b08f288f4aee91522e4140968;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bf84994b372fe55b5f813ac8b77eba8f7fb826a1b5bdb149;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b0ac242d0f2a7c2b34465f8a3bd76d4284a034cfe3e410db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb24e86db78cc9bcdc26b0a13d52eb123f5ea24a52b706d66;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6d5f1cb8c153c2b069691158a6d8b7949c4642b9534e4399;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70dad489d5e4eea7d5b311f297ae2449707ead143c26aac0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h230813c3b4a92a36b43064a2601387ac0fb9e4dc9ead1126b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5798f16cad7163bf12bede0bc18b6eab17479bb843ffc8f91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6647a114b14f4a6aa320a86b4327d14f863bb896890d4ac76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75990c133079ab38338f25fe99f5f38aa71bee5d231dca52d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h450d1629f5676a579b7bed887c72c4cc67a8b60e036008771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2850a30444b246b56537b80c7e1baf1e7de09b951311489b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55d983c22866439ec45ea8b50a9654e4a23256787be7e606e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d1a52d63944afafb9a17541442d1ec3e9bd0b1d399d39c81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2763b88f9f0ee1b15395c6b2f113785e8fb7910b57f233a85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefa273666739ef6d9745e66335fef7282146c9a60efafa6db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8969437668e41845a8dd2f7677f200436c5956b82da098612;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80e814491547abf8e4f5676d8fcd23946b5e904a090a8e995;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf68ae1ae8921ccce77b2d7939e72fc72d1f790f5455e7804;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff7a1412badf6f04a89d6d7210a1743c2633be40ce0774a99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h358b7c12557839dc857dc4e3abcce827473e4c70fbd2d74f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22f067f32d527eb711fa84da1351365ee3317c9b2537427de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d7900e4038bcf3ac5d269dc4ef3006223384ecc55c1b210b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac9bd3de81c23dbc51edfbe19ba232eec3a7f445a9953eb24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57274c9e7297c95855abfe98f6b405e1f3eee881b5255ae19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41f96183169c2f25c0efa2c38d8f2a46895f1ad38d1bce3e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h835af08b0fe276b8108f87181d70c5ad7cbabb288507759e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha086a732cbbe52c71ddaadf1de255c117775f5411fd9d0e6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he99a2bbf7fe563ce6f620754fff03d81a8bdc7144c15cb3ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44cd83c8fea2ff03bedea0782175dfad1c697407faa237300;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha17e2300c425dc74b0a2118c6c1e52604ab9c4dc9371db5de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65230711599721536a673b1c6caa50a0f663757fa048b41cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he14435f3e7b5b6dff8e3dc4618c9cd44c3bff06462f7dde1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5adb2da4259ee2fd175bce46aba45dc18f76b6f878928de8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bc2de17bb0d7c4584e3391d8a0b729c46d669a20103b2c06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd782308eb1c6c367a374902de37a39c14a7def64e0b08e1b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c712729dd48a025b9246a46744f3692ddc03762f5dba132;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53a7442c53b94cacb3856e32dd10bca631854b14794b406d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14816264507b3e223167ddbdb266559d1ff65877c1f2f4ee6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd28eeaf6ab098170c91f6f5cb68643419d8b0815ea7e79290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5526ef041c025953bca376390eec579944163d3d1b595e7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84ec84bbbc6a6706a9d3f4d1bcef66c76a11a13060dbd3965;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56280d9f63852f7002d9b4d05d5793f05f145345f0caa9c7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87a045d90fa4eff34ef4fd5a5ff1c49e819a79af6cca9d73e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea85834dec68b6fb9755d889a201fedf938ce68927343b94b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cfff1ce4fabc60c5c9b58336bd4ef3ff6f72789bb5a2b872;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5271c4c4ed58281799acb320c35b256efbfba6b1ee8e7b6d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47433ebb369b84f296c97b69af41a5ead1d200a3f9c7ef1bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heafefa2c0c039348ac1c761ec982f2b4242879a556c1c05ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d0918d4af48f93f31202125e9db18bff53553ed0db0f775;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e37783757b19d3c046562a3f172bfd4beb12138de6367188;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35404a225b87ae33d764df753fdb49f6fd16b1ed110b6c276;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f03d50c2c174966f38b34fe6da5e276c5f3b1bdc5a55d08e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85ae0c377cffb7838788bf8a47df0658172981f84158aa2f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58fa1e8f2cbe8cbf19e24911ec6775378f7bd447e81e86457;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h654eb07dcd54113f938b63e2a58a85b05e1f4fc366742f79f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9c6756cb789c8841c0f62b855a543d66fe161e89159322b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebd59e575c31846f6c39a165d35bd5eee3ea178567b685d2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1222eb25e1964fe7e4698d8e302e97ccceb2312fafae050ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83b4bcfab8aa69f9cd6f1020b8d8834cee51f8599af266a27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17e9f2c63cccca2c124ee05973959ba2ddecb9d740cf33051;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49f0ab26dd900f9410fab78bcbbd4492f8eb990b7244b0694;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87f210122d56645d9ea68836ee107a20724f77025ae892878;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e87d114a018fa0c2c8ca9000214e5fe2969f770f4f95ec94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89af8c4aef22eb1c3a9143186e9b6198bbd1c0df53bd4224e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7af0cf2350c48e7ce8a379c796ac00df3c41819bf372c3af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1100bac231cfadd2e58f2a63c536792e734674879c48c6920;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fc04459b0c143ce98d25a7684c9646d9b8bc57c61f5706f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbbcd2fe6b81bf8360a435fe57c2808c6406ab236eae604c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h246b23cd7bd3710c341bbcc509c74ab52b347c73d3dcaab9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6af29ba84ce23b12e568eceb1338ef4fea8f98a82762a31af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ac69a467c24412b8d4b9f919ff519c633cfe01377375a9ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44e5b2a6bab6705dae2cd47b3069cbbcb1a180381e175b119;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he57e0b006190140bae5260ec37056e7cd4a87cfc548fa705d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea87fdf82ca2ebb78f8e8166b350309346200d0f7b95acc5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b0240403553cd4c67e7b2e3aa4279e9c7ad560b4e60ff50b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h829284ec67483b17e28c3494fff2acd8427141125a0a138ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4219f049ea91c84c55630969a6532a20ebfdafcba2fb367eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb236a29e79571e388444a36ce39b282ae54f5912cda92ff12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d30939551c4b3d9f9260dc093f8e14b7b7fe2a6bef4db75b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f2558a50056fef201ad53f405c34482b3c81ceac05dea106;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd16b3ef0aee65740bad13fce8dcf75ed496305c6dfbbc3bdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefbf7b89211474f9abec7757a46ca1dffc874e61a420f0b65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26aeeef32b43635d4408474a57d2f66ff36a630ff4b6cc6f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd363c2b3437ad711ff20a16a1d5a8422073880621c8a293c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39c9990572c21cf41f2c62f6c8a2295a2a7f13e6833476634;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb11bd261ffa93142f07639af1043f4c2e8498c4bb263c4178;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f62855f290ffb87fe56bc0f0a7f80a3e2edf0c6df4d891c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h925b48637ebae54004e603b9a98574f23f3f10a17f76228f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54594262a564feb74328e0b5ebfd5917d8bfc70f2bf53bf2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd725515203b91c93811a3419d9ef6a6ac355b566f825a49d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc07e32a3aadcfb4801a865d7fe3fe56f86acfb345ad513eb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94e5ddedfb3eaa5c5e92b7aac59fe02b0631bc607d2aa7689;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h519e0b0cf7dc6e8599faef8770ebec0295525c1ff1f756d8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ee8745180a4b48a677c1bb9fe3669028167153d82247143;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6507af0afa6438ba8e4b1ebeae96c80c7b78d34851632387;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eb526b573cedc1d3f5c2927819ed26fefe438972423cc5cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5acc112792f5f52f1b91daff9868b1aa7c5662fe315657498;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69f4fe0350f5bafb19d1c47572ca6c2f8ea657f7fa70d1c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb96777801e75850825398ed239452cda32c3165c2e5c88773;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h629985b79a3eb0123eab649e18ea046c00a0ffced2deeebed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbffb00e079c8a1d12532ae93f6459dfff19edada5d67f8411;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39ebe1e3f4dd246b0d069a74363e8b999e9b28574cf6ecca4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37873502a593af4136ca16ebdfcc4f454fb087e6a12c27504;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6596540ecdfd149f913906a9de50c9f7f567e84957ae20713;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60b9344c94cccf2d0e674bc6040d35229f8a4a230ad72e24e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6cbf1a10f50ea79a24344a0378173441987948c389d2b44a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58c53eaec4b865d13b7a9a810a995970b8aa83a1c6043ea36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75f917b63f7fc3eeb806cd91350254cf3ed7f16bb4b683835;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h963aa5a936c58cdbd8bb8d2e7367405c3a86d4b83a9336813;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h959104a3064f2e7cf54b323ab88c391c19181bed5f2229779;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b30d5114ed6c2ade790b02620aa90e2c12d5c4c52650e9dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h802788da658d9882506831b5aeb2b0167b35c5a38dbe8cd77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h170909b1cc2b34b42412a77ab0f497ded088106d2d1e33d15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefe25b1a724e5953e9986a9b2ad4f7ed30fe4abec836dba14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45ef7d075174a21a8133414c030c85565ca9bb423b4488a25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7216facff4281ce4abc6a3e5e161e93a0b33bb3e9e8085d29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4eb1324794a69035954a7f0ada3481ffea80d70a57344832c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9574d5e58a1e479736fb5900c0c0ac78851ae912754c14973;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47860840f8cfc93cbac78e8c01b9c473815a6be3391c3cdbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3aefb147de81970752ae2a544a653295f59c493fa685ecb28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57411f0ee86f953e93625f5e7235b37ac0822b08862d5817f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5e632b9e9affd4641df4e94bbcca6bb05ce239d980067f72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0a6aed0249afbf6f8a177d3484695eb56d694eea605deeb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a6827052cea3ce5d70533e34c33a8baaa5e80c56dbad69d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14e279d62fe48cce7dd416e4ab678559fd8ee4e3a151404ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h275949333b4e2e30e931f8324765c1c5d792192fd82028746;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82c876c7da1b313239e6f7b046f752aa6de92c5412fa5bf25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc73060b023794ef07ddec48f54741e9fab7232edea19c3748;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbbdaaa9ae2c602a767f0d0d2a3502beaa114cbf8fd54fe7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h524dee3751399427f8f9887c37ef55d4b05bb5b4caceddb9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ef9178623426b2f2e960cab4e8c742a39b4ff2e1b129c58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b0d5e66cfcd8bbb005a4df88ce04539c9ef4747441647182;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36934a5e7674b35360fe8d32cfe55df453910010aac8a8214;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce2414c9c3941cb2cf1cfe9f0c837c5b0715fe30f9632c8b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fbcf31a132032d398671e0399be32770c3d473041689bd21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h300e0c768f02ef437ec566ea8c8b01426a17d235e1ed4f1e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc067800b36f4a4e78aeed0a69fbb516f604389b4b8ebfb1ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha70169339eb55f27bc05ae5501b5444576f0976e0a7e83fcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h494eaaa5d6aa1703457e614ad0cdcf136b390b801b7957a8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbef673cc13003f481ea50fe629222ee8ada929e1b387bcfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1910d61eed0384c5556f461c951c55a2b5ffd3dbe6fe7d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1792fa6b48ef23d4d8d8c40ca41bb45b13a727df7c7ac800;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2846ec25df1fedc2a2fdcc0cdd264e52529d41def61c5a501;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed9784144480e660e446a6772ea44e60703be5bcc61345144;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h375af6a47021319b176cddcc63b09e86ae6475e258edf8c27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdaac54069f2095de3aed11cb6a0e9b788a10cc416a8e0a0f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ef3f233b808777f5306b6b4043b1dc545f2a28e9cbdff143;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5958f40043626626c20aa10ea5b7b8b779854af4f8ab014e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he99ef515d08d41d53f93a2f9cf23c2163165cd8da1855791;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b98aa55f1b71ad8ccd1e55c7ca15074e427c98e3bae4c8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c808787e25bfad0680ad11fa52d4c39e756c29c6491d707b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56bab3ac886f577fd28ff987464ea99df975c103e53dc39f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he90fe1a4ae74fb252459eff3b8e54fce3b9081fbb4ffadeb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26b73faf25fdb3b6fa8d435681db65f886cfa08a241e599e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae24823b68f285c440f68a66c48bd3312a350ffe0eaf8f07c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed65c91664aae1c3057589960de624c9d81f830e7894c1661;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c883c3120a9834140c304b9f6307177a3ee0e22ebb6ee0d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2add0dcc949c3b932aa34ea4b93379f0e0d9eece7c648f17d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7bac0cd8baeefd3519bb2e053f6445288cd755d3ffa44be7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2793578423aadfa68e45962e3f600bb3fbfffb4a9990baba6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h895d2b0d32cac985290d56dca5a527453429bb82e564f4490;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9d2b6b8eba9f21b70aedb6194810a250620e925d1a65d927;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee7d53a586e7ac166f990d90d0db4452237aa7f5c457b3387;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f2c137db9ee260fb3db0a36d86f062647060034db8cf562d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ea83439fbaa05de723f39e9cf144ef25400dcbdfc3983099;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h973db0d7de8524bb018f5877f52fd18051bd2b4aabb7bfb48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23b699da8014f38e14ffd441c478aef8772940f63b016b71f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf05cb08d7edf4798bc2aff9287b5491900ca2631f821696b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac05a0e5e3f095d4a5d563a8b0122b46acf9bcf26479394bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4873cb86cbbd140ff0c722f1555e44258ceeacc26d78b1db8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40aff1c1b890095d5bc2eb522334e70518dd8488a425fbe4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4fe05d1620235ce8cce4bf32baf9288aa6928b24cc5d9f7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6fe79042d43b85f61646f23e918fc9fdb8e7ce9401ed1b4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7837786910ed65bb82f191b855a81c3619a502342ae407dd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57f7eed80691df3295da540a5cb7bd0fb123901394cac01f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1947e96ce4778615da79f4e7662b12ab476eb6e6b173e6c4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed041bd1305da99289bff20796dedc05cb3fff218d007a93a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf47e4cd5ceb5e3293e9e9b43ebb7b4a870cdeefdb8a4acf04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1361abc4633e5c50a3518aa9d16430d27c11a7614a1cb683b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44d4400987ea228cc2904a105e7e182941b75997ca328ad46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f294027880dce22feb92859180ab0dcf1660981179199c75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h304c77f47d5f4f5754d84a59698e67034bcdd2526c25f7471;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a3b9c437a78aceea1a9152f58633b611ca2cf93c38810ccb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h586a30ce45231dbd63fa0e82990a413e470311096cfb1baa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70e981364719e68e4837c91d69fdaeaeb0479316de575c748;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fdfe5b4e20f7431bc96283556506eed8db4b1986dee613fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42b7ca14a05abeb10bc6495db4e81aa3ef6915bc70cb44d6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17df501fa9d8c4a47b316bc2f77b36db95226f0cb68c95789;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8687ec79a01cbbe2ec5369b7d1b492cfd05936c1e221d5d31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5d93054e78f12957202746a2134527e523aba73026229281;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h310182c6a45243975433aa2c45aa0635cfb30bff0533f36cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf40a086b0864f65a1e914f3351e830857d509e6f9ddc05c3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15c24acba3e6219a0045e1a2c1d6ddae0b7da03312955fd6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf13319f25efc079d7f70f52dd96390ca2ad90b6b5270abf7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22174e5271e93b15a13da084e71836a3997f78f8584b2fd44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5a6b89cddd69a2abcfa84ff02a14abeff2e08147582eedef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h385d801dda302687c1ed878ec4bd6fd2cdb79d22812f736fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e6fff931947db7140775f5a5596f1648f7030113e9d63fc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbaea828c91ee4b539013dd61d0ec13854a99c50981079b9d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda8be7d7cf8994db910b57fd19b9796ca09a4e2134a6b1266;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd6e5a9be6434827b13127a7874f74d7670b3a0ef1beb2265;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h296456f03c2a54c76f19e775c7ec4fde408509ccca12d33df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32840b26d0b691af9f321cbe0d6931cf06de774a85b7ee66c;
        #1
        $finish();
    end
endmodule
