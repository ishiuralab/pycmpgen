module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [7:0] stage1_0;
   wire [12:0] stage1_1;
   wire [16:0] stage1_2;
   wire [17:0] stage1_3;
   wire [10:0] stage1_4;
   wire [5:0] stage1_5;
   wire [0:0] stage1_6;
   wire [0:0] stage1_7;
   wire [4:0] stage2_0;
   wire [6:0] stage2_1;
   wire [8:0] stage2_2;
   wire [7:0] stage2_3;
   wire [6:0] stage2_4;
   wire [9:0] stage2_5;
   wire [8:0] stage2_6;
   wire [6:0] stage2_7;
   wire [4:0] stage2_8;
   wire [0:0] stage3_0;
   wire [1:0] stage3_1;
   wire [3:0] stage3_2;
   wire [4:0] stage3_3;
   wire [2:0] stage3_4;
   wire [3:0] stage3_5;
   wire [3:0] stage3_6;
   wire [3:0] stage3_7;
   wire [2:0] stage3_8;
   wire [0:0] stage4_0;
   wire [1:0] stage4_1;
   wire [0:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc215_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3]},
      {stage0_2[1], stage0_2[2]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc3_2 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12]},
      {stage1_1[2],stage1_0[2]}
   );
   gpc7_3 gpc3 (
      {stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage1_2[2],stage1_1[3],stage1_0[3]}
   );
   gpc7_3 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage1_2[3],stage1_1[4],stage1_0[4]}
   );
   gpc7_3 gpc5 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], 1'b0, 1'b0},
      {stage1_2[4],stage1_1[5],stage1_0[5]}
   );
   gpc7_3 gpc6 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_2[5],stage1_1[6],stage1_0[6]}
   );
   gpc7_3 gpc7 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_2[6],stage1_1[7],stage1_0[7]}
   );
   gpc7_3 gpc8 (
      {stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10]},
      {stage1_3[2],stage1_2[7],stage1_1[8]}
   );
   gpc7_3 gpc9 (
      {stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage1_3[3],stage1_2[8],stage1_1[9]}
   );
   gpc7_3 gpc10 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage1_3[4],stage1_2[9],stage1_1[10]}
   );
   gpc7_3 gpc11 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage1_3[5],stage1_2[10],stage1_1[11]}
   );
   gpc7_3 gpc12 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_3[6],stage1_2[11],stage1_1[12]}
   );
   gpc7_3 gpc13 (
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9]},
      {stage1_4[0],stage1_3[7],stage1_2[12]}
   );
   gpc7_3 gpc14 (
      {stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[1],stage1_3[8],stage1_2[13]}
   );
   gpc7_3 gpc15 (
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[2],stage1_3[9],stage1_2[14]}
   );
   gpc7_3 gpc16 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[3],stage1_3[10],stage1_2[15]}
   );
   gpc7_3 gpc17 (
      {stage0_2[31], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_4[4],stage1_3[11],stage1_2[16]}
   );
   gpc606_5 gpc18 (
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_7[0],stage1_6[0],stage1_5[0],stage1_4[5],stage1_3[12]}
   );
   gpc7_3 gpc19 (
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[6],stage1_3[13]}
   );
   gpc7_3 gpc20 (
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[2],stage1_4[7],stage1_3[14]}
   );
   gpc7_3 gpc21 (
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[8],stage1_3[15]}
   );
   gpc7_3 gpc22 (
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], 1'b0, 1'b0},
      {stage1_5[4],stage1_4[9],stage1_3[16]}
   );
   gpc7_3 gpc23 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_5[5],stage1_4[10],stage1_3[17]}
   );
   gpc15_3 gpc24 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0]},
      {stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc215_4 gpc25 (
      {stage1_0[5], stage1_0[6], stage1_0[7], 1'b0, 1'b0},
      {stage1_1[1]},
      {stage1_2[0], stage1_2[1]},
      {stage2_3[0],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc3_2 gpc26 (
      {1'b0, 1'b0, 1'b0},
      {stage2_1[2],stage2_0[2]}
   );
   gpc7_3 gpc27 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_2[2],stage2_1[3],stage2_0[3]}
   );
   gpc7_3 gpc28 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_2[3],stage2_1[4],stage2_0[4]}
   );
   gpc7_3 gpc29 (
      {stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage2_3[1],stage2_2[4],stage2_1[5]}
   );
   gpc7_3 gpc30 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], 1'b0, 1'b0, 1'b0},
      {stage2_3[2],stage2_2[5],stage2_1[6]}
   );
   gpc7_3 gpc31 (
      {stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[0],stage2_3[3],stage2_2[6]}
   );
   gpc7_3 gpc32 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[1],stage2_3[4],stage2_2[7]}
   );
   gpc7_3 gpc33 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[2],stage2_3[5]}
   );
   gpc7_3 gpc34 (
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[1],stage2_4[3],stage2_3[6]}
   );
   gpc7_3 gpc35 (
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], 1'b0, 1'b0, 1'b0},
      {stage2_5[2],stage2_4[4],stage2_3[7]}
   );
   gpc7_3 gpc36 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage2_6[0],stage2_5[3],stage2_4[5]}
   );
   gpc7_3 gpc37 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], 1'b0, 1'b0, 1'b0},
      {stage2_6[1],stage2_5[4],stage2_4[6]}
   );
   gpc1406_5 gpc38 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage2_8[0],stage2_7[0],stage2_6[2],stage2_5[5]}
   );
   gpc207_4 gpc39 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {1'b0, 1'b0},
      {stage2_8[1],stage2_7[1],stage2_6[3],stage2_5[6]}
   );
   gpc215_4 gpc40 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage1_6[0]},
      {1'b0, 1'b0},
      {stage2_8[2],stage2_7[2],stage2_6[4],stage2_5[7]}
   );
   gpc615_5 gpc41 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {1'b0},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_8[3],stage2_7[3],stage2_6[5],stage2_5[8]}
   );
   gpc7_3 gpc42 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_7[4],stage2_6[6],stage2_5[9]}
   );
   gpc215_4 gpc43 (
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {1'b0},
      {1'b0, 1'b0},
      {stage2_8[4],stage2_7[5],stage2_6[7]}
   );
   gpc3_2 gpc44 (
      {1'b0, 1'b0, 1'b0},
      {stage2_7[6],stage2_6[8]}
   );
   gpc1_1 gpc45 (
      {stage1_2[16]},
      {stage2_2[8]}
   );
   gpc135_4 gpc46 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc7_3 gpc47 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], 1'b0, 1'b0, 1'b0},
      {stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc7_3 gpc48 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage3_4[0],stage3_3[2],stage3_2[2]}
   );
   gpc7_3 gpc49 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[1],stage3_3[3]}
   );
   gpc7_3 gpc50 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage3_6[0],stage3_5[1],stage3_4[2]}
   );
   gpc23_3 gpc51 (
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0], stage2_6[1]},
      {stage3_7[0],stage3_6[1],stage3_5[2]}
   );
   gpc7_3 gpc52 (
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9]},
      {stage3_7[1],stage3_6[2],stage3_5[3]}
   );
   gpc7_3 gpc53 (
      {stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage3_8[0],stage3_7[2],stage3_6[3]}
   );
   gpc207_4 gpc54 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {1'b0, 1'b0},
      {stage3_8[1],stage3_7[3]}
   );
   gpc135_4 gpc55 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4]},
      {1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage3_8[2]}
   );
   gpc1_1 gpc56 (
      {stage2_2[8]},
      {stage3_2[3]}
   );
   gpc1_1 gpc57 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc615_5 gpc58 (
      {stage3_0[0], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], 1'b0, 1'b0},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc135_4 gpc59 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1]}
   );
   gpc1343_5 gpc60 (
      {stage3_5[1], stage3_5[2], stage3_5[3]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1325_5 gpc61 (
      {stage3_7[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_8[1], stage3_8[2]},
      {1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage4_8[1],stage4_7[1]}
   );
   gpc1_1 gpc62 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
endmodule
module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    wire [0:0] dst0;
    wire [1:0] dst1;
    wire [0:0] dst2;
    wire [1:0] dst3;
    wire [1:0] dst4;
    wire [1:0] dst5;
    wire [1:0] dst6;
    wire [1:0] dst7;
    wire [1:0] dst8;
    wire [8:0] srcsum;
    wire [8:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0] + dst1[1])<<1) + ((dst2[0])<<2) + ((dst3[0] + dst3[1])<<3) + ((dst4[0] + dst4[1])<<4) + ((dst5[0] + dst5[1])<<5) + ((dst6[0] + dst6[1])<<6) + ((dst7[0] + dst7[1])<<7) + ((dst8[0] + dst8[1])<<8);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src3, src2, src1, src0} <= 128'h0;
        #1
        {src3, src2, src1, src0} <= 128'hffffffffffffffffffffffffffffffff;
        #1
        {src3, src2, src1, src0} <= 128'hdeb71b5e1075b0571d50e2524e540702;
        #1
        {src3, src2, src1, src0} <= 128'hff6968d7fa5c5bc0686e5a4fcfcf36a3;
        #1
        {src3, src2, src1, src0} <= 128'h58233f3b7a6fbbb7fe740fad91805cff;
        #1
        {src3, src2, src1, src0} <= 128'h8abea763ff53187965f0fbd0ee042710;
        #1
        {src3, src2, src1, src0} <= 128'h95a5bb3f2c9898783ddce887837eaad6;
        #1
        {src3, src2, src1, src0} <= 128'h758e9daabdffb6edf0edb1b677f8458e;
        #1
        {src3, src2, src1, src0} <= 128'h9d31f08e793fd2c362479abced637639;
        #1
        {src3, src2, src1, src0} <= 128'h66c80c0e088abe389fb7b0c37f1268b6;
        #1
        {src3, src2, src1, src0} <= 128'ha542e71cbe352a0a3a51eec901493f53;
        #1
        {src3, src2, src1, src0} <= 128'h86d946692f995b36ac9eabc430a71628;
        #1
        {src3, src2, src1, src0} <= 128'h2b3f13fe8c7cf41b39913e39aec9e05b;
        #1
        {src3, src2, src1, src0} <= 128'h3c6ff23fca913844b216486be8dc715f;
        #1
        {src3, src2, src1, src0} <= 128'h8d9c8f4c98db9b556b36351c67b4650e;
        #1
        {src3, src2, src1, src0} <= 128'hde883fc4557ae951c16d856ea0ae335f;
        #1
        {src3, src2, src1, src0} <= 128'he53bb0f4f8b1b0672523518913461b5b;
        #1
        {src3, src2, src1, src0} <= 128'h664ed218f3b66ce23a20ef1782a60efb;
        #1
        {src3, src2, src1, src0} <= 128'hedf8d1cc5d8a4400f08241b0faa229ea;
        #1
        {src3, src2, src1, src0} <= 128'h732e20f4112fc5edc77713824cf77237;
        #1
        {src3, src2, src1, src0} <= 128'h5bf7bd54c9405478101e8641ef8360d9;
        #1
        {src3, src2, src1, src0} <= 128'h77becce62e2ecd7be365fdadefc1f61c;
        #1
        {src3, src2, src1, src0} <= 128'h28187e5cb74cc6f9cc14c5142455e5e2;
        #1
        {src3, src2, src1, src0} <= 128'hcddad66240d8c589022d1bcb7a0d04f5;
        #1
        {src3, src2, src1, src0} <= 128'h731c656842c055a2c5909884b8ff6836;
        #1
        {src3, src2, src1, src0} <= 128'h69fae163581385a4cdacc8274e7896ca;
        #1
        {src3, src2, src1, src0} <= 128'h46bf6be9366b915f8ba46e3d762f6363;
        #1
        {src3, src2, src1, src0} <= 128'h1cc5c35df965b67d3ca370ec1ded61b3;
        #1
        {src3, src2, src1, src0} <= 128'haa150be8b5f73d8f599064a683a01527;
        #1
        {src3, src2, src1, src0} <= 128'h131d71ce80ab84e08e575bb544e59be;
        #1
        {src3, src2, src1, src0} <= 128'h3e2fdb3e2d8e30941898b6a28b4621aa;
        #1
        {src3, src2, src1, src0} <= 128'ha63b497ead28fb87d07b990272c0e593;
        #1
        {src3, src2, src1, src0} <= 128'ha50fd97499ff319483c849ed6d8d8f35;
        #1
        {src3, src2, src1, src0} <= 128'h84dd1baf9941a37264915865b498cba5;
        #1
        {src3, src2, src1, src0} <= 128'h57b9f1262db93903b038fbbafb49f924;
        #1
        {src3, src2, src1, src0} <= 128'h7f3627f0ea76f2592a3a3a4368e586dd;
        #1
        {src3, src2, src1, src0} <= 128'h32d72ae0f450f7327ff7993d6c16c49f;
        #1
        {src3, src2, src1, src0} <= 128'h410be4c27edc37484943448e9dd6c5f1;
        #1
        {src3, src2, src1, src0} <= 128'ha5972d187e0e64e8f0836cc557e38c5c;
        #1
        {src3, src2, src1, src0} <= 128'h3f8286c295031fbce0c66527aa47f766;
        #1
        {src3, src2, src1, src0} <= 128'haf981f0ca7f1aa22031493264806c7d4;
        #1
        {src3, src2, src1, src0} <= 128'ha00ff21134c53fb9d37fb672652f290;
        #1
        {src3, src2, src1, src0} <= 128'hdee94179f129d89a83967c7b657d233c;
        #1
        {src3, src2, src1, src0} <= 128'hf9515ef115ea9c2fabf5c3a7c1075cc8;
        #1
        {src3, src2, src1, src0} <= 128'h5d74711fe96df4723292b2747575db0d;
        #1
        {src3, src2, src1, src0} <= 128'h2b28913c9ce8e9bd946ecfb317ffc9d9;
        #1
        {src3, src2, src1, src0} <= 128'hde9d16ceb1932caaf925043a1bd80492;
        #1
        {src3, src2, src1, src0} <= 128'h80cad31b146e5b29c5ff2bcc9214d4;
        #1
        {src3, src2, src1, src0} <= 128'h435ff98f00972d3ae3bc1284554a2407;
        #1
        {src3, src2, src1, src0} <= 128'hc94f3a4d6ddc5125bf61cdca6aa94e6;
        #1
        {src3, src2, src1, src0} <= 128'hfc8b849c07e252c379f29167c7c93693;
        #1
        {src3, src2, src1, src0} <= 128'ha8582c427b1e4635fed655e18184f3e4;
        #1
        {src3, src2, src1, src0} <= 128'hd29c70425740c3facbba12ec20d42285;
        #1
        {src3, src2, src1, src0} <= 128'h95f81d190757d901961994feaa504e19;
        #1
        {src3, src2, src1, src0} <= 128'h6e1d17b1a3382194de15b88681b6ba6;
        #1
        {src3, src2, src1, src0} <= 128'hdc2a5ab4cc8bf0bdd8924b9a1c09decc;
        #1
        {src3, src2, src1, src0} <= 128'h6ee10d4d9613bbcfabcadb25aadbceb8;
        #1
        {src3, src2, src1, src0} <= 128'hf3b3107578f036bb7be4a923ac02b23;
        #1
        {src3, src2, src1, src0} <= 128'h3d2119a7e74524714f1c58bc40f3e4e9;
        #1
        {src3, src2, src1, src0} <= 128'h4741e1af9ac00f86d76d77b363a44864;
        #1
        {src3, src2, src1, src0} <= 128'h7bdbefb5ea9b0734a9fb371189135235;
        #1
        {src3, src2, src1, src0} <= 128'h119ce5a4b942e84068048958fa2390ba;
        #1
        {src3, src2, src1, src0} <= 128'ha3b26aa6b0998a87c20f29c125887436;
        #1
        {src3, src2, src1, src0} <= 128'h6c467e797a80db83c4b63aec2751114e;
        #1
        {src3, src2, src1, src0} <= 128'h252fa79f2ce52c6d30bb223ce8fcf060;
        #1
        {src3, src2, src1, src0} <= 128'h419c5e32cb4b65a3e881a9d9cdc2adea;
        #1
        {src3, src2, src1, src0} <= 128'h12de67cb3525c2fc0819ab7946c0150a;
        #1
        {src3, src2, src1, src0} <= 128'h518603d3c6dd0f05e19cb2dc64aedf6;
        #1
        {src3, src2, src1, src0} <= 128'h49d5279ca3d2aa2fe1f522d0a27d0002;
        #1
        {src3, src2, src1, src0} <= 128'h15bf8f1129848818d73e7e4dc1b7a444;
        #1
        {src3, src2, src1, src0} <= 128'h44ee549453f35683c08e31ee63b425ab;
        #1
        {src3, src2, src1, src0} <= 128'h5e211b558ae0aaa3511747b6542b8e2f;
        #1
        {src3, src2, src1, src0} <= 128'hf910083802b6cdd8814d103f652d5ecd;
        #1
        {src3, src2, src1, src0} <= 128'h7c2b2d798c05c088f3e65447e51d5722;
        #1
        {src3, src2, src1, src0} <= 128'h11be3ee0484a56e44994ae1b67ff192c;
        #1
        {src3, src2, src1, src0} <= 128'h7ad3bb26b1115933057efcf5ff6da932;
        #1
        {src3, src2, src1, src0} <= 128'hfd24399a85e529678a31d93816f87d03;
        #1
        {src3, src2, src1, src0} <= 128'h56694b10bbb24861f75c96734d36997;
        #1
        {src3, src2, src1, src0} <= 128'h1cc8ddfb1dcd140d2eb945316a3d32ed;
        #1
        {src3, src2, src1, src0} <= 128'h282917277e39683c2df75a93d7ad353d;
        #1
        {src3, src2, src1, src0} <= 128'hb736bdcfff71d4def047372f8241a3d7;
        #1
        {src3, src2, src1, src0} <= 128'h1aef56dc3a506668925bfc7f34804fb3;
        #1
        {src3, src2, src1, src0} <= 128'h8038649c21aae075f1452c9d9bc57ada;
        #1
        {src3, src2, src1, src0} <= 128'h31fce3b10c18c01189bcd8bc8103568d;
        #1
        {src3, src2, src1, src0} <= 128'hc98a39bbcd3776d78307e749f17c94b8;
        #1
        {src3, src2, src1, src0} <= 128'hbe2c4905ade0db8ca675454a11c18f4e;
        #1
        {src3, src2, src1, src0} <= 128'h8611dc01ea78576cdf304d957c27674d;
        #1
        {src3, src2, src1, src0} <= 128'hb53ed1ea0f27d1d25b786d9dab2598f;
        #1
        {src3, src2, src1, src0} <= 128'hfee2ed04b6adb49ea5766c94c4b1bf5a;
        #1
        {src3, src2, src1, src0} <= 128'h5d97417e360f2e2a48fe8ad0b319260d;
        #1
        {src3, src2, src1, src0} <= 128'he729fe353042be009f59c59b79766a7e;
        #1
        {src3, src2, src1, src0} <= 128'h4252595ec5b8d08bc4c96ec34bef4819;
        #1
        {src3, src2, src1, src0} <= 128'hd029627f02d8b1de26b0af7e470c727;
        #1
        {src3, src2, src1, src0} <= 128'h41c1e8cc96e747bb5b0867f434b96c8e;
        #1
        {src3, src2, src1, src0} <= 128'hf83d10a0a7066ba5675861e45e3dbfe3;
        #1
        {src3, src2, src1, src0} <= 128'h94b5cfa4d4f9b3a6b9c96ae1d748448a;
        #1
        {src3, src2, src1, src0} <= 128'hab8bb83a46ca974c206e7896d88d0138;
        #1
        {src3, src2, src1, src0} <= 128'hf27a60f2782da956198216a6842fd26f;
        #1
        {src3, src2, src1, src0} <= 128'h4828ba5b6f7acc620ea56f8274e398bd;
        #1
        {src3, src2, src1, src0} <= 128'h48a8d34776574f9af6786b2118e8457c;
        #1
        {src3, src2, src1, src0} <= 128'h5ba8a5fc9eb8f285fca795557f1cbc5d;
        #1
        {src3, src2, src1, src0} <= 128'h17e054acfcb2cd269a6aa9105dc3394c;
        #1
        $finish();
    end
endmodule
