module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [17:0] src19;
    reg [16:0] src20;
    reg [15:0] src21;
    reg [14:0] src22;
    reg [13:0] src23;
    reg [12:0] src24;
    reg [11:0] src25;
    reg [10:0] src26;
    reg [9:0] src27;
    reg [8:0] src28;
    reg [7:0] src29;
    reg [6:0] src30;
    reg [5:0] src31;
    reg [4:0] src32;
    reg [3:0] src33;
    reg [2:0] src34;
    reg [1:0] src35;
    reg [0:0] src36;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3])<<33) + ((src34[0] + src34[1] + src34[2])<<34) + ((src35[0] + src35[1])<<35) + ((src36[0])<<36);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd519fe898f0c059b2b5aec1a9ca3fca85ff3efa0dad30cb4cf0a06778be6880697a79ea5b03c0509f77dabed97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1542dd537cb6f6a655585f9f65742755d14da0137e3cefb0925ff34c359aa9a8cfd754a036e2ffde43835afb473;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188224b3d4e37d48432c8a7ae1c7da8c3de630183035fca199b78b9aeb946c21ad8e50e8e50ddf32d887ee2dca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136d501415a9ddda2c8dc22c6fc87e018a7fc0df1285dad26e0f32156233cb7dabc0678821385514797b0cefb73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h629d950323a529beb6faf64f70dfbde2346f557744e4ff156266f2ba2e196f542273ea16ffced5ba3a797da940;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd4c3158d90c56d2615dea6428291c251f2e1d23387a9ba79979f0ad90f3589170858868361f0fd51068b399cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haea42a5cdcb5e1507ac65fbde63611c4b1b284c55713dcf9a5005b83c2d1905e297128bf2406eb8a9c6779b9f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccadb519313a75b3bf1eb710cb9bdefcec5e14750223742dc4e4c4b335528a6ce83d2525eb69df5456b38028d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3c1f76ac8f111b9b72c6f2d26635d717150ef297638168b13e9fe7c31c9fa4e9e9a9646445c5dc8343feafa28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146c321b3d09860388a5f11c3b29fc014c169219eef4d90ee3f2302508dfae0c5b2aa84912a56f4497013cd06c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f99aa225947c4f4819affece69e097a2cbdcb4e25284e166399b67e62c393b965017b1bc28692ef847d61e0466;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114cd4a17329f33656c9982cb19f0b18762551069e383a5ab823b6c3f2c57f31d9dc07e1ba45d855aeabe667660;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77d3ee6f1dc1340db80b6a609d2fde322085c4139642d668461618fc4ff9396f69a76c7db76bdd61437f5ee57c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122c53fb50497068969d93b22817855f5fe09d0ed12d75057abb209d9111475bbe9601a780b7dbe688237d4dd0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1499bab59d01199d31586a0d05a8f9f56b232301516680a9153a0ea40f1c0e0abcbe544f943e3b13e3dc3355c33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1839b427868ccc11ccece3b0715ac75bb6ef19d1748eeb7f839f3cca6344862d3607618064761de4102f870c9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ae7aa296dcf94e3e1b1b8a2e7034c90d1620946dbb74b35c01642833d0f6acedbbe0bac5596d9dacb545b3bf0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ead3641d6a5ce9a03ee57c3a7921d32a3460ec495e3b5fd006fc5da226f518ff6add1e8a7f75127aaa46f06d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha39916ccbccbc867af2418358a84ed5d8566ac3dc960a9603c6d8c3ec37bea5f720af025d58816b2760bc7bf42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0b5b07620adf5e0997bf66ac267d029fb5e619aaee2e04562432dbfeffc887c50d35e84eebca8b2a7f070da67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbeea92a65b32539660ee3bc306c16df26005b981a6033a6c393f340b08c3db4aff3924016b1da2e609b209e812;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68489e3224a4e92976824bc6f68cf7058bfa2cf5a045d5f0941bc493b66c5732b8d0e6366da9e4c4717559cc86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1708163f0a9fa5830ca0edf1969decca3080d2e6b2562f176b6a94084c002ec3711ef4fdc4e9cb46fdbb76b18e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66fc15730938a117843ed7e64127747bfbdb9fa5360ff7375f419102b8577f265eaece02e44b66d0d5421cb075;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddac78b87e428b009abfff313d9b65963f64b2f38d29a7c82a3a12d807334a3f6eab887efc8a66422909a91d70;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h809cef5e004ff79675df57f63c7152fd06e56ec0ae73d49fdec177fa96aaafb0eb92b2cee1ab843c4acb9a364d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4f0b9082b4aae11f5e453f107d2a5600403c2726b961ea972c493f388656e527676a973f95e69fc425a8f828e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaca372c716ae0b05b09349de47829ca609f123a7fe724f9064b6ae85490ec6a143a966d9413061a2869e67f29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198e9eb0183667156a09556eae2c6a6ed3eec182587104b638002ffb407e3ef5072279ad88dcd49052e80634fe4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a7694bf3701e74965928d2937972de137f74b8219e056feab27cb46ba982732c8f2b6dc4cfe5f7a24e77bd58e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17453273b482e0a4aca65f2c12b57b460c46db21b198bf33f006ce9850a0fc3f4561679feb5c30b5dfef544afb8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc3a8433bfb539994bbc82730206e948f36dfdacd9f1000b0e48e6e24b6befc89c5d292002171210a5ccd30739;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf874b3cfc354c929baced5efa26ba2a4cb9f19a8715d7823293c2b9e18d30bff1956efaa5581500b3d7cce1f09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0923d8218c3d1533874eae4a5876c8efe86b9f4ff5548a7455a8f1f8142afa9028cbd35e0b7aa97cf7ed74a7d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd5360ec86959cc95d8a8165b5112f52bc0560a05796179aae4c36c7ab25abcab1188dbc2e2d37ff0e77137972;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19299053eaba9a56525e8bfd7dab0a4af8a1d5b8dddbe8bf3d6d65faed26f972b2f4607497c6b84ab84aa3ece54;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ed2c882fd527a63bcf008f47fb66bbad9c0049a65aa5707989db4ecbc6aa7f8376825acf98bfb601bccd639f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdcb7bb2b2956abcfdab3d272cff1c3bb9f1cf37180d64038d92f1a7a8260b0c1754391fcec4591959e02b19de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174dc606c6a7cccbdb61ee59973e10a97587199d2fb50d2d36c6d2f2bcca46282760d7b501c45376df8628f429d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2772019298fe935072a6af1fae77f54dbb6a07f37cb59286720d212927506e8c3b01f6e61c2819cd06017fff1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f6a1cef5730d5c77033de9d4e182f2ec599bbd1557d40302e5438b3445ec8e8e2929cc4d9c05aab5de6e4c43a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc41490803ebb0ee1644ce5e9f6598e523cb66ca25125d1a5f1b2482e18c57e34bbadb7dd3b7f5ccf03af25b6ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70e882773b432c30aaaff06d030f752606e1be5a9765eae906a9b56688983c3c0fd157c5f1c8fabea9f1445bcd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1beff2759f4efb05808935d20db9926daccfbd4cc12fd8f6571c7351f605a25d086bd905c72051731ee10893a17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b2a33dc045b86951775b9463a1739f8fd327f5f3acc6616aae90a709c01e8627409e01d70fd92ebf0ffa82e0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59dd2c0e874ead8a6e4568f90212438c9e085610824f24fd841ba841adb34d418e27790d8e413144d52782e4d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bd4cf919cf9243828a5cd437496283cae13a6884dc5f24393f7652c4b2b7c615c49060b4895391015e74ba31a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80d07915dd83906bcbc49ce4633480f34b5bd6d68705e5e662f0fc0f5b3fc34963d024f27d4ba803a00ee40ba0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1384d79cd20410fce5bab8bb0852ad68ca349ea2103f51fe5d77de911373217749521b8e87b32f19b7fa2fbac45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1936c7f6aa0efb2a86519039e9ed915e6744fb35e8253a878fb441e58128acbeee390ae18c20c45b947099e2271;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ef523e5218d4ee110ffc0238d3974ba611615211a96f5573fa7d5dc4b4170bd49252d8f775ae40a9d89a87cec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3269805a7507bc68c136790c10f726fdc2a63e977a7121f4b94bd04cbce04073a84f66ecd6d6b0934f328daff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ccd48a97f012d4dfdceb55aad63491456ebdc53f82bb8ca8901fb98e79ca54a1191605ab26328a4954bcb0e95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72c255092b2cdd2272eb97234dc5f6d38b6a0f55b7a4048eadc3a02965f3ccba197b4ae752063ce1f04722309;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e6cd4a92fb688a8dc085383d91570c9003588406ff50d0df72c28abf78c2cb56e25ba8191ed03caabd68c3554;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5fe7baf839343a5970d58f98f5a22e23ee6fe57ab48ebedd116ebc688585add1ad2f35d11138a504e92d8f173e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1191ebbc5f8d05a515a32688e1dbc88dff1570bc30fdbb33f7b7655ade164356810eabb42ce814a6912e893aa11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1342f6d9e15016f60925ec6aebb979f80d017468be3d059cc74f8590bb9717929197e3ff941536aae672387b491;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55268efd65b899241d6bfb8137aa2c5d88645992837eb99952a572d8260e2b89a81295332e0b9986e1c7432d75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1644640c5ae7c9faa37b93b36a557a27292c3a26ce723fad299996c548f84bd0c8045fa6d4968c024fcc6b115;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc44ec9bdf5133f1179aa498951420551e2957a48522ef3692e5a7633f0750374b881a0402189c69674cbe9218;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7638b1b9c945b0097c84951d7854d99e6b187f6095f47a4137b559f6121953d9db35c2740c15d3c5dbb3a98914;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8be42421258e16efd2a5b5206a95d7bd6b1ca8301d3140045afc3d73f1a63b1917c20442f4520ccaa3b7d14014;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169af783ab1af1efc7a19e4666edd3bf9b2aa2c8a1f5c226e1c127f2657f87951b19bdb9349c1b547f77c20c4fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da01e4acf369c71ebc2fdcfce20dfa5a60c61f5d69cf328d824d7a5bdddec0746afef1301ec1a615d4da3692db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0d960e12c141a333a079a8f86810d79e8b9387e03919e5b842a4c1217437ab7c9349f54c5d2a038a260d28c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e56ec4e6fdc73e6965202a89e9e961bbc5f43ad8cce312bfc767359c87d117e5a533e88ef4682b5802aca009f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha859770ba89627d8129bf45008290fadbebca7373183862feb8c83a2a03cd6b04008ae53d4763250f6dc39464;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156502300307becaf8ece8573bffe1a0d3c007ff185d3a6cbf4cf317d090377728ef56098656f032c037bfdaeb8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91f3fa9ebfc3ec8d5cd174e1f2db8fb621d855c377672f6161d08063ddab96429d3a123dcd55d914410fffa682;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae46f85155ede10747c3eb9794ffb1c5ed990c7806f1a3ae162c440c34deece3c4e584c1097e3858a600477e38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb232b51f33eef3a833ada1e244f119a83431fd18b80667903ce0c7fcba6f06b61f307ccc9dff6a3dcacb25efb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae3c4568c7958b44cc65bc678bad0c57876f2b7bfa0af92d8b58d0d0b19e7e73b4a79688c459c868e7be48d6b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f928e97e702ed993f2929f643d19e26a82774a2fc0994d714552ce4b6b391763c9bcff766361951e9c4c486b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136d0ea21bbf7288b6e4f0815aed26ad6f5371f6adafd99862070a83e9fae79f1142952bc22e4828878d7e82591;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc16a1651195adea7c843c2d360c66967a6e2fcf9d02abaa31e81ac448ffb689aaac2767948cd14ac98c7950c16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f9b08f77bcb4bdc4e70da921a0933abbb36dc1077674e64f8c696027221a12ed147fe97fb3d2375bc2cb0f70e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3be4006881ba2b914b1b33683e6d36951df420fa351276ed53d41e8cfbf0a12627534c45414a9bb5cef77b9697;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110afe043713c27a66251d5fbbacc3c7be2268fa678ca22ed283638ddb6ec031c7bc2133cdb255815758f25c981;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0fa911ebec03f50ad3656dce4055fde4f97d860d223af0c8f540050d18bdafece256d4cfaa86b1712b2158a43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfef82b750b25f016e4921d6e8d77468742a3654ed8380f10281eec077821271c4c734926b8a9af2375d9da1acc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a14d22f17c59106ae5fb0d93b1f126321daecaa27a31591186b104da27ee2bd7eacfbbb195d84c4721a116e1dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b8a43b5b263a49d42402d1e3372d7b5ed7e90478c7ea5c1a7cc22ce39556f961ce6ddb4c310312f0dfa1a0d43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h875a3dcd9df9f22d22a1155eb9b4abd94c978fd72a3c6f7a77d40dc11316f39a4de2457f3c5c57f6e0e6325354;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffe5be26aee8dcd52565a267f9f28b06a9ad83248a47ec360d57dd5ad199c9adc929cef963511339938a91fc04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66b0e04e952393c36b0e99d1501e97ae16ced943ae02e9c28a87f73f776d8c0fa6be49adbc695e42412353f9db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e8a98d3670986840ec12d9e70ff39708c28126439748777e6470c966dd822b6e08e9965d4c55238af7279f591;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5833cefb8065b4b16b0ede4c059f98a4e91e5fc704681df2c844357aeae7e15286c9ffeaceab8cfe33b022238;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e5445796b1fe454b1c1006c3ec8de2a4fe3bb33c8af3d97358e100d991e268924e58d49c6b94923f8e8a39482;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0cbf88c961013d9267420d593a94c3e84b3f1dbb6f6d40ce6561b59457113d96894f7bc4dd85197b819c500ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182b3218661bb1aef74d9c5cc3e6d3f73d7527171faca25ab73fe508229e6a384729c59cbab089f1c7a6193b6ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha178020e54657379dac45990f6f858380a9dea4c89fc152508bf71f111029b4a6250515673f7cdde367be35314;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h796fbd27c5792e2dabe449bf596a3d36848a58c131ca0560f36f469c8078cc4ed7abd94d6fc38e1566162ffa04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9020b4e695408198b79114fffe16662a5bc225c15084ccd14819f8c361d6d1dd9997a64d6de7f4658fc65562cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1351cb20f2f5eb1a3201e2162d07a2415718f78cd51c24a0c87875162c3e1bedcbf0db49c03fa7d4c88d0afac0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101d6a6cf00b29751333e1c42ffd999bc87eb8682abc3116b681fbd8657be37e4f5f9e018365c3abf40c4469c4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1024239762c28f248e8dfaaf52f6f945dd89b2480b56ae30a9f14008efd4b7806036fa3d050793d689d0751ae89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2949f4aee45b0374732fc55c03e581c40b1c6d242e07d9fab1742eeda8246648199fe5b61624f0c1d9e029a50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10079fbee698c86a7dec3ae6640243d0be7c7e0a8a634235c3e5bb751c56508b39a95baf178ddaee9eac03bb649;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13477db63a0a5ce6a34681cbc89dd3c21a3f66379b0b1aebfa1c67bdbfc23e49f7f068a2cb5d3c86f840192fb2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h656128f122dcb41b98f7d9d9beecd264f4b551a558ec8ac2099a59a5a2ea64e44fe2dc08849fdcf49489fef703;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187fb3b27aa1919d6ce3c176c569bc0abd9b2ab9fd546d4cbe019f8747e3df232dcf04997b17762a7bb0d8682f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133cd7ce84519711f2f5e765cfe0eb5d39fa001cc1904daddf9e6faed17f4a950ea30ac6830df3ac51c199e602a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd724ba96efda52fecbe5c4f321afb69b7ea6ba58aeb2dd1a751ff01f9f9587addcd7dc52550d3f3e60ba754cdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha87431a981885ac40cdf73c7c019a2039722403ff5d53a2c0ec5bd02a59773c57d4337618c934b349566b3d229;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3638405d6a88dda1f8aa64669a1ebc958445603940b4d7f86468b71d610b88a26ea417257301935b9a302261f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149beb6fbf4203daf44d9412881938d100b593d6138011a0011c54b51d42e840dc577ce41e86075a9a2999ea97c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1810df8b9559c05b711bef76c93922279bb4f4328e76b31092360e4152d6c1e23f6155611d6e4c8e31a2836cb1d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df23f74fb4c79d72dcf9e8b8e7d57b32a14befc75d6d6222a6207aab57789d369cb4d495d2e1c390c04f04708f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd55a6416bc29ea28ea09f0f58b263ea195b331a4c1e2c6456c17ebbdd0425a14f003c67b0232262cfdcdf14cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172fee160082693f2e016d06e07027b4d191b49be88e4a479c1bc2b138cd37ea97d071527c9c4e773fe0af8c8b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cfdc2dbdfb66c184c84d71b4fa7650fbe1b504db5db523cca6bfeec1c21368a8d0c95d7f63a545f361629cf4d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa8df6acfe3c85272fa65460c7719be4bd97f9b3bee7a68c9ca71081c09bccde4932a22b4dcfcb855fb2ca8204;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60dda38c0f2889268176156145987c5109e51abfebe4aecab39d9da13e297e9f2654ceba13e22e5e16dbfa915b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65f5fd7a36962ae06c6e4221f74b96a6788571478f687b76f4e4314d52e8d9eb1d2bf8a41893197d382cf9ed5b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6767fe97f33d8fa5e0ef70a4aa93c5f67f846bdd9c6000d353422900c8ceede5cc8cf63c3b867707a6ee0a1803;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1001e74e3ec39965f96c1691a209f8682c33b22633f88323960845993a2294730ebda03d25d75689180bec3cb00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149225a4e87d56da976fcff769b309b07e7e7f31e6baece0688151d6deda8f5e6e99e6d6a075a2fd873190c4e39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9605469e78572852229d88136932ad6f362f48651942875eb3c50caadbdf0bbfcc5fd6706dec5c6c5119ef88b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h897c229d9562780ba841f2f10d22469a2a573f19ac9b2c542790122bb0df16dfaf8f152815b4e1da3fe41bead7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2845257ad1fd3ed4f482d99bd8005d70e7d22ebe64fd083cc1d7e473a3b570abc19a743e5b209f9758fade1d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16587280ef0f604e8692b6f9445a6f11d563fbb14b842426f8e11f59ee421fd172948b4b9874c1b227bca13f167;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1857a7f1abe6e2929e7fcab0913a1ac2fac8e9c90b2a061c3baec63a40a8fa26c0740e8b0dad802bdc548051db6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3409a3eb1ec076f69166d2a96bdbfdcdfda3cece6972fcfe55cc4452ebe97f7b328076fddf00ba098835de0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ab9fbf91b1fa8ff511d319f56df41b8f5a638e85d62f873495ef8519f518aa5d38e31a787c689bc47f8400b0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98893a321c06eb64d7da636a44992276aa42ae9481dcbb8a4f62c96c61a1c9c32181f0075c71367b287b4e8ad0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfeb9bcb82e82d97f8b2acdc60c14e32bebc977e4a63e0a08b2bf62ad1f5ae51f5e2d62432a1b137a550b2f02b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfe37b13cccad3a2a5b2e9922ff256bf11d47214d3266f8cee5b38e8ecbee09249496281b85831fd7312772cc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1564a69751e7e20f385b81bb7bb1f9d988980c594cf1a5faecc357cdfc7889eb2f3d54b9971c751bc74ff981ab0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26df68aedcf943c1c5d28baf40179c733cd077c71ffc8e6c0fc044c10e17127ab3eb3d81454cb1e18a33673c21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha21aa44496a4024f42a6402e8d4b10bac2d97181a29d75c5b421368449a373f3cd968e6c809acc76ba5efd1c0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b0c1d363b7a6391dc973901268e6e9f4077516072b7a91c42c77fb5b2dce82e8c28b581e6f5954c30168fc125;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd01a41ba97a6b3e0fd2c856fbd886f7651b00d6950794e3ffbc2ca5a44f08594905f4ab24752356596006bc52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15cd127ae8a28bb17a206f17da165e5f04bd55ee6fbc9f58b2e7aeedead72c5bb28b05981f09cbff8756bc56043;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c784cc6ae27c421f03985a6cb44a080237cafe5f2d54cc5e9fc6373c70af409da6c568b78c2cd06cbb95c3bf6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60d1cf6b7ba191f56cad749e3525704cc847638a425ce46e62a8cb4a65ce1afa0471971c2374b3754dc07818e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bc70ff5e78888ae4dd567f0bf4fff8d32198cf6d9a8fad1fd0175039d93835a2c9d6c71ccee4e4fbe5d848aac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h655eaee02841915c987192c4e4580b8fe8fa4c83fede29b0938bb1558736fb104f29dbde5336871a6ad53b8805;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16180a7ff29105f2cdaabaf4bfb8baa9fbbc6c92ddcdb9218b7ccacc837255dcf722d38b89da76fd9206f729162;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b83453ec780e188a0b749acc8b8a5b3bb73a913668fff2a0c92a7826d903fddaeef410b04b31a964cfb8a0a2e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df0084dd14c82bf20386f6d260a14bf599ca2b56537d0ca2931e1574d93dfd62202a7c88771803624f40780e63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24726c7c56dd3e2ab2ba6c2fd8083713910e9922ac5cc93ff6f157ed2d301e1ad1cc10696376b3690ce63413a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d2bf6afc7fc168e2c0a13957091f3aa21122aaf97f05dcf5accfddb05e36c64c67e364e049c0688837b85f7c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6ebf84fd7bd2b6bed99c6b64033efc149704cbe698f502469f811a4f39fc2eecef6c355ae977c3fa5de326e89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa55fe1b4961878dc3ba4a6134b644608d61f102bed59406a467dd00b781a882f581085586ccfb560b960f9b68;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1951c2e64a227093ce5545b5cb3480ddd8ace4d63fea494d3b7ef26dce5473e406f24f888e205e71310c777ed5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef1a97ea33eeef29eec43479270fd1ba0c36954dab2bd7964f024b413277974af86d138fb339e0bf42ddb92e55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20c578b271f2096151cb030b03fccc85a637b4c62468a84ec44bccddf2886ede79e5468fde0db7bf38999af046;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb40635b903d19ec28e5b33c7afc5fd9a557548723721b56d413b7a61fc3e01ff83228ba77cc7776d340cf49aa7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f116af8726e1593227a2a2a11f9bbe736c81de314a8da0986d2566b1efa99ccdb6b5ba80608141ac31aa0d808;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc218cecaa84d1c11f8e2155beb7840d12d864379ba961e609e86188e850b20dfec5b2abb4bab2e94c6c29f1596;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a7ebbf5129e7859e670b0abb60eda8299b1f47fe96ad1b7d12190d238150b8a66b3ba99174619f3d1c6dcf7ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1515befe6935d19f5dd30c5a16e970bb396887a9958c5471d2f4ac6674f1e6d1fcadefb31522413d1d1cad45b43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d0eec64c80732df93d7148694b92c83d71fdc9bbbd9b7a5e029db334db9032ac04392109af3d259b0f4dc9623;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2c8975aac61fd5240807a5607fe2d4e3ac8c6e5c36ff97de28c45236e7bf7441aa4405d256cfcb7f9d129f6a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b28a8da72d011401778cda11324ac68a0ea2e7abb95bed64fc90e2ad30bb3bbc6237df3090aec59a81579fa61a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b90ce37d2a41bc140e140b227a39127a28bcad801430906ea99250fd283afb25d85f3bae938bd1b0478484213;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170fc214dd04ac10888254e2585785f6e59d938c2c1d97109e12d5a33363e2e882a3c1332ebd3ddcc53cc51d4fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18934206e5af00148bd2780a2849bc97a64f52814b22540207f2f5ec6a51ba92c93028e382740f3f8348109ce5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1435855f0bd7f50866ebae3edb99ed994fe3ec2e3cadea167d746d16937244402c27c2d91e6ecebbd09aad31991;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bfc6365f5647f8869e1e86a6c2a5043da1e2b8fd0dda7ff44f669d4ad7381c49e2cf6acec82400042b4ff5dcd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e73f60c9b3555d68cb1a30438684ceaf1259b2982c2ad75db136d4a4b9c06ffb6e578963d50b751d67a3a2c94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c3bc45522950dccea7e11d06a7d2c9de78cc2c96e68293304e46cce24f96b836e846c787d83c77ea191e38ef4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b3302393e66fbb584d021466f8344a19a17c7fb1f8eb26c09fa798eebf4fc370c042f99c05d91cdd3d83a898e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58892a3dc8f05cfa0ad81d30139704dba568e8852f24003ae6d5300ff9700092e004b5a3c1796b4e9039bd054f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1879c15a1fd529a0b4a457c88096cc06192b796fc7b358aca2034ecbc611e6ef78e1aa21ab8aff1bcb38dc877d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9bca55fde21fc35180aa52e33589d417d357bea73740d575d0a2375ba4b80dba460e390b109fb6992c661b5e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1944adcc04cbaa9ad312dc23eb81508e828d0519b8376db4bd08a5e69aae1c7c9ee309dd8a6031c8f30515aabc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a7ba6a55546e1324db5caceb4a4c3e83b55947baf22c8d33bebda514009005bce544dc423f069aaf0f3b91954;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a541c78423ea64670222689cf9e054717aa88ee99e9ba3c5e6dce564ba35d068bc8f56724aa57d42836762e1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa5566d148a6049b7c70452cbcb6ed8ea32d51137c4639613b7a7a064ecb382b732194f8d088d0b871e09310a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1989c427bc453f59f762ca1febc6d8b9f2d13cf42ffc6ab925c3fbba8497d9b277a9a656e6e3696446de8a3c2f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca18ce29aa298eda05948e9150f1b73f3fc654d292d5cc5beff0b62c391034da116f9ba2415b6b1c6183177dd2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbda2c4d09b6d3d07b740b6f3568950d2585f363670b33b38887fb80106a4125f5ad2e2fa0ac2b8f41a1dda784;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2f7f8022f1d3b6efabf1230fb7bdff5ce5ad2fd57c54f3313bd42a65b6f39991449e1e6516785ef14ec809c22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10283dc5f026c448b96f929327efb1a929b15fda0f42960d0c8b02e8de3c9643dfbf54d5e60d9c70793f51e5456;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f14ab73766dfe7c55fc9f388e0b7614e2d2e2eae3c31256ded2a8e0d8e7a18c6f5fea34d6b19905228b69e9d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17347094691711a095f4fd0a2f10e4c9e9d6b398724adf5dcc039ea743c1edce1a2ad91f10bde870be6b19ba376;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd765f1411225e8d8dfe97f03e7508f4cf381e9ec30aaa7604a76ffe161d1aada0abff4f9d94f1f49b0e68fcd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb78a028a2a5a021fe362b603d05133d54425162cd25854604e2a01191707014c64f5206195df828a87d798ef7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcaeade45572bc12e0eef5d88b4638bdd0c9d173fea35b48ca4ca1c541f84f91850e075a087a30a33519e727b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f77e092612b294390bd33a20631f836a15cd1f34e70beffc4324d56cfaa27de772632c14b3e592bebb26576b3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a046e6ad7938e76906014fc19894c463e9e55b982bf8907d583851ff9f90aafb8c1eec0ba6409547464d64e326;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e5487586cc3d175e692434229ced2ab9a2e643305a2df0c612810ca8a949dba96e598718b8a00f8576c330edb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29875c425f973d6e85946fbdb9cc850edcd86cf3ce6c721e561946204b863e47825245bf6d268dfc4849c38ca2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab10adb93e0ff44d02d50b3d00e1813c7129b5c347f42d7333f85704eed07dd28e01f652398fe29d650d2a8b62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8adede12c994b23b942162c549f6902edc6d38438b0a52b0666d1ea2902a5916812c64b008ad685f3353759795;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb1a15fe646899d52bccf92b0b2a5117a22f444ed57ae3eb422ea8b3704d39274780597096cd4b82ccc3374982;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13780eabba10e8922ff50dc4d37afa357a6ace8f7abf57df47cc94a5d2c81395e8c2a47d99b3e32e7d98c565e83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164a4170c9d0fa1f367ed6cb3244e79fe419352993240d34e241ecba377ab263d6ee99e7c53e55d77f412f8b9c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1150b634822f5767ba47c57c4a5897aad1cc72a53ac906eb99465d2581cc2dac5ae6b6e7d4a1d2a0d9c555d53be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a8b45be6ca1d058cdec82d60b23b4503c935a292d8697312b1f4350e13fe1d53d60e594470b9b38572658404d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha42b43a62fcd01d875e37da518a9099eb876de4134e7daafe04dcc1454bef75868971f531d37e322091ad0670f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151c90907875dff328b1e1a2f242622acf9be9770a4375976d730a65f697336b0256ec5369eac5e0fb67008a01;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3b992f6b49e0842b5bd481ac2488c58f69d09e3844c5ceca1706efd012327b0bfc74f459732e8e32bb40dc181;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d16ab8165f839ba0c43d70e7a7de42b85cd135b986592fb47790aad896f419b4b84d22eb10b7008a1d913ed662;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d02718e4446aebaeef743057e38f0575f582aea014340cba4140be1a5b9d7cc1963d22b71dbc2942b895639f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae50906d47fc125d7ec1db651c11969d39b481807d6bed3c89728a4daa4bb2dcb56f8f8e6a69e89282abe19645;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1061831f79a82ded1d51f72ddc4b2ea52bc66c24565fd4fe165af8cf8f0a18e13b8dab403acbb7386fbf92f7349;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14605f33266f2621e536b5a639338869adc9a6ecbbba3fc0b43916147c6fc36bc2d35270f973b13b5cebedf78d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1115174150ab966816450ebfacc4c42e295f0e5fb065d227cb5fe94b4abbef804da78c80d42de2856ff26adf833;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d854f17872004adce650e523bc8cb7cff8eeb44d6fc5524d9504c5c2e863ce90cb83644eb3bf34bb4b1e1a3bf6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a5cde7b0f484ba878d1f4cd80384c65d075be34d48328a340b77d4e68667e05385b7814b092a58db4bffb201e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf15796f966cf47cddfc5c5df4f7f38c54f3c291d8fe87f1f6c79f95a4a87132602d31978e29be5622ab73ae7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h433ebef39ee74f8dd13bdb3a3f2e7087f4b290365a26d1068b3c0757129b296bfd425800aaf8fe66911013d60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16dacdf2fac24b9605dfaeb8bee913c962381400142f04773a9012c4d87b4bc3007847b931385b283ff635e0e73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4d74a98a30a177ce5aa5870d69204ad7572e04888db91612d53b9cb9eacffffa6e208cb610e57dc029861b32e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf951692de792a9b2243196baa0dde8b6d3c3a629c3c4bd7ca17b80dc9bd145ced0da7ed823d704f4540e8963aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184284997af21f552f79be534876d94d0aff5ccd424e2cd7849cc5448f13a5e546938e629ebd58f2be92d666279;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1040cd10f1ddb86f7a05418f0df955b4a7c37af6d8e628bbc2a196fb0698057f0988ff06c15c60cf716a0cdf21c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55f1c11e72479cfc6f036befed16a10ac846a67f1582a6da760fb0de74a5515bec99919be12461b50d4908f77b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45cda431b886d0ba6160a0c090d631b3b1ad10c34507188ddf4555cbcde973b0f55b94786f16d79439efe35b73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6bb091a51a9550cf9a76baee495fc9cc3e097a4c768e4b58354226716235b23ed2ac4c38215969df156731952c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd167a1f6dd6dc69ae62127be71c632945dcda191af95fa0816f052aae27ece2bc2d281219b7506c672d24a7866;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e0b7400bb19b7c1fb04215893c9ed4881ea14661bdc3279e8fd14000f4ad8ced75006ff6fbc0c3a4e38530339;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h350b85acafc3eb89d71ab8532d0fc3982a3f26c68d4a39d844ba5bd03e0c9cac348a6c177ad332e7aca1b2ed45;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda9d29f752759dc9df28a68a9a1e1649d84e881fcf84bf56f42f5d0c3dfc6ae4ff53600b8f4ee517699655137;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he6f90202a31949cbf287f572b96e4eab966b1c7f55c25f9bfa2522594f818fa9a521202bbe132cd724fa52a9b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1908d73d3b1ba546c1dec822f9d9d80da7988c41263c385951e3bf490e528508ada29e1e491246499ccac4152a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92bfcd7379935905af3d7685c402f739ac320e78e0f2a4d96be25666b5fe4dec1083a4fc42799abb4ca7d2ec0c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a84398802679eae9f5df1ae317eb59f36c695097f09c45657f1a8919d4244f753905e90bf9f3db7ac761ed140;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53a9c659794b12f414a79a294d333e5cadebbd994bd4b5692cf1ee077adf80db7afc2535fae7488087c5feeafb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69d26af07fcb9e7625b8bf530aeae039cd7742aa12721a6b19eca759fbe6d3a78644541007e7db7b4213e1a338;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a19d5fb91ff4b6e1f76f90639f4c4d593eff5d33cfe72c95b3e83f472ac66df9fe2d3cdd742c50fb394ee453c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a5275979fb87c870ac7e5e7c3d6062aade6d7c04408167ffada9dc6d3d3bf62b63cf30bb2273643e3fc209cb3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h660da7a2555fbce982830d0c34f3e9954a0904cb1eab85d4020a07e617c6dc68785b9bb289488fb670a62e49c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19817d079448b5e68670c57a4276eb4728694f45022451b42d1fabb0e77a8888cad61b2ba97626a045ec71af780;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae8810022546f0a01b560ad0d832e3b8f90ce9b4d6f0d764403b138ea9cca96ec74c2570553bf7cf9854e09cf0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ce71eae178793549487ac3d80ca23887cdde38e723075e46df2377dd0162b30b419b1366dbc43e70f3f6078d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h752c45916e0d2ea4e8553fd817ac5c48fca01a92fede3a6a1a2291a4f8b55ad1f53f04c25b5112a8f283273fc5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b55aa0a0633bc93b82d671968fa2de63855681d3db6f3e8cf50577b49a825f1d6afee41493391f3824366f6d86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1249530a685cd8af91339cd96770cd4c0cbe5edf1f1e303d39aad8cfecba508f2c27f1d723953c0b3235ef3738b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc37e09619d2ef02756ebecf74a5f6a6f322cbce0fb8450e793699ccde8bb0929bd12765bf619d4b490b5fbe8d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76a967664721e92401a7b4e91de7d27a6d8d1ad82f2d533b5f39b92589aa3f05f0e045bc9956cd0d0d4f2c7103;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15de6783e7f6ffdbfbc0167c5babab586bd4a0acaefa98d9ad091585015829d6efaa3c302767ae3e6a66b12786;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180ab6ed7cb960e89d6a091d50fb797a1219f497a1317f334c2526b4bed16486a154b04af1deaad08d09e646801;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f59743629531e510322c21fec3172bc837b0414f510b9bb61b6a2d336424c9a0ecb351a7fea5ed63096aad3f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1f13efa9bad6dbf1c8460dbe877ee9f7a755d9bf768d8d970587b9cd86d2df49194677d094a7b7aed0a7d0aac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ed04cceec6c848aa0d8d20099a156462bc146f5be807f9dbe41dcb5af8350feffd7c20e743224cc5cd7beff8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bee534e790a9a725bdd3f4d926fa2cb833c38377acd775ed6c31894551bedb9408637b692b260e9db23dc66a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h822b09817052739d0d28ffcd037813b95d79f411b2fda5657a316484285ba9b8ab5b6ad930e785638200338d0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57733b22e0629018949c0a56af5b4aec5f98bfd5efd02562a8cc382872746ed2f07b95ff995b8a614f0d3a5a7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a297c2debf2d8bd203b5acff1e53c64c4152464a2ccb4ee7f29426821250d21d8c5534ef337628a5548ea943c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ead505ce1d2780cef547049456ab7a4e4837d03442e4b7633991741065e0811e39371370cc00abbf58fdaf08f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191cb6134c838e8785822df22ff30d081b5897f902db0f8ca5453921196a13650d44b606191891ba720c2725a72;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb02706f7894d53d4cb19b9f5dac4d345a229b1726cc9ece7084ab6bc9076e1047c0bbcd25aabf66465d35cd356;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3f416e5b9934da52019896f51cd13c6639caacecbfbe4bd70ed1957d255930a165a1031ea9ffdad16d0b69317;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152f583990295dde20505b989333dfe2664e98fabac87b4757e0de77910e717b4c7f0b7a0b2a4e7b3d412068edb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6d901739edd38844a0f38c6b6c9db59748078e47290e5f003f553c6434905733de99ab93f14cf4a8d9fe023ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he684dfe5e4488348eb712570b5d08f33f7e65693f0f648e75da22c0cf59438c7666f823d35a665b77ffc867f3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6b1d0d180ba73404bd0056aa26b90bc4cd5a0b1651d31d5fe0d9a2ef19866fbeaeff2b6cb1538d2de6b505687;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bbab8e63197e59a78abf1d4bbd32fd02dc95c1ac28beefbb0a515fc1aebe6cc82fd9cc86bd7a2579b152ab8b13;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12743759992e637d26748d971ea74c4a6f2f8ceb0f59420243351d66c91f1942c1425a6f259772ccaef70bd8c14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16158f355b95ebe15ad8987b8e692ec82797df5fe8ad1b734fac406a79940ba6438607a4614b997538f843cd559;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda9abcdcc19967f9a8766100e311092a9dc9b067be1a8d79d15c4dcd4747977ca20d5df93554bf26ecaad299b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79d37992222a229657d77db801213f089ff758616a7b26ac511c1656a5070d2eb6a97879f15506e434fa672e84;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ec1b59be80d5e392b4330e9a345c17e968c549a80ee5dc118ada97d53b6828a6a15ea63fe711b053674be85c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43ea0e9dd6c81e220f13803bf7ea67566cb577ac2868292a6b39227490763c2813eb94d71f5cca6b31b2610c5b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h627ac45278a3bcb64497ba34ada83c02c3c31ea047415db43d13b1a7affcde6b8c46f489cd6be2ee1d71588cb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h157dd57385b0875d0eaec23fd15b81aa36e43870661c662de2414ed401d6aa207faa6b5bef4736cd6594e7cbb56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39a8b2664d80ff2c342e3b44db1934985c78bb2165b2f906bc34fe5f6f0d3953bc6be5e68db29cd91a0631634;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbf41ab895ed49db29d5a3c4bc3081f044f74fbd191db8b2ca5bb3b1c8c6d2abb07bc057ddb30946e2d2c867a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heafbaf3e7301c865e9c6c297bfbe735b38a8da75821289243f944892460773dd6801cd4d349d04849e51a9bdc7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf787d7b7d723cef7e0eb9a7504db37d9b72a2e9b1a20be19054e6c8940c49b36c997a3b966cc5818c62fa2fa19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbdf344f749a97801b8721c649f5f4be8e687534ade3b70fe5816ba0cd26ac3c1535102119226db6b001adaa9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed63abc62278db9fa49e84ed8883c0aeaa66148e168cd31d2bff8d6c39071e64d41059f02a44a84fa5ae4c833c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd62266457e00bf2db319e4f9810bcf464b41db72d6e777995de6546428c2ed75829b46eb417611d1ea249121a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117282104b1e3373db2745da4e53f6213ceac7aac0d2b4b9c864e4865dc6e39c59334fb2e9d600b97eeb45e932f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f185ebad18229e3c40a6466475b8a1e1a89ecd22b125a2bcc2c21f0ba26607ba606a784f9d8af8be0c817da3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40dd8da7b934e12684dfd0814abb33fa69786685081d69bce88a629a6bec92e3eeb08bb11e80141770d51a8663;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha956a10970be4e55e45a3b16e11d0a4fc5c9303efb45445f3817d2ddc21e9800cf774e48338e91aff41e683c56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e631c29409f97ea7d03ca7aa4ec954797e1bfc0f4ec2dee8304c9c56db8baec4497c618e5b04e3636a4ba2000a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bcefdae64042cb57e6b7003b45e61118920e854e172574e677e4a651c87c36a246b57895e0551438c39f49b4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1712ed5afd1b45cce5c9378f5ffb7af488a454367299cf549db79519e4d716d0477df9d470f4f977b2f3b48d176;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d6011ab4f04cb2461631f1746fa700e2f1fda7967eca339b80c000e618ab55a55c1e4bf323344615161855122;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddb02cec06413e721282af87bd450bb587a12de329e5b97253ac379798e346da39db44a1bcd5761cb8b98feb39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha301e0f6db89ad2b24d3aaa12f9fd10e582de0b6b289e468647d0116f026f9c7897388c07b53b6e01f467d212a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h267a25f296b32b4a8dbea467aa6a825df5b19265865e13faaf48e424639ea716a60af920692017faf74cc90a7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178f6a625874180747286427660ecdc96173551c5c2ed10775178f8568a2f5aa6d330ba9268ccd197e667dbd073;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8af0079cff3bd67975bad908fd40537aafe6c96a5a88501af9841633c1da0cf0590af7d439db10bb81544d2e94;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7292ef9dc84e633791827ae641f2e5aa469612ce6df229797297f9d09026e9b4e2fadbb774ae1034ce3a7117c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4e8193c8552733d538b7211e01638605e01f6ea0c4196c9c32e02f88610b34466177a7815d3db66848900126f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ce34cff4d98afed6ad6bd19e2493362784e82dbe758ce62bfc68856509a9c5fa46cf28213d0753b54d8cc6e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7fa965c85853db1e454ef58845ea29357d11d275700d5c79fcbdc4cc09b5b2408959134a8e488b04312b24a96;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1293c452f17215c1ee94ff8d3089440f0ded5443f89345b707b13f25f51e98a00b5d1a3e4b927dd6088c771c2b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h937bd57146a3b6be609974a26746eb409183f1047121cb16121837f504bbdef77cabb805e8617220149f11f1a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bd88332e0a188e1e0b348e497322836eff78ad81c24704aa8d6aa930fc809a671d2c33eac0d5f81e453383d21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3f240a969334270b679737fadf011db8a2d5af5ddb52c80e46c7bd3da9b0d909aa0db3408e407923df5eca8b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd78136c3511079479dedec4b54922af81319fe87629035e220b74888853e0682f27f9096e77de8520bc16b60e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cd0789c39c30330f46461035cbcb0fd0a3aaaf8ff4e6f98df13b9d188f540a36a79d22f267b21a42997d1ff88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4f86f9706764c49769141efa7d306e3648dd8e7157a119ef9974f88738af479cb3105ff7bada568c258535595;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1c6de48907379dc5a378b05df9459052dd800982d0d12973ca0bf3e1efbbaf3b232b3c386968b32cc86b8e354;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bfaf97f2fad850bb280f4979b1df9b95de48b5fc41b6f6b71f1ecd62f56725ce60dd9ef7c2a00ccafb0ee7dce2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1029e963dbc227c3cb7f65477fd4b2cd38b544e890cf322c5fd7bb9a57aa14a9e1416086961dd9cfa85be822d33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hade2bf7051e7f51540aae332a72def381553f37f220245de517e997083104c837b37b36f5c1d1e7451a4183162;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14221932beea5393160aeeb2c256832f4243dedae3184c86dd0cf52549da6f6b80422c95c3eb57770fb7611c816;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff9ad2002a80230f5b0d2fcf0aea245c97c362ef2ad40772eb0ccfedb115255cd479f749f20c24899f070df193;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9449f6535e4b33d8741ca9693e095104a4cf2a0c412fe476650940a06db5b7c883828df13539edd1afe468c7d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41b090b74e6816c827f33e084876ad06ab1ccbd4c4202fa7585fd397ab2a3baf7f259ae70a0e0d61856c5ad8b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c88a8f34af80a595e4b3fd32e98172ee884911ea6bd2d061aab94e5278b2bd0b7540f5d4965c28367b0aabfa1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ba01e136609b86be927001970c5d5a0c2967292502ca4211eff26cfb5e297a4f1a6db9da2bbc5290685966d67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h552d11274a41cae4339f8d96b1545779cb239a1b91f5284f758e35a13cfeab00b2196a31f498517e3f4e00a91a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13097fc05e9cfdaf53d8899b0233d37ff118e1388f984a1304b42f1cb32b5859b95310ca058fc7c070af9789745;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbf321a6b9f8739161251301b66357f7a1cf21d4367692e38659e10af35717bc68d84aa8966b4834ca6880afd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he027b0f2959e91ed63d8e034990bd11f648168ff8a2336805096addfd46e757c1a33cb583f7d29f84339a82561;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18998a2fbf862d41603ce10dc378aaa189534824966c26c3b76c7f9de1589ccdcd455aacfbf35119084178dac2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ff1fc6d0634fe7d7701b67710a4d792cf9138aebd9bbf9cc58246fb6799b4a463cb99372a2541a1a2d9a5729d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc19c1ed58563137145eedaf03fb2b7265659f43acabd8e087eb96da0c26dc59189db2a033fd9b9701343c8c582;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb58691f532689672343bf29bb0774f3547e95685dc7278d8b98f2cc2fb5a7354accd3d9bb18a0cd518477f5c06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15815cc21ae0d2f8ce3639a97382554cd017e03f9bf2f1530ea732ed1e5bf0bb277309ecf27836480e204a6b63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f27e44f3515e1fedf2ec44b4384ff1061671157cadc2287e5bd9969ba52f349e83e6e13fe65fe7953324e27547;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c7ceb2b02ddea48d1196b49021eb94ae5b0bca6ff097151b52a9d322f066495733f224e7e0296489971f307bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15192737d2136fac0c3fbe5a9d03f90da87a6a36b356a04f525863bdbe0140a3315b9f26f48b605948fbf766c38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c22185c6e15fec56d0562d316c61fab8cea2657c31cc7d00cd7d9ebf0acc74972bed85cd30ddd0d3b66ed9f2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ba0b924948f031b4cc2ebddceea7a01cee00f629dcf1f9392ba7c6c5c018cfa37df586a74b369fb889c128dda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcff7af42b4a68cc0fda207127f72a7e2cdbbb6ab970cc062b826c81d402c20c3887a39da508b10dc501a7414ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87d15c396274bab9c5ffd5ad6e2b6e42be6f6a91a0a909083edfbcb4d825964612365162227bfc0e8cc3905c16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d004dcb17e65502ad4530b709fd4a376025cfce6745db89c87f08d29dc3b533e7c1aca36d49590b600e634d210;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he426bb61350ed7b2098bfc069f6c9a969687420440eef842e9b7ba3d9412bce42c0cdd058828de2f664e150ab2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a98b780ae13206254e93311a6847b74a1e611d80a405688c79748004bf7e293c199656b84d870bb8c9f0ffab60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf5ad3b1bd983e5df8ffebae3c90699bed813e323396b0378a75690d4b6b0965dc4c81f91d8706c7fb3a0b68d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e1f2665a3ba49b8fe75524229fb36a49a4771599f3d45acea35e1a16d42efea5de805eeffa4e49b9768e00579;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132e33da567434d663155721547d6d0025280630b3b658eb312cb5536cfc08f337019c4c9c4a5e6a13a2c5652f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ec50c2e80a62d13fea8c4f1d4dede0ca3413d1d9080efbc953163a2315846565a54bed3bcebcd581f272cbe52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1b5b8c774942a2b839b00e44bdb4f4bbe336e90da5e39a11882e92fff5557796ea58d17e2a5a4751376b5ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4acff210b575e7da6319e813351381f2f1cee30a532e6f788413590085438f629748bdbdd47d524744bca16ad5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ef8cef958c7d7d0bd583d80db882eeb1a90313d962c0d025c1ecdea5bf8f25ad4d911e8d3b65ab836e2cb3261;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb60857f955d7ad46007c0b9a6523ff80abea3b1e6a3abc2eb9f0b3b292d0c05f689e6b1b1e27f94f0eb5b4f38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab8ee2afc182e70aec6a92e1782756a19c6fc1c0e6c4cdb591f3be842e61acc50939f0e03aaf915f0cda2b4247;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13aa161d932f59a3b109d8dc1d054aa2b01adb50e3913863dfa0de0dd2ee820f56ccd7592011d432e292337db98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he72d8ab7806354f02870ac9308a9db29d94d99a5bb86a311b5d1f79c66992c66da8d6133f803a6effcddbd4267;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f0994d8243bca9801f6cfbbf537bdc1e2a5aaa56e415c0beab34431d77403d4c71bff0a07af3e2b4de36eb00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51793657738e872470202a5911139cd29ed594a0f9a01b036499674e05f60b0303b02c49e59412e2967638e1cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11aa3e4453b3af1763ef1c3558e8193914972bcb62781e95b9a3558f25b62471bb158529a6137d0746901760c13;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cca1aeba7b93438456e0bdc7f345638e2a628a3bb36aed3d05ca6458b9f007f546a263da3162292de323a1943;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9edf78cacfda6d27bba5e97e51548530be6cfa602ce4fe0987294b03a452edd3ad41e43f1f44f4993268a8d95e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1074fca213b83e98274ee18e3f56903299fda7b4ec1552daf8b9047c99ebbd82d834b49b999f741169616eb1303;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e969f052f8a7024df2cfa696c2c01e57ef78a476b2f1f86e516299c8697fe2ea83ab325458d10da4fb6ec555d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3e68431c621b5a5f667aac1fce7df5b18e2f9163fe4e00bcab66bf8c0114fb5c147196d66fa024cbc5cc2f93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e32d3c0f31470463646daeff39d0fca91065bd69a243158b42ead2a4ebeb2d25a5ff48315ab7848fdf40e15f5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e60e009ba78abe8ae82792eb9802d2e718327202ec255aaa7724b4c93dcc7f00c304a32a264618863e6bed4931;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd72da242ecd31489316c85c8f877b0313cb26dca337c708402a6dbc583f6049400a8fc3d3b00c7c515e4b6ea1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2a5c70e9739b715a933f1c6170bacd7c415364f9742dc9fa6148c6cd778ffc84390db10ad08e07e794e9d4fe7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb38e2d7f0b4cd178a5ea5046a63b57c1717e7c85cb38da820c370a783a97873bb4462968819eb5fb23e5bdc5b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee0da47bf6ebfc9d52a257a4713337c5cc56e497efc78b8557bea1048c2a48c36675555a35529c9a74ff5f1c00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd24016ae85d9c4dca9b79fd9068879075b482f7ead46d4521fd6c4d6694641fa9efc188d12e72742d15a03e9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c1c2f3012e9c863fde062aaa5941b646a2247f29f21c43e42ef963e64cdb61ac855b19447dd6525978463c8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a66f17d1c0cc0052baaafaedc5c7c70ada912793bec8a8342fedb93ccbf8c3b4d22d2364a701d4552b967fe149;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11939153476c6ab82ab37f0ccaef205fe908c0d128decc1907c7828bae8da33425d60bcda30376978a397aa9db8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1321dd71b448b03d49f1ebdfad947b67bbb97639bb8f0e1b30610f004c96ff787a183821d489e99c8b0d73b4c0c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0f5c52ca0614681bd69d3f253a90b092b42b3eebdea4731ae567f4673887c440aa9c74fa5708a746dc35755a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae4e768669673841919108108e4cf056ed740d7d63fcdae4043e52014ad4faa501f6c0da4a870c8c9b7b90eb0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193960ee5d2cc8108bcc9a745ac0c120acfe486b24cf7a00bfee887818fa0f133d2a7880508946cc0752b490aa4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3bc48780e3e6e7087c60b88caa3c01ffee8ac3ca25293f11947f4fc464e01d71bda744f583c97a22f2d7df33f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134930f1890e7e56eb6e815799cfbccb0d6f3009eebf649a425df47181c48223374055d9d06f1eed81033b2726c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad0ef1bc5c19b1416ffbffc355e9522631626d3204ba684942986bd8b40e033ee3f056bdfe2ac57e47fad94b0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfafba7e387faccfed5b5790941afe21c3198daaccae81d93d44e9f3a227be6697640f161a9bed69c7d7ab24cb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2f9dc08920b01ad0bce199b8c2c0f26ebe42d783fe7f24801577c0acfbc6aa594c8ecf2bf6affd1ba1db78fc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b863ad2f5bc776aabd2d4542158db133e154fe9cd168ec8610fef25f2337f9830c2dda96922e597a46a7f7a88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16da998e82bff0bb08c3f5d4aefe175fbb85e17884a9dac04e01b71d00e6139cba0c05f2448cef1c32e5bf4d6ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ca4cdb5af24a73dd76abb010f66a0351d68ac066f9dac85288d4f13437afd3a22b8f95c90eb4915573c1543c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133a34d7c1c1cc87df2ebbea58e8691f383c82d4503e2a248e6c4bad6171d622229265db1c3c50aacbae1edc5a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14596204c5692d67d3ac8f032b8848dad4b002e6e8660c86b2d0fa6009722f547a02d59c4d7d32c073b4cdbd745;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5627e0f664d93f230567e3a563a456a60065a33b28510e8a3249847c0ae1cb2b76b8e17d63ac547c2fc341a69b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f3ef48f6dedb2b71d171c5d62033a6058eb9e80f290530b765602aafb77ae9b812d0187593d4af643a9809028;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82d18a4d69c0a9f4ab5613251c9137ed364f43886970a4fe1c711179aff9ab515caa5e3833785b69e9b390d7a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f694717de464d890e1acf6c7633bf76f2f3efdcfa750f62c3ec50eaf58639e0073895b9fc8ccd14c5750100c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135967b2cf80bd5e2cbed489cda027f13ffbaa86ca0a66dd71688cd56e42ebf93652fd356726c14f778fb051e89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3e4131867a599f38b04d975d4d7c138ba51b237ffeb8df831b39a106649c3b41103bc98ae613a815816276d3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a6fbc91e4c9673dbdc27545d7d453dec2b23a249937c2b33116760f5062990ec942427ed32199c096e054fc8c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99e890cf40a50f001921b297b5e932f4ef899dfd9112c2eca24aac3a1cc07d80a9d828bffa0fe53170395899cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b560d2f93c8f7bc6e203cf73f17ce5472d64ffc9a3066eaa45b247e7dcd26a12d5d16bc144b11bb784791a17a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ad1a8cc87bd2aafe1fa93e4fff8ea02e0539db0ffdd0f698b5603ce5f14bc2354ce116869ebbdfd400229cda7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90ca0ed1a6e2d6f061e2f8af2523818efb5f0d4f7702fc27921f83e5bd8336d0901aec21c1474c923a3648fd09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h669121ab673933eb881480ff15315255ce5580f0d88e264e044285a7e1de3f272a6aed5b26214d3c8a600b12b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61e9d009552e09b24864b85e883e420466b812a94cc0dbfdc2e67a52016e53e24511f6264018a602c5c25091c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10cbd9126733f8439d08a7fa6c9b3d1494e2f77df7c5ccb9ae017804930954175544e4c7525fc4c4b80a29c7630;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1518b833ff7e8a5bcfe081b90d74d07c2e99ee59b221ab9be0b83d3548a3c1352715eaf41e9afe8ab9a8f24a9ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b602645aaa0411a3ec0420b38972d2592e7b7205b9769439596ad681873772b5c5e742208b4025f76814af24e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91a48c073b59cc03a81cbf164e8c8f388cc60427822e2314673e9090fd3a766e14d42449d2e40bd554809bbfc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe197d0a9ce3f9af0def3f16e70cac1034d801dd14789f80a97c8ee69381148aa49b10ad66df29c100bce9885c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121bcffab75360e5d527e0996370cd4915728544200601fe495c0251f71a0945cd03bc786968fc747698bab7fd4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h704e2fa25958dbcac254e330a2cba032f3749ba4e88c6a2d28041766c335a4442be62173aa0a77880215ed0518;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3415cfdc9d860d8dfd15916c40c7e0b562c8d4f39b92b2041c19d9c4ffc3bc9d463c38666d9b783a5327b61ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3d619154e998f9eb654e0e913f7a239f21781ff9b7a9e532f55bd59fbe9cc6a95e5bf4c1564c157d0b97acd62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6437b17ac6ff94f728844bac4711c3d5860cab1250cf51c546d63f8a534d89d206814af4aa729008c18448b59d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c192bf525633e0a396f6eb6046cd2794e9f124dacdbd43e25bc71d7c0e84a5c63f249fc0c754a07dcc386643f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78b5283cd43e37bd5d4b2c5e74334fd168e7efd30fcd09e4e7581f244b49246484f51d8bce514d1f47757a2a81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6d8ccab230adbc8da67f0cd471bea95e76ab225f05fee46fa606a10489a6b196cde62db63e9d82d7686a3f043;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa7278f76fac48a6854b9fef92f20512e336571a018e403ca032e47c974bc2ec079e9616daaada7305ead03745;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e13a607a50ad2b1f1cb6bb79de4ae4d1990b76ebfa6218b250f6aaff55c7de0df83cbff45150e0d5b1e8b43608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb73c4b5c53be4eaf6148d654978816de6f2f77103860758671f5bd8329d998a5df9435e2eca328f844ba9ba10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4309ab32d261faeb1079940492f972c5579e3950e901572a69eb2c11f8b95c7224c368f9d029d0177efc190d67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179095a46702ecbab5cdb7fe520ff8a0c0af70ba0059d0fb1fd28d451fce76f1f6362e1b329737dc6e4a81eeeaa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f54f927f62fed0188a38a6d1e71034bcf300fda11d222e2bd6fa5b8b3d687417a9311961c2f81e8743a7d43f0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3214d3120a2358f86be64b8861f0aa38f2be5b24f005a85beb174357adeb09013b794e4096439ffd456c42213e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0361a3b8df87afd12fd2f7bcf17cc63e34884e59633ddb937befbb685318471d00d76ad0a8a212749bffa2cfc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3534d2dd00a684f5ef6f4860bda483954f24085ee30e99e5ac70e79bb282e67d799e48f8c3bc4daf233fdfc2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e51047ea74f4853437dfe5d3ff88cccbcaf569dcbc8b933a4fc46abb58fee44d45213307c8dc4ade0cb6108d71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5575b4c6bd3f66f21efc834a311668bcc2281b121044cd433d7ecc3a9042094843caf000e5e0a36bc7d3323d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af4f31f0bfd8bd888d430dcfcbb5303712923e0d4a423bbda91d7126d4e5c4fdf13708c7ef8d60f75bde9d6cea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166771834aa553e1b733ed7e8f5dd37e6704868957216addf71923fce9938fb3fbf3526d159e34963eb4f8df731;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22cf63288168f01e400c1fdefdb638a5c4e34a3fbd78c035030f916199ec5808a607846acf286baf5533adc968;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd933f99d09875bddc8bb48ac3a13e311bc4f9f99ade19297bf10e3143a19c1d46846604eb56bb02b273ca58fe2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc32c98124f723b9bdcce703f03673f77e7f0e2b4b45d4e7aa4f20ef8a691a1690183be9ff7d1261f05d659dd4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4ce9d04309187eb7d70d9059acb4a365e4bf2246f0b29de88add810910525e7c3ac3726f8827d02ebce410c02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3ceaf25e6cce84340c9ed79c3859e400a4964798c30851ee31c4de275afd091a10b8ff71b293b0e7f481179a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d784dcfc0df1f74174b688459ec7f87cafce7fb8791abf9f4713c16ffcc3c7d8d26933918a0650036c654aa6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab2220710c2faf628b6006d0ffdbf8ae5d01197d466d9b55e99e384990b9233148cea7da5dfc0636f698e00b86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10094ddef108a7aa8b7c962680e60b075cd60ba19f550d2e322e5c61964f7e39e3bf5f6aeaa6b52d3f22223dc8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9084b9279fa6a674de99bbbfe2ba3aeb59f95c91cf89a8b08667718dc9b05de01a66f6dd9282b3612be3587554;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27f9781c5d9b1a3e4bbe8501dfff44176a92356edd0d9dc6dbfe0314b331d28ee6adf826c27647c90a511098d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h677a93edb3f0e5b05da5c88ef90f51379eb860137e523824330bff7d7aee7e5cf577b746cdd0c7d6f697372060;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12467824ceb637525f293d8c8412586a574c80d94c6dcbe70b4792234e882ea799d85a762a4c096c828ee952d04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab017e414e0159fde8514e9017879a474fb7c46fa91d4884f5effbbd7fb8b79f68c529a3be49359e533c8de170;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a6593c8a2a08d29adf05ac73a3e7d5a405adb16248ae504343f98ac83703fbe35014a049438282c308b08fe18;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c216565c2d4bfcf64bbdf7a9dd9c0f26805b93d8649289a32c0636988873f651ac3fedce2327535b40703ed13;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65d1db69fe939a3db67a9bb05b935dbf67bebfadd8a8c3ca26ad0aed4a56bf9d1568a26fb1046c6e1b1d19e8e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13323a0720d7b9655a5da5734a515ce60010e7fd63d7402150e1d1b2a2c07f2f57a1e649768e37b378d0a23d444;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d1df7eda81fabe0c5886df2cb6dd624585406d25ce989dc33962140bdf16c12ae7bc32c729c320df146730d04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b415be9a89941b5f35291ee51b14ae5198d704d09c9716ff7e45736bb39983fd97d638f55ca657687ff297a2ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43656774cecdc26a110701522024a86cc5e45f793d64e1a377536baa452f6ac92ebcb37e68ca1fd848b80853dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121ad3a647786325822b097db7dbc1951cc0a6f2f628479fdac271fe24cd57046cbdcf21bc307a9eb79235253be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1597586974809721fc723af38554cab9e3f3b79552e3600b9915590e02b5a00854cd254cc1f740fede98f98e9b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had47f30e0023d6cf37c047e72b16f67dae4bbde7ab1e7498c8b5c26b2291be1bee5ce348401f29b187e1467cb1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131abb9f19aeb681d42dec2d2614cdc7b840700be07e1f1b699e23e4b1a8b328bbb204f96517b6009ac6cbde0e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b1c0df52eda02ca5a7ef3b2677b068571e87b6fe7939d70784afd1220bf01690c0b900c5aef74c40f207a3832;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128a8d3760e27d581fc4f1e0cba9646de83680d18049f76225b8ba3c49885aa225fb77f15964effb310d872a09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1711520a99b7824156cc653ebf078db056849ab62800718cb168cddab31b66caef9592876457c28d82880cc7529;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbeeb9d4318ba3f059656787bbfeecef459e943c6b670bb27a6d94cdd69540d8f55beec8ffefb19681ff998d335;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1e2f50229de22a49add6a3c2a16ffe689bb19f44afaadb5828f3c6fe7ea2b06b445eb99ea6093baa500873c90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb579301add3d1c43fad6860c8337f96a15d6ca1ab0253d1f05eeb252a342480c4549c31b62d1fa2c9908c648b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17aa79339ed149007bd53b0914bc506a962e8828b684d9c25f9128e8d8f0b400bed366f412a859ff3069390c762;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1d850a342e561cd613c20ec9852b3897b8a3bb1f55f63037d3e364e61aaec96e606938512d9fa9ab1f6b05f04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2daa1171cf307eedaa008b0029c68c1ca31ef436e23a54616b9d0592262d46cbc743394e1c76b2dccc15c58923;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d044e1c4c3d8fb15a524367a37858bb05c93559df8cc3c488f461c087bbf268f8257b355a0dd39e67d5104cc4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e48e175e8b37f786965bb1048b82298b4cfac5dd935bd411a0abd33db167a09b604038bc5a02ae9270fed4820;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc30b77418df0d10bf763f8e5fb6c59aeaab8c4dc0b3c905d628f342f9ccb97e05fac218c50eb2a5ae5207d531f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h211414669d142d0c09e6ba2ea929fef217ec917e508203417d2232f8ea908475522cf283fb844a0ab65ff18ad0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ea5ec10aed0e28be88ab4a94c63e98bd2dc00b76c3366de21b46e24165082b8384275f39d0e73cb221ffdae10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f98d3679d2b816091a6c4351bd7e63455cdab4755e770f9fd9e5a11669f5a34057c90888510582fd9c6b1edc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ddd1f32cbbd375f4619d0f24025f61ad8ffba3937d3305bef616854e313572764177cae746d84aee94b839a4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b5d7e1643195798b28640cfe8f81cf4c7ad6c969e76ef31ab810ef3f1bf170397c320d07f979036dfc6c9b31;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0bbc19cd98722967f615c589307a9e613350b8917085018d526aa9124758c6bf558d072ee0ce194f59e4e5937;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa7bbac5757ab578b2568c44da037ce1ec070943f832c0f9e5fcf85fa7fca86b9696020fe7dde20417d7eae7da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h651714247f65598c3cbb7eebe31ba8654574fb795ed489568abccc30c2e436afd57aceeb748c62878ef723a6ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5774391d0b661c3a6169d83286eda3f7a4a9b6d50c3a6e0b507717470a602abb5c075e6da3408de5c5fc07179f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176c3a933b2b55beb782d48accb3f58357d601c61bf4ac8ff5113c6c02cdd060f91700915bbbf15f06fafd3849;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80cd8d348ac04a76c635e0e51ba4a386aa760765022693a8738626564cfeba39efe1bfebc4fb04a8c1f2bdc571;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168ad04358af7867dae34c22918b4a42901ec68ed88ba659b804f7b89feaf89a9f3e650c910de3989a0cec06eff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19deb3fadd983d14a55f91073a380954011e5a6fa73101865a7803f2bd744a1e0d9cad9d3e8a41e94a444d811f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea361b922815137d0f3abe6f44ebd7bab0ada882f1a375ccbc9dd76bef69870e50495adae7f5d3633ca2d7f8df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e37642fca7215ebdf7c215930b4de95a1e63d4a2427057db469c5ebbef17a1c6fea079fb51a0fbe44e91a2273;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1768536317afc56c3cabc6c52a2c274802dac73cb7a4fd41afa825bdc086da872a1a150fb4750347a238d83bf46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7759e422dc5236b321c3cec41b0f71926b1bb7cee2cc3e19e0fe70ce0b045d427dc3b1e9db2dddc808b6309f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70bc905bc7e019b37a62e8a725d8735de2012229d74cd2b7d7ab1796629053948783f846bdd0aebfbd05acf7cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e1e865985227a8d6515dbe50ad3bf03677619b410e6a29abb6d4c206113f9ed5c10c84d78d9ed6b96f296b74e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138321713c9671df3859dadcbd161fe68b28575da24cbe205e1d8c920eed45abc06dbb9250ed8eb5f5b16ee5bbc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f162fce5e70ad99454b220a8f283bd33b97f091e97169fab6ed8dc496bbe183b0b2b1bc8c15e5757cf2deeb241;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee96d8d6e8162125dc7214f95d90bd06114d7445cc64fc953d956d9f25f0771366c28092333646a9fabb0d6a8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfb1771e91b8469dff9823479bb9b4fb4605da11203df934b4f945254e15436c524a5380509e73989158e317fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10643bc5a92796b4ea4cb83df9a5099419bb986ed4262b9356450c9eee9a464e77bdf16c8202bc4eac43f3d6ef3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c666e11706cc7790ef4485d94db669c509f07e2290f8e60664df1515717f010ce628779b988680ff0d31c577cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ce9aa72fac7c906ff7a4b98dc7893a0c973bfff62a14f5e6f668a7c7a8d0a721e0f5bfba23cbd8f5d8ce4c7bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb806323b2d8feca52e3ea11516568ad36b7b5a5eece27338b66709291603626c871d3f11b51ababdbd5c70571;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8e45b019215cd34d244f46f4fa8cd7b4789c0fa87ef5ec156c732f4b8195f5afb4a4b30fb905d8956dbe975d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a5aa22eb5855cefeb6cffe7fc701496dbea5838eb04e9360c4e4baccde1fc61a99a09a8e74a7c8c67e5ab84148;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf13a23ca81ff2232265e8353473b7d69c8c9619c5265b12aec173ace20e55d57b267a5eadf61d15796ede31d8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8163e06206dfe2b0ce62b305d350b0f77921c3660536c22918bc0150193832d849a74b6e02ec2100e40ad2d3a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h569b9bafdc740af95d901d126d97d00fd61d7efa374c925b5b09d1fb56469e72cdd1216458c5d66f6a49339137;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16bb0efbab74863c007bc4ec4a74a0de57bcd4c3f85a8d46ed4c83a81379287fb7f0f021c6cd3f80ce637765da2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1607ff8bf20f5b988bd0537503fb9800eb51ef6cbd48cbf3b2437684a7d509e5314347a834f1a41f794e98e04f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f2b26c8c1334c9ff73b412fb79d4e38a513180d6ab8d9a47344c3e22702280ff0865096e199547f34421fdbf5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce4c40b7f939da32d149db6f25277607fc41bbab5287b54436bd4e53ceb201d061d55cabfaf339c431c17893a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ecd381352b7bc1e15a500f1c6dee735a6e8ffd5805b6872c27372250d50ee4aed20ac1357ff8ca3b71305cf76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4ce27ef8adc46dba395a8e9f5acb325d3797f78744e8bbefb4d98650f6ccc8ccbf72ebe4c2610147a4b9447bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1173db9a8faff717e72db53a49c2f13d07a04302f5bf9c555a805521dd7fcca9847669d8ff5250b5e55b6c45946;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe6a26fd349577cab3dbbab0f6ad41fe8ba9c8f7cc410c947edbdb7816c56b6640c28d74e5c69c65b24183f2bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2007a6656b8691ec4de8741669d715648973dbefcca579115b94c40bafdec3f0f7e1aee7e9a064abb5fbd0ba5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b9d809ada08c7b779599d77c20ac25dc41bd94a52ca000ae7eb12d53cbc98676886b3e7aecc03178fa5d28fa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d9d7360960f3e65d1a79790555f468ef9e023bba8631b28ea40fae4d12947b7ee38be609d3bc61c145e26c44f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1678e9aa9de991d0dff5027c0f50fc9fae4b0d6efd0d275d9ee9246740c38e9631de9255b217b384dd76fe73266;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95a65feef764fa12356f5f43d34399d017a9f51720d9d6ff6135f40ea172351a204be76fe339350a2228559c43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f4c57df39a9090bfcf00d4ac4e45b9a491c4d2e064c9cffb73eefcf2746d94d2ebd58cac0fd1114d6dd37d4ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h667fb5ceac7106ace06197d7b45d557506974ac94199eb100f78ae01deda7daa0834e18734c8721f9414008fa0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ea019c06dbd88d11373bc5148baf2c626c1231edf6f5e75c126440f0876b6a19e16653dd96eac3ef20ed1d87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c76cef21f67bb161c8383413939b6682c3d3603efa28fce1639d45d8076303c091bb9559acd2d5d7baa16161d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8f4ec567390699ee283e729731a25efc6b31286762421ad7aae6ccc3d755f8c04116a49c480824e961f77f85b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc60bd165d1773b4f9319bbfaf97667928deeff531e25af97d76d57fba3e27f662957c3d8177a91fd88a72bfd1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d2ff4ad1507848716849697a843395252b1939d6a9ede2d598e4391feac8d85f871e4fd31e764b51631cf9800;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180b0312075e6c312e098bff5ee439c0638f78711806c60edd5524d70967709519a7be19e4a1d9f84cf8d92fc8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16832abfb572d5368798c5e9a9049309aa590cb4b5b2b7e2dfbb0ae41d92bd2abe660c6ae7dc9b0093ad0f421f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h129397fa837235ea7bcbbab20388b7b5963047de11d364a4174f6e389ac2ad836d013a6505b3f52dbba3db678ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cf690ffabe23c6e87185fd437ec4df1d65fc8dee733e63149102fdd4820bc147e78e59432103fc05fc135fd4c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c2f2766f07a7f9cede4f236e3df95c48df270cf965a80588cdec32e5239d09b2bdf3551fb59363114e937ab22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1729165a2379a89cbe0347f0e15fd3ea1869fb94cc58762547db5eb62c2a5c8b868e0d4627246c892506b75cfb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c3dca5b5ffd9a72a9461e5703ce904d997975b72b988e63b843d1610032f32f446ecda89d003d5296ced80eb2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e339dccc328028b0ef5bd4b585dd8d36fe1b08396235444c511ec4f70995a216511d30f48225823de77786b64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db35195fc4de5040fd2468a0de5a73345fcc940273703a8a600f3d67044f417faf914f528440c03a91ea574739;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18413f8f4b6fa6c28e7a21c02e175c1ac750fd071c7eec4b91e083e1111a2ba40871c6fc172354a4a6c166f75a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3718bbcf63805848b8c03fd18858526fc3a067c424095fa07a005b3541fa2b40f994ab761517ba752d7e52710;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h251424656c291c62c7fe554b2b75eabbdd728e6e53622e32354ed0d2bd35b65b91895fb03c4d6be3004ae41d19;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1493b35c4b08928a37f31dce20c4f264d3733063ffd498f36737c0bc55413f815a75f1bde6460f6dd16002ed321;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa461f14b0dede944ff20d316150e6ad20efb487738207485e9d7bcb9ed598fab9e3a29a4b176363edb4497934;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b41ebe2dec9afe042eb20fdc6a04904ac1d164767d969714ded1e176d1f9ef3e379d7a548a9a56fa74f7bcb3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a33353746178bf09c1517b9abd7afbae9051c1e756605736a5f61d4369457c2143113dd1cda16941f4e99bdae7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24e74aaef0693936e9a8865a60022ce4e687b587f3f277ac1d5e2006e0b5501b71e8069b0adbbd480f60346034;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eeaf428747d28aea72dee94d87b38dd0ccb0f97c6ef200708f087d6c54d52298085c4842090e6bfc85e93dae18;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1301e677a8fd09cdf694033fb1db2638ee57e01f95b857a426b6595711e96a146cd14c457006f78385ec90e8463;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fac6724b9649eafc2027e818ba84739fbc9109537d84336c9c15ab4524149969fb03504c47a90673989e464d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112ff975f8289a58083dc0098164d5f1c488bef814edeeb5eb94b4155c8b7c07ab9112076ebce327ae7d4242aee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1924139f926b321ea9e43dbf2ce00c1f3192334cab6ba75e5906480451703eeab5db736844c4b19ea32ad9f2c73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14eba272473adec7b53d6abb18cdaf99174d9ff1bbe583223b1191bedddf030425679834e1cc61eb592e23cb4fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf31c3ba63e454548a9b4ed8df315958d0203fbb9e0a22b4808657f8be59cc3f2f9faf27aa49c0d59cca46dcf68;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e36d6abfe1c8f90237f1af9da75b6eb6fdc309ed55d492ea94f159a6b076137a19ec56fdc3b1a23fd60034715;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5075dbf0e2b4adfc97ee5da2b58e899831e4af6e5d569dd28180210335027cea92cc0921be7e16998b6de3ba4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc20be0abdaa84e84c26c78b2ff116f803ca41cfcf07f47f9f361840dfabdd621b2f529ae1df07e08ae878768fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h843d4190019cba85496238464768eeba1a77672f7d7a0451b7a31fe429d1738749da3b510001076af0e710e8fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb077874d04b2a0d0fef3b64ef130442656d80a8368f09d033eca744ba3327f0809cccf13f24e5b4770214c2114;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166756b7cc15dcaa598c84816fe1ec2ce640e870f10032075500a518421d13e5047530dbe3068e09cb3e6ac604a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1ae0e19dd9ae5e10391e4203708a9b94bd2b803a4d1ae5ed0fbce46e92d0bf062135dc6c431dd32c9cea0a6e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6d3b3c1f0274b007e834dd2954892410923bebd7b1522a1b230895f920ede2dd6ccf5a09bca1327a684340814;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54a4561db43b80fde27645eaadf38bae1651057a280f206ddc997b153f5340c3ddb580cab098ce7da67a869f67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1235bffa0c80480fcd4f5446058d6a0f2f8d901cbdd38584d35efbf9f6988bff30d1daaf1ddf02064f2dc0320c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb73be467c5207e04e2c7084b1c7a9d2eafa64d2f75370176852707774e9943f4f344fce9b87fde6fbe3e24570;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3502f05e57e2150d16d678d5ea61e8c099a7e96d19ab6ae094afd094c9a363f2f79104764a2aba8599c344f92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaba014ca3a72ecb9a65628fb7715d296ecfa6e8b8dd458b0d669da36219ecb2ed495796434d05f188cca37e58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14eeedd515b3db31b23b7ea405cc7aa41f1d5be08ca69b0da42f0f347c043564941f4092f91b3b664ceb399a301;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3819d1a6a1a3271285336bb2ac4bf658abbbcb95aeda7e156f8abd4f70bc35b3fd74fef5a5d243c05e17ad8a6e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h518296d29b42dc5ac04878c9b83ce33c0ceb9b479fbc6c5e0625ca231e865431420957568464f2c2d06a91de1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa2171d45571dea59205f44b04a95f900f36b6d686fd81674f6a63f908d53c9e1823d61011594230f27a739242;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10814bc1480d8e0be8bf357b868f2ee4aceb61d70598abd17763612ab2952e4910a2d719ac0b23c1e9af78f9604;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff90c1e9b692ee8f453168448e66e1e02fab6531629322372d2f99be5fdd3ab5e403f2f300f190883416cc22c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda544469925af2c135b0dbe819de35d14571d48c156d0961b2b333d385c50c41960846c209cb459b2c913ca431;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8869271219072c610920df724510d320aac6dfeec0feb1c61dd5f9ba77e1cac417b7d9efdaa968d21b3f9146e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19908e3dfcfc34999cc63557ac4c041948ae45f09b3165f4c462a45ff44efe776653a5a37363f173f5097bbc054;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a57ef954c649fd2c16f8e4e112456cdec01463f73d326152dd3e080d0600744ef250cb15623330cec097b76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44b3cfe8f169568f26635f2e6ee650615a09ac081b101c8006331a4a5a0726353946ceabab08a2181ed52471c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189c77ba4caf5d6dac0df6b8f683989deb521540bab1a3685f355afae4a10923566c2d8871324c0ba9ecc6bff38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51a6612dc6038c01b367740ae8a3e4909471d7056ace5743f68c1d652e00fa2dd241da98b6d70a0e4482308004;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4a47cfb0433ec8c4899cba32bbe0ca2b884b8ac7066538b6c07a958cd9240f5c5e1d4c8c6273e20ba04917bf3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a5c4cd1905459bd443691704ad8eb7914b8c2fb20f848a56c190964052cd6c9dc04357a5a0a2d26292e118b92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h766449c0c2838a51986654b4091e3f7c41cc9cd2d54fea9ec465fcd186db9daf100f5960a7621510c497ddfa7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9ea854aea1001179a14ac4c3bb4c08989ef1c8791f449eacab00e9eac3b7477d73fad7bea6ca15eca00f8d40c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174cbcef78cf3852cbb066bd1ebc7ba2a62c879e69d2867039cd457ab8eef7dc062baf9a3fa31c899268c04b592;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bd22e011ff279fd78d3e8decc706372b915075a28db04315e5c9b702feae3816039ef55441024548bf413cec0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1456ba0742bc6289fa5f4a44e813c908fc0c0c8233af4ccfc1a3da7da115437439c80075fb94d21ecc09ac6b38c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7bf88713e686cb3856b3eed9b73d97673678cee95c4f857d9622c08e2d369aef17a623d7c9af88d934c042072;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bed8ae6bb7803e86fffe02bcba86467bd0855d4bb4a9fdb4298a51b92c239b6c475a1ffe8b32b45fe1bc7775c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8cdf49a465f52b257ec82a98b24f1436ee4f606ffe421fbd8811f79ff0c873c4585512c230cce50daf2390c95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127e978dd2814dbea2405febcdec982ddcdbb640b27071b3aa3403fc3706f9ba993aa6e5001b805ab7ff6d47f09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb42d7c0121829101732486fc313407209b0c19f045051c0492652cea6fc65998fcad0225dc6860cec54855862;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c90c595de87324bc2ed2c2c88fd716cc37d4e24e77e7feb1a7fff66afc8cebaeb4509ec547a2604c4fcb07d5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb0df7952a855d3fde603a507549d4dc3e41f04a81731472436df27101dfd91eff111c97764d0aa2925cc577fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c49bcd9a7356d2721736491da754ebac8b128840396fca3cedf481bc311ccf79e0f75e06bf167eb77934432c4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188d72786be6f3b97457fd3e7c924974ea36d2c0e72115dd7b6b9c495732a16f1deedf60862970ad00732f93e97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5a5f7d814ee8135724817f2895edf94f867745a7a136fc5fdd5245809c8313c93b06749efddbd920c8a1a3622;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc532c163e4efc7f14d9e699314f6973f6b2e58b9c7fe4c24b3ca56121acda5988c5781605118fd2d55f3d4b9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf41d60133ae88cddb5e3784c1dc57852c650580ccd0ee699b02f73dd3cc7f915935a5ab4ff426dddfbedf22708;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hedc5ec7f79723cb5c9a9bd11b29208e1ab360f41f4c9162617fea4ab829ecb163f72e952129629ac6b0346a85a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135856ea5fea5f19b4a453eb17e59e148e6e7f8ba80ca4f08044aaa55adcaaafedac26e2f94a69ec4eb6e97739d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4059fe3281042eb27238c022e44335f23b713b5a54d6503b82f513edb0a838436c52db6748b83d4cec10ecc86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab94aa36a33d2ecca41d7b722573ce7e733463d819ed6746db5afe0da4e9c5144309f6010b8b05c3aade594a80;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1258410663872b1a2dde214b368b55ef0aeb0f61e4beb7533486fb303a616cde22e149ed21a48e051cab7d43e53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14247ee8d715359da07825d148c773860ca9780fececb262ea9b6c1953e9597c37380e7bf15340f41eec6bc6dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1193301c788a64607891e19c9dc7e8a4584df37fd860d986228ab8da6e19592e878f1d96faa2b99455b546f4f6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d05c3b017f25919fa989ea9a19e94fa96a2a8102c3c66e4b6008d9e0d33521c4a251a36c8d91404ed8b2c0e11;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2d061000b8177e6fce5de01dc4b83b039890369a19333ab1a66c66f9e339bb2a1a289d50ccca60fd324b4799c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb764d0de3e2f3824148ff041c8d7dd901cd11d9e63ffd7aeda72facdea9387539aa70ce6129d2c64e60c19acd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c4de44b86a15dd965e6a71f51c0f3932d0669fc46330b824e3596ee347a766a2bbd9988a5f6dcfec6b3fa716a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h139c19a1c32e1abe6f14fce77bebbc5e2e3e0cefeabc96306f977ffd41f1beb532f6b7e0f1e408852a960621020;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65d7ed8867de6c667c7bb68c7445c0403e81602fad4d11fc3b77031bae4863f844b3061204c8b6073803a327b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ca031d0637bdf23fac35906c646a2f750a90b271c5d838797cab36dd18c09a9d96c5b0a31800eae13cffa6ee7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132e2eb41ba73a5167406a8dbe680be4d451fa216760f63e89eba672c13465371e2fddb9c99b53e378af1f8cbec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17675b50af8ea997c5d756ccb79f88863338237035ec9b3cc7aeeb4920c213d0dfd3f893b31e19ffcd294778b89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b45d013c297c0bcb3553c8a64715801f42e9ec0c9b91c4d1f27d00bb8c846866959f335a4e138ec09df7cfb8ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf079bba99b450aed4de6e4ef607211c97a65b6c52ea292393d6f6d13e9c1c91c44e6f48a97c39b20d0a43d0529;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6dc324f870cc1867e5686d683c6731f2b6b0b7cb9725205e9b1fcbbe91f46d3755f4bf5b62bf2402feeb525b3f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15116782ce6b53bf02a48ced9ef89d26eeaf1022da917a689f6334d6206336b38b3d6de72507c84b80212fcae8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf6612ce91069905c7c768dc79270ec4251c7e8b397ac4921fdaf42507b6df820c82b790eb8a86cd3bced79e74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d664d0105a9ca2b2720aaba457cfc7131926cc8237d432a4016519fe2bfb81a550b52764bfd702bbb179fd4de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5f0a2d51b581a1b792d58f3d17f1290edbab2e8ebb83316ca065721154e828bb1a4b66b77ab4580f6b60c1f55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6e015ef0039ed8990f421b891ac7be9af97a9ca2ce16d19fbba8ad327328ed31e693a5bb52ef658c39bb8c58a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h585fcaa7879842e067a509a746020fa8e3b2049c91fad319e3fe2bd118a2f951867a93ccacd821d224d171886c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74e2e9b814bb410e3cc2dbacfb21b7936cd63745a823c9c9f3c328db3cddb62f7de32d15f5cc22c4789949cc6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe7d0e98d6a604f6e293fa018fea7d81246a2f81c95f54cf24268231c2de56f878e05fb46b0fc208a691281d40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b7de1013c0e82639ab9c02b89b14b6bcc56a3fc52130f128cc8ae5d0a064c55e1b04447f420a17013c020a0ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f631f0ffc11d3892bfbdadbd57e7cc0de54593729f6f68ca8680843ff8158401d4a5b316f19247f121377c4370;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1839b3fc1886656b26dc93420b4cd321229a4fb665c184dcff3ca6de5df9b39df3cb7bcef57571f685b566591c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a3aee23f7423c9d38f5250eda7a4f8eda3f80b877ab039cb40384c0cd470e565808f224e5d6761edd6beae026;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ed02170a7d9efa8ea70d72063ec1910d80149dcf464ef1fddc80ab5a43acaa10c5e7323be01163971c7fb8358;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74698551fc33906c1936e927357490ba6addd6f9f1a623484a120bcebd412d49ef9cf85627dcbdbe278f0d0ef2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a563cb3ced20542f70f579ac10eb5a077915fe4bfdb8ee4e680853d964338fe95aedad9c487441e6de4db8e55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11dd48edce382c0314b1ba4ff725f212236733df30e1ee91e78fc33d5d15e91e6c5ce74672159b0a571a1ab8f8b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha489017aefb0c64129394858b6a6eeaa634a1e86f32df1607ae0bf032c2fe4e262cfbaff5cbc0f8164d6129648;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182fa9ef3b8c026a60db16c7dbd21eec4c93bc5c45639f71d508cd6ae4ce815eaf311b795d42557e08f44d507e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf9391e859663cd1a8c2166e7bdcae31b4aedf8ea07248b224c1896174754c3bcb8f9b5d7796c4c1bd4395495b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha65253bf7d0f8e9ed9b7e01c7394fafa0e90eabc426804234079874542f0ccb95d3702e95b100ce0f5e51e4674;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1980f2a22375b443461dcb5b65a4c034bb8d1708f0ca226618d2c41174bd1b331d67bece3edb7400e3be929d197;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6dacaef1a6751ea6829057aa29c0eea99d9e7bc48d397e0a6a67106ac48a4902a67a648c70e3f9c45b102b7959;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e08a0a04593365910fb7282d59ebd77c7083d02524fcc89264e01b6cf128e7d70c87d7639186fef19be2da71b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e0c1d5655976316500b7167f38d448a2d7bae685071fca9ec70b10f2d66d734cba90d09093a661d5b48b626ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6f3d6eccdf82191adfbf0a5b00bc99dd275a013d3ded56a3685eedd91dca8d8e460b69c2bec188b913445ec1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105a52bf0481e58e17256dec27a99b6c4b67309f49f8a83aed0bcbb835bca5391f310112eced80ddeac4b289c3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5e83451e11b734807d0d7202c7bdc98d15f30b45415a791a080293abb614ada2e205aa977302fa9550d8f26a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ba2788d3599d04a95ba7387bbcd460a6d510c361e8f6304a780509ab4520b64ceecded5ff46e62b8fd4e81b02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119180111f53ddac63e65c034b511c66c5cf804d0c6ef9eee507acc9b75cb5e1f684f84b1925341f53472911b3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f0d2dfe6c67b78bba2fe6cd87c2b4f7d87a36a33c220389ca8144700595117714229de7b102160d2ec7876152;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16265fd4ab17ba478b8cfe5290aa49725f54cc3b03a132dd9a1100f259d43490143c9a5fb58310070093d160e3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d50789f4303c87c3c3fdac784f9b1a902af0b6f6d3a02c3e2557da58b8fe443fa4f82b0beeced8a1651b3789c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be2b68e30328b0e8fa02366a4057410dcba354a591f24a50d972d14eba4183df9e2059ace972df6dac88245cf7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3137c748b02f50536bd0669544d4419579eb533cc89c08e9806a0f629f97ba74690b25bec9a71c0d8afa0f384c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80122218a72a29d5027530ecd9a9bf935a01c673b7906b842f7b3fe28750af69a6daebab6bff99ce12642ba18e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a431b9b8716b1b71c42765c747861a0dbed8d9543d36644c897f30b3e97dbf5ecbac08c49102b7c9a47fad304;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf7ae46c197ead851fe464e6a29225799210b2de912329b229810e307eff5d574df17b2f1fde0bd6d99df2b0be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c7b04f9aff146b66ae9eb62194a24c28e29e8469e980568a4f7b141c2c7daa5a27eadd2cd70b3b28a8e880024;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f41894b48044dcb32c80b6190b8e9a46697ae7c34460c0a6173ca1d6603b11628935620b8ddbd406f13ef69264;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fcfe76616963101384650965baf2f15a31139924dc2e8d0a26131d826a2a6bb9e7b7393f7408a06b9f8056d50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd113e844654ae86660f4b588f6e13a1af39f744dc74acad66a25333a1def843e9b1b220053dcf318745168ec9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haefde3f374cb4cc3e12c144693e7b7938dfd60bb8215a5bd7ef8bd012995cb5d5bdfbb62620d3c31f5f5aa463e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1debdbf7d54d9475dbbd12d2e3d24ab11ce44d2fb11c8c8e5919ec98c7c7e27cbefd5813aca9281b32603ec4893;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5dfccd3683d4057f411a43e770851e547fc347161f3d184237667634fe13e95ee079f11bc3861e5cc01a16f5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f7698e4a138f4d3b115630fe3f06adc9ca6151c6c608708dafdc403ab802f7d1accee37c2ab6c21fccc6deabb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcad7984ca97d7fe4c06144d86d00f35ea7478a9acdc527c8532cc58f230b7ed15c7b77feca5adbfe96cedfa5d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3091922fc30af66f1adf07613e3ecedd461e7ebe6bd3b33968e1d01c23fb0b6933d4a5578aaf891558567154d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c19cf11ad50d2aa790345f40d361334b89792dad48d9e2e4df1aca855815f99dd0d29446ced00798941589180;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b631d0d0e656a16c0d6672965dd2aa5615fd4c20e0c73bec64929f4474047bf77ae3ffaa2ae9253ab3d198b43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cbc5b1a1cc1b1795000c2dfac359b94260eaadf7e77a9c6f43dc6a4ff80581eaf7f7f5461640b4ffe0ec25d24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18729ca198ee34c51b36f6ca117619132f2e78c93c44e3b4bf20e01b2d07b1fa2bf8d590a71ec015a38c8e11e32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fec5f8978b0a27e6332bbd658005839a09d9e18f8041185891dbf838e7ca9b6170aab1bffccac9fc1aa8c36120;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha40f2748630ccefa728b83fbdfe62a8d38a41cf681105c8fd846d4ae893fb9ffa10920de6cadc882fe260d1fa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b25e074383bc020ad86f5bbb25d4fa592bef851a1733d53f1d50f9dc41dee435a6524140b09c85e03bed0ed7e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc53766c9435efd12543d252c7ef35194aeed258994ce2a8194fdc6bf058a9f8fcc88514b3aee3f29cea305c24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0e211f34048f5ba50ae07c088295b9e045a416e19d22f9a62e3825a13d9ca1cf564b11dfae30a0069c4935ddf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d85d3262065ca226dbc44a6ababbaeee054b5d75a43fdf96ab7dc51302e612874cc35f0e949698b83b66ccd75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dab1c2868a01813fff0632b9eadb25b9114ad4ed9de90e4ef29b04050bdb579569233572bcda61d858e7166c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d6c43a48481d9447c05c621d60d15789e197701f64e5c3ba600cb7b7549675bb2effa343120928afc8ccb4da7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e0b38eab8ad94732055ae441867967dca2ea2387d5960edce56ae09a10694846127a5b5a302d489a8652e4929;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46e996caa78868114acfc6cb3315534ef720f85f2c4a0daf064f4b9802caaffe35b3110ac324af3afafbaa839f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1c250008e62f34af9f5e18025a4c1744eae32ae19fee13632e8a922f3eb48ab87167d6d23dbe2a4ca33c349b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3614190f2c84109653e9391bc3668d6165e330d69d4f9e5e263de0caff721a8cfea611845a1df25fe2d79faa67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cf08e1fd6b32c45d25aa62aadc6b65083d369dc105e8bc1d870a3b7f1f151b44400feab6d48a8cd580a958aa5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcaaa0d7151af7cca9faa0ab02b5bd08c21f0b850e196a4c59c8a62172f3dce04ad21a91e917555c4bade3be0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114a1b0093e6de2fa8b1b371234efaf915ae5b731b5ad0199f26689cc10fa963e881e15a761590378ec4080d658;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3efa9ffe3b68d0e292d2fc41059e16da768b55708ea70ddce0160a669bdfb0250186d80bd4dfa321355e42d83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52d4a5622f928ec255da478f3f48591850e7dd32ccff5881653813634a20e951898f6988e42c702652ae8913f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e54a0bcb625b6703911b0a1b2c454f2295f13f705fc3d0dad3e49aad1a4df12c281d005cf168c128250745eab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16756d5f13aa7521d550526828416f7db999e875e4b1cffa9b130a5efc631dc5e59d5a9a32a1f7b26ddad1f0596;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f7bec614d319be20355089cf603e365aafa0f01dce7497d74271d5fb247328b3b648efcb217d6ff5fbf29a2c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15273ac654bb6dc4d39072d4bb2afa7d346a927c245796f12d59242db423f0966358da2418ecacfb55a9a6ccba3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db440660dc4b449d8ed7038332f387c3f97bfaab88fd60f88479b11d3407df88c662ff56269686345414a9fabc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc483173104f6e53d92eb77b025a13a09f68f3158a250358779f793edc68935a922b632cbf5d36bf63630871e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ece869010f226ee8b00e0dd5feb77164b7bf188b6e7f830b15ec7535c2c16f5cfb2e26e257839dc01d337f511;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h942ab7bbbac535d61399fcf33749584bbbd4754d135e9470ae066028108274d11dcd6fef17e9e7453bcbc9f6aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ce0ab40a540df58f1f45b5d089f1bb1013838a7e85706745fe92a3294dc09979b8739009c826aa5ebae3d4016;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e9993620ef4afd5753d96e77ac187183d54d97134c5b9f667c71ee0a85586479625e0e6b57ac5339834f7943;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c23ed5ac61214f8af114b3358ce4a3e6ad75602aafffef38f9c355e6b4b931c3e00be0640c40d70941a659c0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c350478c4cae0f54e436f5e662cab43712b07e7b2d80de6ede9d95487a922b49a94620140443da938231ff2bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103f0953a3642bc1be7e02fbade993a16d5e854ef8c81ba63e2a25408448031fad1458c9ce161eed5f05cca1104;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4372bc493e41cd6576b6305a908c8b0b97f48b90c2cfe3dc5239e3ff96ba2f9fe75c4c709ea84715ebbf4cceb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fe584a990cf221ffa2d86c16abf9f9913b0ede4d4af4f492250aa73ee334871f8c403e9936247064d6df1d121;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5420317d438278444e8052353a431ec508855d8fec14529859530a7d0827c7232456645676703e6c9d0d7566af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha17526584aec1d2d0046a93118d68a42c738a4c821696666ea74b6dc5f93d02ca72ba95d7a1edc4bbcdcc28de6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h409ff38f7fcf6998fc6c9b5dd1de2800aefa13372c1fc148c3c94ff7302497b09f5e17bbdb1702b74e8951ce2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159597ff8a995d3eb7220753bdbb8747cbc823eff270c20bd3fe604102cd3432466f6d9dc3c656e8470491342f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66676510c76d89f2186b019835f8821986f88d8311a090361f2dc7336c006f875fdaff1f3b1e5b57cc729212bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd02e93085fab81ca5e156d5837566d6a183a6faa5c0ee35d7f2419c54cbc16bb84c39e840b158777df66b9d12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1120e61c7674db7d634d418cd6534fe5924e74cea8f05d0c6f89df5480f48b450582148f09410222428710b2efe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca9e693aa3287cb05556d0209f339f85833dd9c75f2b7af1c8c0d3f966e7fe2a00116abda76080a7015255ad12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4762309ef2fdb320322e03ca41d15d8209e9c8b7fc0348f1aa6e34348274234ff4841f8cda2fd6a79578b8300;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e486633ea087ab84a5cdd4872a6512aa34e1abdc30798c456c3f69358c57a65a838d08ef839adb87c4cbe2ae29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f8f7cb27e32b4f9350cf91eef43dd171a0c6bfdc38b887525c590525fd33b788d0749541e2d29b9d7b0008b55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0a348519d7a550844d23d8230725b591816002c967cd7099e4b4751452fcdbb90c29fa94c6e53cb848ea815b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ab2547a83262924dfec3ed7b4f66a92f16953c77c41ecebfc7ba19411fb33f3642279182559a282f34aa10090;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45a8184530b21a46c2df2c9e6141ccb67cf846108c7baadb8bee00797a4436880386e00d5634dc0cd5e92d1801;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ab42242ed453bc786b8e21900d934b59a8fcbbd0d5e55087636cb327f0920f3acc89c93ebdee401cbcc5624de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha853eadf37416cf8ecb6846223cd72b7e02df5a89d12c0f38bf5a1d66c7e2d1ad829c5411c1202178ebb6f1924;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176a472b03f2cec02c44538413ab164da7fdcc68ed64693b390770c02fa2dae0fe432837e6a781a059cf3176b8d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7faa4fef74d4dea3cb2a7999b819e5d705099c968e52ceae1f079ebdfe9f268a8e03ba041e091a9c1d6a0b9cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbce0a0eadf6d2cc2307d37ab8b13c05407df1b3d465306c8f447c1d7649029353f38de5ba19705b883c094c5e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b0b41bce07914809d1780468518b76a160200dd814f9f95dd0a6bfd0b9f9615558f58b8409d8038c68d5d40bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c645d2603f36f1950907044e748bbb0d3413d22339db91a5e248467bf5bc966e7007af107fe84255295f3a8d23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a182645073d88e3c4c36d4647440f179cc8ab3fdad059ca263e41b7740609a7bd581a1a0d07277f56654c5ab9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd25b4e25dc6b9a52de773936f3e7414335fb3caa83a4b32f990fe112d034c6c3ad2e77461f8da59eac10ce5928;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c7056e894be8d8559f3889c8508fb10a23dca12d295c469b538a90ba46c227bd516811e815438920f0b415699;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75a0f42bc6d7012fc22253b458e878726397a2d7a6a7cf8d6f087dbbeba8e8bd49247327e4ea943e33ba582f2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cec6246a2430295fce31e05b7e2048a61dd5c51e5fc2c0b49b0cad246e0f1f1fb0c2c28016bbe5396aedd30ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b4a247625fa4be17ec25f2f7b45ec4c2a320b85ccf20ce619ec439a6146cf4ead02aef7a4201f000d1b436429;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5310920e2ca9cce564f4a54e5126f80a4865e1f04e75d48c7960661570c3b2cd5e037aa38ac9f3bd1b9460de3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b647ceaa60893e6be0eba3fda130a271ab20b8368f66242fa2174d026f8ade3025526f504b2ff8020e1dd4f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b73feae55341c449dfc9ea056434d624c4f38d1e6d55e38d8a344899214c54909604f8323dc5b4adbc826926a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba555c3d44b6e1870a157962ea0088f05c44010f0c10ba443da00517a024b0e6d60743e559e3680b34fbb6656d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16eeef7f68b939a2eb611e4c20127dc75713fa18210ebd1ebcf36d25badbaaabcdae2f10cbdd72fd206d5b70b57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5507449411c7dd41f634134c6cde067bdabc863d4d5bcc2a77808c818a8eabda86ef5d1a4819fa555ee32c6a55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b2460055056d449ee6e7998f8ac72743b347221febf7950fcd0b8970ea67be928935a83654845f82dac5c0e63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164c3aec6eaa7661d61f1da6a76a8393289af66ab514640b70b7291bd6478f70e0f84a917fd4c65d995d08c9428;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0ce10be3c811c3233e4a5b80039eb599563e3eafaebd8158e2baf5dc399a849e3f598157ecf61a8ecb9ec98d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d6fcaf12ed450c0ecb3d2d35f87915d5710959bd49ef5bb84287e507bb9464b67eeb9377fb95ef07eeaf7de30;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb51c83435c1e907676036c4d9851feecf98d6311118ebfd371c490791305a813302bcca0e2188b02a912efa3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e673cd49abfedde9955cc8c6b5cb0154a49f286048c70128a24e72cd23ed660ab91ebf063ddafec3a16305c059;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1270cf2838615b6f139e2b282d84609bcd4f150896af1c22c833ebf7e149018f7e1d7fdee261a7b66d52de386d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc495244f1a47da3fe1729c2b57c328de41c5c870da7095c3f20173d721dbd7c051648b3738003088fe5577a882;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f60d403defa798a104005a691fe11ae2c18a341501886bcf023412f1c4408911e88aded014425c240619d31d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cef333b2595d247fb544e7d98d490a674334af71cc751738567e4063ded19b07f2015f7e8949250be251fb4b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe5b689691060e0d439dc9fe8bf099c01af24eb795061d6eb10c7861e347f85c665f4caa60a7a7d45e22c223be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cca953987efe38d2257c262de417e4fb07b796fc6ea2d3b95779932584b7e6197252c52727c6ee40b71c47cbb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1941df69252f5ac9e7122d5a585b8bd911c92e5095983fe1e13c09b80bd944b4e8659140ebde8c6673c7f5b8d9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ebd33914326565c5972c071cbb1dd8af0803122230742017188a52e66751fce0a572b1c34bd00ddf582c82843;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4c16e8b408d2d1508509e087e3dc70c8dae34684928c12a8da890d26d50618d96c7a68adb9d58fbe14dc05ab4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112aa7bde16fcace1516ab996cd88f29ad660b50bc021773e5cf8f9b55a55022eef159b4370afc72e9f179693cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198f1f780c6f8d0df536b0816486359a46eaa8f6c03df40def44a883898f24663b33797437b051d316916b3c14d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cdd8231bd55782421bfcc4275112687bffdeafc34d0b9b3d2c77095170eff1f1b07d8a24fd95a0d1686ce2e669;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6461c8566c072f7fd2e03ac9ef2950455880b6e2dcc8a3672173410e76e84c64dc9b417b9abb2ae4a5979c7269;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19fe2b87b9dd98e9f88623cb7bdcdf2194ae1d2c1260ca3061369f8f16bdec56e0956ec3585f59197c552938489;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha510fd36a37a42ec7d7411a54a06337c6b2b573b16a87f5eae00816c51ac0161d7de5522b108583bf99ab2dd87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc4f74d8cfda49febc1e79ca4484eb471001b21f3d609104cd4dbcf45aa46fd35d98a9eb1115b1805c45976247;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94365d345af25f57b2b864c710a851c374f794e485609a93c60b37f0cb973d3a4a399056ba4bf36f00cc9da7f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15971537c18c3f7f12a8da845ff8e2095289bbe94259f349ecf6ad46e8bb08410dd07e6f60cfad1d9d2fc54a523;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7fc95e146536282cf9896b5217c34b81a5e85ea69298e96160a2d6f6de20cc63afa39374ae5e3462c0cd45566;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h797fa1d01440d8dfd7d30251ad33907867b0a1e8c28569a8eec675d7a647fb83ebd9af58adbd869d3baa3716a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45a9d1d6b5e058a9e32409f37dd71b5ff3a351278298a69fd3d1ba1b1394e98d5bac5c33d89fcd52cda0e7f648;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bb5285bc3a2d5d9ecedd3583c718cb9c09818ee397878635f8bc046d1abd54b73347157450613e3000f03ae79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b06a28447761ce31a53cab57731c02e019a6957df3e12186fda87121532fc5d40910b70cdccf3419d70bafac3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24296084b2afec9b7b1e412646a17aac1d86c7368a6ef54eed25d548c40ffbbc4f8e672af5192dda9f4932d621;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha69c1873fbea9d7d421bdfb3239778845801d5441860f46824991c8af4259563f13a888081fe5037595b263fcf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b0b102b71cb78d2808c75c661148d2d3b96862489e4f969e65ad72f239e8e6d46699765297b3a6a71b4a86607;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1215d46a522097a76a0e9c1dc2905a3083d9d957a849274f65ad7e18afa4b0718f3ef3505dd7e1d428bebd84440;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11455908ea343a15dd2da2ee9b12c7203f0738a04ea58bc40805a2501c10abfd8285b05cb7409ddd5ff364af996;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hacecb7bb8b214b1b437fd460ea56998132b1cae26c3602f8286770d980ac783a8ccb4c8f9bb1cdb1e81f6cfabd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1442a4d3373f4e9e8f2df33f364812031c580f2b672b808aaa4cf6ce42ddd7b9e5146286d849a3cd06c193f620a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dbefcc6d21c74f1ac9b9332eef54a9e4646874e77b221af43e284c61e329de9f07011018485d23c27c062e9c06;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11338972c6abc0c8c22dfb697269b63d6c64b64303809f304c0c9f37a38f1de2e51e5ae9b4d0947d53bb77b1f61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfee5c80732a9fc5d1f22781e455f36c634a0dd2f58cbd4b21e96f2379f60d4eaea9fbf943bb46531841b5d9caa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he323bf1bba0551178a026b55d4ab943fb6a316b12ed13efa5ac351f0ec468bfbb81b4910bf01e97ae9c41f66d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37d376cac4768f2c4e395d01e474da5f148bc17cdffab91643b5a2b8bfdb6cf5126136ee454e072d11abbb67d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1522f0b4928906b07b0d1248e776ade4c0769e8c1a5e6a899033ee2e9bf6be730e2b9a3ae04e00c19e59a975621;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfacb1942dc3f1aa99a1dbd9c3fdcfa20fd9b67f75d694d72cfd5e9a4aca790d341d49553ced39866bc22d2dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he84c98d9c64db36966641e07fae4ff587935a33931c6dd72c9e90f980ffb6b1710c6c2ee8364254be0580d2189;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1513c60945c89694ef85c1a7abf1c0d427064cf7159756e56ee55d0a88b651a957e988c4fbf7cee6623ae3ed58f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78de496087d2b3bce14299d47247bdc79d02423179c9d733bdb067ff5892db5420d9c14755feea440e68e1a829;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6cbca4bff5cb623857839ca12f9de8a8ccbcb5157dd6d0300fcc4d6e8f119fedb8a1dc4871f1328a4dda79a03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha84f8fdb11817a765daddefe133fd4d8d3146d99d229c80122a0c71f229682b0a170c048ac7cb53e3f641a3896;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2b15a0bd5bb2e91200722562f4d2f7de6ccb6ef85e562176cab3f240179e83384086cf8fe4945db3af9f7c3ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f97dcf66ff1e388ccb22cbc710a38cb3fdd0a239e03609bc400824f708a41d2cbc2450f69bd4edeb80deb44567;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0a7d3e66a1698e567438bd96dbecd1912dc1f5cb360dbe40f9ce4242ac05ea4cfe446807672ea6bf6979c3745;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbb61ba857ed7b08e11dbc3f19f6daf38807c8ef60f2ae837d336e19c62bc067a4da4eee91f599d281a7ce01d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc00e12ff7eca40dacb0da6ffedfcdbbc78f41d3798a7845edf9c757907f4a1b03649a1043735a6f4981827efc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd555a555e31cebf73be57b7a33b5f7bee4902432dcf1d3ea01c11119162ea81e882a20172703f3703859b55715;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd800d30da14393bc61b983d97d8243f8df5bb659793054be861b2920f23cc48c9f5f818ec7326a226c8850a3f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64afc2c4e523131ae4d561bc35cb358b8e39344e4b8080edb35d8e92cb8f9330f6bd377dabd053a77b99f1cb6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166867c0f819e80fc1dfd751a6ae2ffcfe609a3cd7a4071872eb24f8c94095c2e71bed3e0756796f803a8d2b6d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8e0e0a4cf2468ae997bd7f4d6a1849fe61578d64e3ac13c2890b5e9cfa301a17690ce1b110d89cd754ef76bdc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb7ac2649ca3a91c2b47d39025ca2d02dbedbf30ae91844985b068759270d80dd5e18960af5e1fccf6e6470db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a2e24e32ec1e1127017780b13a022a52f4e7fb68af53004d7a270b97440760003f23faf26ee08a94048bf6796;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ee6a260f669f2135a2c23bddad00b367e834da5e2f5667a082a39191dfe7a633a4d09e5c71261cca255b4b49a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dee75c56b96070ac921f3df80518f551d56e6018d313f633da49be50392e8c20c52570d78bf0b6a562db9c68fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1282519e8da58a5dfd83c817ce5e2da92800e64e8317624d14db6940b564ff5a3f13ef2772a68adc64eee1ddc4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf2370dabf2906b30a4b42cca77186ab11b51cd97adfdabbebbeb857e5b17c99251b8007fd8acaf4140a316766;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119349bf41633578bf35088f59b7c5fd78ab1bbbdd3af716fcd8da692c7ab5474b67af4ee23dd7ddced1cd55ca9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c943e3871d09503e7880e71658eb05d2c135fa9cb73eb9cfd4c6963dacc5d20137d615d6251e51747d382c434c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a97e84bc345f31cc5dc053153835c20f89c2a821b88c24fa651253e5d786c549037924e6e0ed9734d8fd0a447;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4f8d621d7fb3b1bb3b52cbea21a7a6c562feb6f64014068788329feb693a910424333abfdcd98144b72b8727e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c951bc1a5770c5479ba07e4e21d8ec833289dd2ef788b8cbbcf3bcd28e16674af730dcecc5cdc2e33f8b7b48a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec4bbfa7140a5fbe7b1e39a6b369b6aedf09e39c24afb6bb60c588d4d0c0bad6fbaa25aba940eabebc168f68f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d26e673aec26bfe5b4e4fe140f5664cfb7a5ba2d642a14820d3dad071b21f57f37bc034dffae16e6b5f23b9e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184f6be29e78a1ac5d2607310d4f2af3b0db67412ed1b0358111007c0cf03a16792e8d0c91840ffa4b579713c8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f5ce44d2188a2650b2b399573166c6d712f5a28eb67be0f6eaf0e1b6eef5baaafc533ff1f2a925c331d305248;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha53c0aa0aa707f2e2b5958a3593857f0929f5040a8c9eeb1a95aa54a5b3184db43bb522943c97b959645aa593;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59dc2e611f95dfe26cfb46106db6ed58a91e769a0fe8d7808f2ca232a8ea961b9080c7eb102a76bee2d88ec507;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b73ccd6b0d4c75e0a40088d6dcac234c8e4509a4e43a7cbb7279d222a5b6416855a4bb2751eb806e2aad929a77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa6e60505dd01ef4226d760135e74dc05e30d9594888693928c7fed7943b51ce10fee028c39c5243e8e0658d21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c41593f8e789403d898b617c3ca8a8cb6e22296033bad59a3c44c630e5db7b4e098d1e8edd4d89f968fa8e711;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1594728b68148e48bc859da2dd09b03b1835fb9527707aedc55b031f416c28554507861c37df55720d3e1425319;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125b07d78aae037859997626a0920539278368ed060b398b1251b28a902731207ded11a823b92254b1cef39db6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143e71c42615d126e5d48a6f5db6858bd9096c0f59d030929a52de05f46b78f10a8cfd700c90e52043734c5c1e9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd4151db46044607be4da741b23670b5d67f78a02192f0903af9f2ff5c7d167d2cb76ca91cf7ac1520ce5b3b62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97505fef843ff8f13056b896f83ad9362c410f4a0244fc3b6750be23d194822c5424fff0cccf5879637bb5063a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e7d5c7a8dbc9d0ad5ab7f913d07aa94e7531f3ebebab10ab7bc4b4673faf4ec7db2c3750eb50f40938bf27b67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f0a26082bb1c070e581552d8f25656acc2c7fdd227c42a44924395bf6a9bfb982404ed2732ee4c133dadcedd2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbed9fe00138f919ed38eb80fda26ec2d1425cc100333c8c7564b62caa5a99aa2ca79fa59f79a38cbc0e0f1f660;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d41a09573818fa3c1f471e3080629c0b22904e8f7f5f87ceadb2c61bbb0f1b60975518ab4f7d4c3eda137dd0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c714be759dc814909cfed0263086fb44795e59cd51e1e2b1bbe68ced54f524d2c0ff2730548936c7a8374c8ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a64c9590ef1fc5b5a282edf0306d851e2d0dc0fe41d6c601298da5d0cc032690ca908c65183287829a0f8f7de3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88767bed25eb1d9040282d76204ab60f40f451e8af80faf95bd341b616d6c4544ea369e739e2e1386bf2377c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0a0c66c8e6139e0b13d52c976e17f7a5ce297a2793ae5e7f6362cecc897596a99b67fe38f8d901680baea17a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f5fd1b3521838c7b7bfcb18f4464e24b9fa035fb5085f0bf6dd9f56629cea0b9901d2f297ead734910940de97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160195089df96a138e0d3a828d3cd9a8cda3aaadf84857fe0224a125f235162bb9ca7782a41de96333a8b517583;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9720c0f2c738327e610d31f7b5701cb238ccda0c1057a11058ab8fcfcaa10efb9332c52c5b8aaac5d9469c71d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf8d62e9a3885c00bf39c86c9921ae15ffa86303ffc138237f74b0fbacefdac26e1b309ee9582c81527586f5a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10120beebc751445af780247c8ea4ff351a8b1516fdecbf337bbe025dd1ad22767d8aea98d365ba9c8467aab4ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6587bc7e992fe202ae315396adb6e04d290ca9c09bdada8d567723db55874ed24d326359eaf855a6dd69273b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b55dc059ad48f72d9e116eda709fe07cb3d4e3cfa1c677cf3113bba867cb6a2e6bad1c60d7790f77ca67bb2ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b74977130dbfad5678b7b88c0e0ca303de6e1b30af757d05ec83a372d8f2d278805f651663e8cd187348712a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed687914c67634bb0a5eaf94fbcca478c7ad514d54d69298542308c2bfc33c6c7e5f730ce49e07f7f7cf2219dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5837ec41aa82faaedfdee93ad299871c699f2f45758480accb36594b293131559519608741747187ad79a8c7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0e93b7235ce049277fe911611465ba77eb6d1af4a1473831bf2b2804de3bf278184ebe5b6501791908497c3d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a34dbd006d0d96b2ce23ed1501bc8dcbc2dee32c1f39d966fe3008abd9811e5c5fe4f2ff201ccbe39161b41d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbaf8df91f832aa3ee4d8ecbb78d229ce2b0d03de0ec2363de8e373843882e2a784901bffc74bfacac2cb6c8c7f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ad6649147a084b5073eb91bd88cf5d118c9d695b748623ef81816f8c25fa68dd86029f9770555ef9bc426cea9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h910d993f2fa76c285b9679080636a65fa4627c263ff69d99e625221478dee3bdd3aea29dca8c5c78197187ba2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33b672d3f5468cfb29476ef3dd3bd3ae77c09673fadfca043a4a6bc2778cc8af216fdadea2be2a0cbb6d74ff73;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5b67f9c8f5badd1f76cd3307ad092f6de783f15af03edc599d27813d893b49e78c210aa20448d33c872ebd337;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b199392ac1bed24a1e87d3ab08efd235655143837b644b5db2647b63bc531de81389e1ada093e34c0d68b00f35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f3ac6127a74321743386ee25ad8f201903a401a00430e79c161ed6b68b2891ae8dc4799860b9da44b403c5c2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2d56ee7fed8dec65e703b83dfd25335bde878b55ddf9fb4d1fbf5ba77e806d19f00122bcb81d3508ef7ea560;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0895153a73a29a1c54a402809381b87f7a7d4a4e6dc62070183242cd6ceffee020ccdea90a91bcef45a3e8973;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a5483884f3bbe640b7085aabdfc8c2902f1105b0444db669e70324f2453b2eff59efca8058d2739e2d2cf83aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4ff6e364639b633b8eee23c659b84cd0ae7d22fc6513220d360272e85393896d5c6d312d4214e3ad96d4f27f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5eff539abb7a73ede902273e55362b5a464cc324e77c39e3a413244399b3a89ee42361a229bc21931f719fd168;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1065fcd676b97fe600baf7a130a257ad83a90ce1df455aee6f84c8207f029e59140291f4da9e201ebb0f0e18d93;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18017271951ed38d938584e0bced2cb7073c7042fafc0ecf5e2996783408f9f98bf24051b9ad1231b4522c6aeae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1e435027452a761d3a68b093591f25a44eb2588f24e6aedb8d9e66bc449f6a9898f2ce3b51db28efa0d886bea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54ba706576f4e0f6255f65539ce70879acf67a45ee246a74fb26d7bc2a1ad60cae688f60e3056251d06ff32bb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbbecbaafd609ec0938a0e22f89bb20d953bb8569834d89d7b424869ac7de2830f4587fc471d3151c7ba5bd976;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd66952988699a08f0cc75dfaaa796c7ddae71d20a1bd23056257505e2c5c0bc09722e0e85a9a2dc05c14dff5a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2e200740d79f2cd4b4e2eed4c23dee1fef97e9f521e02b47ac3cd2b003a17618d79fc9cb4cded9a9e901157c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5f0545389e6b7b6bc6281ad4f6baee90e2dbe24d99d1faee59b55c24d8706c92bdb63b190a5ed47c53abf4514;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93fa4a5577023cafa9116b117f64b26db080abb5de1dade933f3e1db56b6e9ad520138550bb80aa5f75c244b3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d95b0608433b00d97b26ed6d2ab9c86ec3c1ffc6f6c54b5233970d8fda18fe086c421c0e7ac609e138ca39c14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b51dc3f90d54bc77f787699d0e904118f24da3694c488d4fd5929ead1e8c567fe31cbafe6bad77b91d9649f1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha05e327f2113e217fccd22ec87429898d80dcd016f81d25676e4fd2b33617b6eb247847e614f34937456686f98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc1c51f22462c51c4ddc3702c074a522506884057d3ee024d7e5c4bfdd93b719341acd4459a5e6b79ad9c62a49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1324414633c92aa06d0099d8f052c454e0df9f480be29858bdfa7e8220aa9b34a9f3014f7c55b7691483d241c72;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9dd94341c34b003358479b193e6eb536bab18fe33d86cc2e5f63a415fb0653e8967147e8adc87394cf5222c5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ebafe5ff2223e8d211459696d68237b70ea1d0f1e770cdf68c52902f30f35f19e4c2e81080530e49c50c734ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1152b2f21debecb92bcfecb0fd74ccf2c811ab943f040e4c65838b75867f8ce2c3b08dd417a952d8fbd1d855;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107b1a6d9eaf216af5ae82552655c58fc76f94e0267142881c4fd256c6c6a1175b26b55c6018992b04d17333cfa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125fbc8d9084b6f39b9b3442dbc9d374e31e88d0378b845ac7d831e6804f38a9cfb177a0b8e4052ca682493b36f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a501490400e8293c5b1b5b716d66e546eedb257afa4c42516f3fc449ce1d749980f330b6a27457dc62f50ce3ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164bfab72213355058282628e36f994e6921840eb75ad54ee54ee7a6014dd964f67fe796909a70b1e1ecc872d23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189031845acd0040cf79335274bbf16d84720a80ae720eeb7fb42f6579faac102283df9c5f4fe9f0acc59f699a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6fcfd0c1a89c9e6e7b4e7244066ac3fd5c19607d2402388083945b41b69bdee2c6cbd588c2c373753c8d3b2c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ade9341818970aa04165cd8b9ea1eb8832de41c151e141e5eb4269c26c92a94fe023d97d85e272d8b919a23f4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcfac04412066ac77fb6b34dbcb17935dc32b57cece36104f1e9616f93e51491055e50b503dcda7514c6283bff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ed1124b5abf58cf72a0d84d7ffdfe7166004a5f2b057c7428ad2c1faefd0c0a74584cc673a022feb533ecb851;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbc7e45a503d556858cec16289cee6a3bedb1b0c77623a73fd74b55fa6a1f78aaeba32a4d5bb028ec96ef02dce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49c74b792dde180c7e4f4997260b374b88375fc07f35515e47ff9cd121c602ad1a02f9ed0e00079f932d580576;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31962322fd0717912a1517b7750ed79344e7c50efe9896b760e47e7677dc2666c1f14f7090dd17c9a764a534bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca2707e9a0d62680b5d5462b2e8fb09d75aa7e90272ba780a205f85383667baf9b5e95b36b428c30445ee8d23e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5877d4efdb731c5e332f6a947772e55fd25f910a9d31de53e34de5446334a43f987f6e6921f9e21cb8a07ceaea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5286966241cff60b9d89bec27ffd694a881ca21d32f5bc72010781b88473f505a87a089cd7c98d54e3e7bd1567;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e15cb86efdb517308bec2b702bd10db1836e2aa93c497afc6f93e63bf6ff132cce93139551c4e9184e800c2b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd832d2b58f3f3ca40e8c1b79dd2ce307375b7ca356453ef13590a0596dcfc1b1d892302cd6ac7851ef46cf10c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3061d5a194726af800832788954d88980378a4041ebe1fbc977a0f5c6290d55121b008fac34393a7ca3409c2ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3a240a0bd1cfeb926a350f2ad4b507c1a23704c6fb6cd9651204ae8a0c20b09554ffa0c2165206305214e4dee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1811adb9d2cd8586588cff5ea9260063aa9670dfb70a1e8dd2c65159969b3a4bed628c7bc9b0d4e85efd023f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88f430b03d0f3fd69d1fb98bf163502633f4b4145d141499c267818f729f2ba5e363f2712e1a2a5b6724202973;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hded448abb196e8afefe2dab9860569c5e8c881913bde622dbdcaf52e5feff11ae9190c5123e3d1cf12c60cb0c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8df2d70f4de8ef760f8d8d049e9fa2de821ea78884df4feed50de21947ea5bb2962207096f21c5c579116b393;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc04e6ecdccb234bf5690ba19343dc217303bbe92a9309082ed74fe5400f3d6bb5c2e27c9ba296480657f98061;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f34eb72d4d97aa3d6c34a5d1563504b1c76a907fa4d2ca9890163c2cf6ce1c570aaeb3235d9adda548ec7e5fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha38849d784ee03aedc298b4a5b0f7048ca007cf172988cbc469eea17b3ded1ec3c5a04c78bd5cbf8c8d3d858d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd80035c6b7e03d7dbc1d45f1e852583a407718384d937103661328cb77a40ecea1290bf393f5609a6c0637438;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16de78b35ed99f1ea25c5eda02f6bbc62d2a7d52ae2f01d87a9dff9220b35b6025091361563fd411c3224c555f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf181f513ffc38facfe105a2278574f4fb422fa46fee2e70af9c59b2962c8610075a1a4b8f3b1c84537ea377339;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1483846a83d03e31d8f4f1d00c8598910d713208808ae13d0213cefab0941528f17f777f85c494df363b21ba667;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d112fb23edc18d4caf21c57f0da145046077a89e85dc3916f90f53cf201ea4ee13fe0a1acc6c346f59959f5e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba84803840f0577d685496e64ecc14c61fd4dbb57266881550ce97f392e4e2506b957fc255e9218d3d7cc18f29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e83317b908e4cb73c1acb5a4c3fdd4ed561efe5155c5d24a2cbddf48bccbadf0293b12bb1d3797403ca9a34cc7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128b4ed09ed828259ae30d91bface89e56de24ee3f73280ccdb772b6a7955655b1243fac171afcd6d596cff804e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df19630c79e12868d51334bb7d49458c37eb7b8467c73d0a0c85b24196d05d273706d2e72fa8d308d0fb05e5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cfedd7d0d7bc1ab9854b67d935330cad56d5ce99c4d7a70f74ca71c88c97cbdfafffd7e9a103c10b36650e006;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192bfc715cd70bd0e865061bb87441e3194ebe495b99cddc23074bdcc2b0da474668df82c53438b180c960488fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdfa7b418873d387d90bd045908ae873cd1bcd0a49c93146c1d7283ff2adc5eb1c7a0508b6d85e9fba0b56d8f21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4756381bfdd2d2e7a37b3ffa07013311332de192c03fa87db82b6f224342ca84f884523eb15464af62269a15a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18da0619b98ea1abad879b3049771ed6c3401de5c0acc5ea28b19892078ea20fbd75b4594a03b9ec574183ed5b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f407114b8db1394af686542a739c6ad91d66ab086f82b408e98ff486aa5b72daa6bfae4c8ec27bbcae246698d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h892ce7bb7fdd6283b41503b3f1a4b63ab81b5ebb3728e8dff739d3d1f117656abfe2337cd0cdb9a029e47939e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4bc7758fc7d5a302ab75cee395f373bb04cb4e6435b6a8335fcc22111ea978ba3917e154d0a0cd126bd7ca6596;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f26f66171f2c19546123b364485fdb0ddf197ef6e095d691afa2fe28aeeef0f738d497e5b880e27816709746a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1cc329c4b1cd7eb5838587fb10165d54b1b3034cbb3903f9739088ade33bc32a61f03f9c142e7ca23f50a606;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d81d5832aba90379f842ce572f4a3ec0f9ba9770b1eb46d905e4dca440a3abd9f1a6478f8d4c27ed7443988e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146dc5fdcc8b6d85b9aa50978d83a56a96d88d2e82d7ba30248541ef4fd3771b46cf8a053cb6f57a56eb1a5f8ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df7a51c6cdf16be470dba2b0d4ca27df53e089028f78f359f8c9e2fd00fc2f593aaf6b07f0f225880f0db48c5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a8ebdc1f56ffbe61bf963777d4b169585263debd54c85a11d204f2afe012e3655549eb196d1e373caad573b3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18899270b6046ef3771414e8c008db9f605e45da8e7d02560784403e64101b701c44726939d44df244221ebf97a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1670b4c9cf95f5a94a3eef05aff1e4af958cccc0307cf04c7ba95fc167dbaca6c9047665d322eec0dcd88597bb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3c2d9218dc8fecb7e8c9a484744293a0ca5b01d7e29afd0c5b09d2840dd4d2bca1a174e0247818a02066c3a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ff2b0953869531bdf572f47723031a7b39faa63a16005cebbcfa97bf8c5b2be07258fdcdae2f3b84c99c319e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b745bf80dbabba39178b79cb4078fb97bc5a5154d9725d11db9e4a05aaec73332c5d068d00a47b4406cd830ab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7064e8dc4ec2434c75c97de4cfeb27a11c183b196b64985d408e0567febf2c728d8be724d7b810d4b61b6d9581;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b5fb3f971be9954761e2d2ed62fe6b1e8837131ec4f13640b5cf4501d6f462192df40eb17de14714f012463ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae9abefec215a6adcaefdcbc8b7d12ff736f69b5bafd2f6500bcb8cd63c4edaeebbe5bb09f458a254441b33090;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9843cf98ef66ef8956efe881e1df17092727ff4144549507e0b8241d7a5ea62478b12e624968ee9342dcdee16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h675cc287d7cd3b49620cf348a82d3326032d3abc7c813a61ccc77ff701c00d03a49dfecc016498ae34eecd595e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5bf127edfce9ccd97cc9345b789d3bb5efc56aaa251bd0324ebba3249b5f9c9f6182ebe74f0c92eaf8df7dd03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f06c1737d5397056654f23ab58b1903d7854a4f2014112d32ae15009d8ab0abddf5597d1aad2de3976154e778e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ccc04f5a4e7401a9d227364410892eb7d74caa6451cb81d464fb9519bb0e7b32067c01cb0377cd4b52a331650;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5dfe32f9243847a6dad7179ac0a30487b549fb9aecf9247ea93b3be5ef5e6fcac31d909ec305243508c1ad82cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126d4fe6f440647e7a59d95e6e690258634bd10756603a7f2e55994e58730b1c5a34d03c3ec171d023edc44aeee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h795bddfa99744645119954b81b0f76c5a527ccbd4e19ff3d8f09d5260168b9e3104791631764d374732c454c9c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b2eb992957ec324055dd551e555390a4cd648312d893d47ba3484d2e1b518bcbb0f3fa3cbe1f4a198cb4b5561;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfdd03511cddc05777bc3cbb738f5ccdf78a9c737072189015ba0423c0ab68bd6df612a65556a83cb168311f98;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dcebcf90ada3a833acc022389495e63c107a85809ef5a6e82a974080967ea2bbc03ae4e8a60e6067310bda706;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e92256f0494df1e261fc24cfb876a64c310d465d50f99a2565b5e0882e58a92c4a63b1e0471d41245cccc635b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb587646dd409278a283b2d5802a362ed151c2d4ae75251c754de6bac4a0f869b8b2affae641a40fba8af80612b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c415967c488a21d05bd3792cb76a6e2920894fb1871eb88f8f1e2abd3a1d41765314a1afe2f95bf04cc5a44ae0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h562f71ef08d601cb4e3e097d9b443f70b09d90a3b227b4fa2def7bd08177845a09b9d61e6520e3a0a56d7abbee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9eeaf1d350f8f4018cd3500778dc3bc67706ba397db694e114e932db00026c3186a88d2883d538733f2fc3e35c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150b0875e559cea47bd4e61b4409e0b3162ae298030612c3ea7f7c56a2ec4d6fa21a06a08efcc3bc4495c21efd9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h786e29ce3afd9343f27aad82acb8707017dd1a3be45122f55a655aa8bd9e9da5187b4a91a07afce0a3b9e978c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19be206bdf8cfc7123808d05ec92f04dfdcee244f05cf60a25cf969217d37258cc04842797f4a53b7f06404fbe8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e8dfe4752155e361368c88d1a8b0c287faf965ec6aed7e6cc53228d317018ac392493d0ec6b8ce32f5739afc9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e990ad95dd710958a78a0ab88d5df6bee802986a87c96f7014afd8f8bc29e34c4214582f0105d0c4df36a8614;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbede49627f92c67b913a1f0dd8ae3b50031bad81a49a0c8c52a716ae78c07f30f75b0f85aedfdf2ab68f483ab6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19486745834d5835d170a09c77aebe4b6a1775db7dc5b3b5d7ffd3b4f3a6b3d524fc79262d0f7e9c6f5c329b66a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9abbda9281cc4105adcd8f26df7758114414540f06db3c1f722b8d299c2edcbd5601882e59fd23e79403d84f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1390637b4e45cb57c67f14d7dda112cb36c12b86d625506497c56212c6fe9961f6c946845d89a04fdf987b51a79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd45cc869004490ea6839afed3aceeb475dda02f024248449a5633dab507b56d0025c0fc8d3bf614b46c17eedaa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6b35a0aad6455f265590dd09520d410642a08987789505bbc5b3d1e0fed64b45c012a191aa9826b6ac9ed9c7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d6297b13319bf89f842defad74e3c0e4f6201f524b820a29ac80f3eeb1452beb6e148b4052f7a69c115e14046;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b7ea5cf8533fbc76d36c47b1d62ba5c3e8fe941ed213e474d3c8c83bafbc5062e1f86e5f2d42101a3d9d00399;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha62e381c251b0527c69e9b8c1f2657a5e1806aab4cc97913da291fa4d59e8e5e7a734ab437009cc6df457aae70;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a63d9c2713a4e161de1849673fabb40218ab08e3e2937ec2954e7fd965b8d88b177ece0e314174224a5069276;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14160155308a8e5240653ef47596b4e2ed57deb152a1e9b87b754161801d46ce5d1a342e66a91e47a589f40ea29;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he50ac5abbfe60eb4bb1063fcfd2ce67907ef7bdf9414f36187cd9411ffa531126dc890bc7a7c820f9da00fd5e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b996b805e9a3b301b8bd807226bfd3bc756b36f73fdbf35ff5d0b205f14c308a580c38bd68f1d4c40b011d351;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199f8cec45074be1b8ff61ebf5ae4fcc0ce4ab6eabe184c6448c2089bcfdb0f75e26ddca3357d89a7fa8bcbc62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8c5a8919622381ad3645c037329edd7a73f782817dc4301571b5b8f3a4220ade40718f8b7db72751b5bb822ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4f7ed3f325eca99f99e4716c440122ce4f242389b74a797078c0c421a4258734d63e0af20f4733d607874a24f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155f9172645e33397a26780a954ed5e238e84015cd2a4a37526c04a4c678f165aed378025ee64dd5fce0c2f0e96;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa2ca6aabbdfb595e3b674ac342305032caf7bede65abd7465561e3d1461327df6847e41edb65045966bb79eab;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14cf7ff54391f1f9cd99b49469a32263cbd87f62765600a8b3ffce4a652df209d47e342b01ac644b9ef828c8aa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1031e74b2f2e8094808f4a2a31a8a4e4fb7f965aff7c312c816affc9b4221dd124f4c76fde9877203d82337e23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1faace73645cfe68282cf77b0b4cd551364c32593bb1c684773e5ec5cdb0c74cebdd87e42a77f6d35626c97ecfb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d35f4a150967a8522c4f8cb65790d86e0bbf440ce609129d610a0a23e023472ec40c312a1b7fd61fe8c13042e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fee53fedfa54d5d58101aeee3da76a86dbd4ae8853586a8482e9798d5e73f6273e075b474abe792fbe80b6719;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141f27ab9169a28c25d6969ce9f8b8a023d2e6a1b6252440e684116f477a68298512ba593c552805a36023a3440;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c27281efd770fd24ac9e223902fdb4cd4c72953e11a0d943312a558e6bea554cfccacafd7ee1ec503e9139b6bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10706033ca36ab63bb7db6c7e48f3da4eff1f3a295bf99e13a3c84a7d8d775b35636961cd373bd7c2f3a61954cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11510a9bf7b14904eb5101d30a29aa579dec9bbf03bbb767dde36ce65b4abb883e792159132b1cb1f4596941952;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1084118ac6cee01c18b654058a3ce4a32ea7aee6355880b4ce9ce5201af1c7927c6d5b6262cd7dc6cafb1fc5666;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140e8018de2782a71d6f660a9bddd7eddbdd2903c6fbd54234b852295b4f0ac2b8e9cc1a2f2309fb6f124c44196;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he951fd64b4c2650b1a661fcf6c80328243c86c3be5da15f2d93bffdaf782e24b86a0fb5deae1d72972128f05b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf725b763ecfb6908ec41ac32dfbc443e37681fab4867e2068617739d3c6f649f984d0ec3d52e2b96f5d8ff22ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10123d8ebf57e83fa2559ee2a0e90d282c02f16688aacf9a88216492450d61b301589d431581c29917acfbec8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda9815f4daf7678f2f40d25453e41be62e430e6929d63db7be8c8a8555ca73b19645fbed4ffc21b380a34c7424;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5cf8491975691274c285b549b9510a7b7f73dd58efea153e3e5a4b26df0fdb80a5ce5f9ceaf1b048110d81724;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81ad6465deb940cee409f08934ecaa3951fb073bed1421d2a7375cc5d2390de7c9c7a01ffa0e777238bfc7ef5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab883cbb3abc45117f0d12817baa26704f0e59bc67183d629553512ba746717ebe42beeba9f0708f2aaa1c2a86;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf0d1022e4b266aec0453b58d5a33b0f0e8d8a8a3028923d1ecda9734fe86989dff5bac5535c657cf30ca8115f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dcad25203afcf0e3b626e9989105761c750b5f1dd77b94686b6ecce109ddf907e012438172db4674fc40f5187d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1973b41c4898d97af0d6c316d54feb91a0decf637d48539900936d842bbb5f7dc966a37d220ba2d5f46e1afe0a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15cba771f04f8b27c823cd86790451be9cb065eb95392173d66706277a396cda3eb5cb5f2ddd52139b81baa560b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb45ae064b3d112669c03f15d178eabafb2c7bebb0703c560d65111c7b087bd0a127f3dcf4010694e6fe3863c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137e3545aeb82466519e2c3525fcd342898ed4a3abfc8692a7c4392e640f1a37e5d3c76ff0a810e7cd4f58d6e77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127bc33bcfc5d6b255db376efa2bdbbcc9b7c6343d084fad1e7523f0e577ac5ec1236cd6f15ae3f7e45aa1d368a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c070178885e63cd326a43f89e0d11e43777c47957bb9d6275b194e1ec90ce4081f24961afe2301cbf9bf32a12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99aa40b68d9754b367bc673f43fa649714d5a0cc30ebff61d011129fab0c1724f7a0bc1b415517c698650addbd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99e26b1c455a694d441d1e7df9b0c93e4085f452fd03a91151f57b02e18bbf91b19146beac20a381193c4e4a9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0c68f1cec9b245efc9bf6c8144ab74d4f7e184cbf24cf8c974d9423539a2fdc38a593cd529365d326660a9e35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10aaf121156e09410347005125208a6cf339b626819c248499ffea591a17b536d2b943264ca8e4ec38f3a6212ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7979e6bfc9b46c71740a7cb3c2ab9fe9ee994e92388ad197351624c5078cae5b5e5eac8b5ae0308ac13a457203;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h844cc847aa4b89af31e6434f853be9aa90028763eda87f86cc0515cc17b7b474d372db68f99d3167766dab78b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfbaabfee99b97b8c581e6c2df7d4936d894a83475eb4f42d680d4d99e36fda23182895558048f5ed2f4efd33c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138e21996e7f02c2397d2381b2e39d10b63231dd6bb502e36276b2f75c05fbcf19b412628ed4723f3df89637c3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2f32ff0f030edb2e25e15e69c2a5d34a62a44a6b38f21eeec49f3586f2c65ee6f6dd2383e2ad26905ff30eeda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0395bbe0e13d171196879d949c0fd65442dac9d001b1c1c5406191137680cda43fe950f8f343f545d68c1432a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc3ed9ccfe893647fd35f366e36a1aa00665b82baf30fe5cdf2e7c90fe7a98a3a28b4f99937d79ff5702cfcc95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f8358c637e5e26c94af08e7b15a32122a0e424b5d5cd05c371b33e9593f30dc9750cedc52e0ce70705ee36e9a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e118d34eb99d39ebf54d1466cbcf9b0c83b0eb48fd4fa7cf0e33120408e0a3f96161dc08777db58a31f22a011;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126d18bf5deb075e1cbc7cce5a755c659a4745119732daef64fd3ecef7c2472cc3e405261ccf8221a3b45db7c8b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd9bb1356f85dfedab33ebe461a2504e8961d3902971d1ae01f28bd6d14050732e6e545f93641ffd9955ccc214;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a19071a3c77116dc7ceaece4491a31928c69a83e44a0b2c742419a9d588e975fdf96d9b044fe2ead13319a975;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121b37c8b81bbfff2a33f348ea3f3ab7e0254e8639da89032793dee4dd431f4f3be2100082af8746d06a702724e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafff0571bfb85c2278259cdf973c0c8f090443a543cc639f4a6fc890d4b85ba24c204dd9f5c8eabf007c35926;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb225af70e053911e04dc889c15328962e86642800d48bb6a905a7cf87c03ebef59a24eeaa5b4ebdce668d6de7a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a560cb979f1831d6b10ad437eb6410931fd80033fa55c904496455bef72a5460eab3be8a478497494d9cd68ef;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52b88b956575087ce0736ad76f22e9cce777ef156377f064beb4a4b71045b1076406cfb92e4ba060fc8d1d58ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104c08ef281079748c4017cee3e8875411ff7c42e1e9c897ec91228d19756ae818e8d8d5eec5d6c9d00df1d66c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h749590730fbd62002f7f4c23ebd2aa46f0be31607e8103eff667e402e523670914386679b4bad76878b64ed356;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d4dd984faf091d5e1acd00b23a53504809f2eb2ac76e5e6e90e493bfb737fea6e9ac9c2081239e206468d7fbf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bce98aa8b9fc2b66f427e03c6f62dd753294d0f25baebd8d9b6a1d94a8862fd79f2e681d37120ced5a54f4543;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180e681f31e08eb3d1b3fba743fdb33bbbb6061e08ba898af2e3d13addc2f2be27eea09121e3a8cf9ceba5e50bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e0bed0f9618d7bfe86902ddc70b3b70a6fb3eb0c4504282130564231e611cf1c28a950b78ebcf6e6d04908213;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130cda63d51c8c1d0681f165dafd12b0717afe24e307ffa84589f07640ae538d7c96f6fc74609c52aee04523667;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6463ec215ac3e6a6a4662621b755662595f30d907e8d986182193e93f53ae73ef05d1e90b62d251782e3d3a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14064a06e88e6b544480e121cb2224c619c983071f632dd44568f55932bc57ab3d5d4c3f6c0caf897b0f3a0a79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1ee7d785869610aaa21e3eac6f56f1280d612580d18d49df6e51c8e1faddaa406bce50c8d816e8fc5a1067e0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b02c2cd1600f737bcb4852fe1bb6ed019a715041c62f159c94b382e2daf26e30e37cfe1930102fd36a9a357b0c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ba0193eadfaae48f690ebdf6b1250681d9c982ab55f6b35db9a7dc8ea3cf42c9a7081ad7b8eceab8b72c3cfaf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30b9de3e96d938b4d873ca25255cf6670368e8eeaee79d3accd657256398d013bcef187f4f9d52dbe50941f598;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13038d74154448dfa7b6b9bf95e492e6e7b41c7c2a872e62318615ad9cbfb6995a332d4ededb5e47d3e479fef46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h444d3124d68f0539f17a488b780fa7152cceda5abeafb5516584f68c733de55b6ce544ba19c3bcbfb1e4c1bd74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117bb7000dd6e1a85b0adae36f9260c9a2e57da7863ae0fa3857eef03266f2b2371a318641a53d3e7edfb3481a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ebc4bf33e83654a0c5f617e117b18b4a3fdbc7172c91e5eafb825a5df889c8155cfc817be1e6a56a73859f6cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a0eaf8ef78f7bc712ddb8622960e4265b5adadceaeb301ed98d2ff7456b7ca26518876dd34eeb627f60e8751d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18af41ca9efd0ec37d126e5d22ba58ee52ad6af659d9016112e1b0b1d4a565f9f0a7fb51a0bd9e66ba611766c87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a0ebfa22404c9b5fb706230d0f8eec6f4b343caa5e3fc30bf16cea1bd8de1daba8e4c15be8d21609018c8905e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1411a0c1fc3a637d28b032e7c26a58e53beb268a03608ad08c7b327bdb57c9ca9dfd48a675c4a094fc7eb8cc201;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d30c35b570fd31afed3b21e5145410ee8d7b857d071c888d71848b838f118d4ee54372b08da72d12cad918d495;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56b596432dc5960ca8ff8d0290e51bde20743ecb802f9b379791935efb991a7d694fc709d530f35446326500c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d8a3c55cde5a3068f4c54d83815d8c67ca7d937934b3616d077d9ae28a711a800c0dbac8018c40eb8e7363c1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e2fb38420a0609a811f5b553093a5a342b1f19b99becec75874a6b4533e41c98abd5aa1f632326a1e9a84711c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e8d94ac48230b117d21ac784896366a627d288eff60976230a201cf523d19a275232d964ebb7ba7e70eb776df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3c6c683f89270a07efba1592465291b0620c43fb2c35a5ed7ed0a8ada1febda4491737d72d347c16bc2132f3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124df90d8fc83c36d904535aa411af95aa23bb24539f21fe7b5156f2fd3079b91ad659cb0c747a8f11ffd4af692;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19411d8ca9e0d4a90f9ad82638764828f10ee080167eaf9532ac7157867610cad56c281b89f8be3849c1aa051a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb97e70876cc704f299e0e11fb41df480cd4afb7a73200d0a4069c7e778fc4637305a296b85e8e4d3a15d07896;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b9ae20926f3e4780eac7a9f7d6bdd0587b71e6b95ca5383de514243e006705be0b91095a087352f0e53f9c34b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165d8eaa62f715572ca9822e3fab7af5a3e1caaa994706acfa0b3202e39a73bf51a05adf3db781b3bdaba31a8c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14adcabcd5f962c096591611730c002a8ff91ae45666629173b3fe5f3a3746487160ae45f7c52e4712e67dcd8b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50ff0b82335911e04dffe5dd5c1fab44b1aa17e3eab4209407755ba35319031e884009bcf99d100f8d475842d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h700e11b04a03f3b5419cbd1a88be83024cce5a093c8384d0cac32e030fc3eb4ffd0ad4072b53fed6e65a6ad4bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c6792aa38bf27bde0769757a58d7dcfdd65bbe27be2703b1cb829af079ab90babf4c62b3c4dbed6325332f1ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108a77fe3cc5bd9e95d7e84a7f85d7261237faa15d2c12eae64c9680ff7ed157584fb8c9c47c7609426b73d5c10;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166d4ddd73f9ae8b4abde64352938f2e22dbd0c169b14ff4502f74b08a0f99031505d6de289ad129a902dd7dac9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4adf138f91866b16b275530abec189a990bac20f01e22833afaa2e5e2dce17dcb0099b1ebc3f99d36ced1f65b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134a207aaa576dd4b9a6a8048b4942ddd2bdb9897a7784ae15d4f2a78412f2d0b59f2bd242d41814063b312c48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17dc6c289d4c5c9bd18281387477a7d965d0405ded56a27e23b0e5b0104c8a71355bc03d4107d2106b3e44e13ba;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0d1934b6ceb8a40f9a5880fc4b739caa9466bd9014cc7d8824e560319e0ad72da028551b29f80a17f20c009c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb244c66c2b5411f0e82e34bd0471563264b2adb261e676a17672f190ec4edb46432e52d7f995b539f9454d0398;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2f6a736c3c9e3bca1f45c614feb824b904ca78244fa5f107ad19f424b5c6c61f88b3741a9e231acc7e6fe815a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haeb0e82d530c143633f5288766b983217b051a85f403b6335511972b8f72a44c90f8ed023b06aa559d342179fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b72a142db986f492ff221bb61097d59b7545d49d4e3da7c6a5af1b84c5b1278c30e985c27de74e1e7f42c34a78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44d23f5a01af71d0658ba4574dd330d203f0b9042440ac3f7d545044bf96fca67453aa9db4b01bfd7f96ebaa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1ae46e5626e91227208a67f02e171fb33c711033b0d7320ebb355f796b940fde687830b27007b833330b3d0cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h451acb4ba6bf9f7b09394b14060b20908b036867de3b6260fb5a4a3a1a9269cc9c5b532b24b8c561fa8478524a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf585f1f90fa3d80b8887363d911013b4323bb23aa2d457096b749716f94722f763f06528daf0dc59c3db22e1c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2a910af9e8c6860d551e15a790df9e0a6d1b1ecb0e8e95c68264277fd81674b5028d8f482334f1ae42330bd0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2fef3dd731d012ae6c0d22b22f696e426cdcc636dac8b7029ceffbf18fcc609cb57d6501bb7d21ce7a736918f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183804f99cba549a7b5b91e1195918e408d86294506f5403ea7c4eaf69eaf60d96de658c03395f7ec25b5d9614c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b40bd176b8358c5bb696fab1954cffc4d24328c72d9d146cac5d56a773875c5017884723f84f79a1a173705885;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee5e8f83f4a03c8b2fc56c3195269d8282a13f0244763c79dc40f4f222094706cc1ff73d2e6fc07075f520a548;
        #1
        $finish();
    end
endmodule
