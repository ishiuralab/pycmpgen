module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [28:0] src30;
    reg [27:0] src31;
    reg [26:0] src32;
    reg [25:0] src33;
    reg [24:0] src34;
    reg [23:0] src35;
    reg [22:0] src36;
    reg [21:0] src37;
    reg [20:0] src38;
    reg [19:0] src39;
    reg [18:0] src40;
    reg [17:0] src41;
    reg [16:0] src42;
    reg [15:0] src43;
    reg [14:0] src44;
    reg [13:0] src45;
    reg [12:0] src46;
    reg [11:0] src47;
    reg [10:0] src48;
    reg [9:0] src49;
    reg [8:0] src50;
    reg [7:0] src51;
    reg [6:0] src52;
    reg [5:0] src53;
    reg [4:0] src54;
    reg [3:0] src55;
    reg [2:0] src56;
    reg [1:0] src57;
    reg [0:0] src58;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [59:0] srcsum;
    wire [59:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3])<<55) + ((src56[0] + src56[1] + src56[2])<<56) + ((src57[0] + src57[1])<<57) + ((src58[0])<<58);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f15d2d6e44d21e953038bdb4623d8e2ffcb2b8031b876c44fbfac7559904894a40035182d8a68036c63acf925661cd8c0b4dcf388771efc7d4250976f284eba33a10183dc8c56780ce00f16e788f73fdb903f23875b22018128d33062d5ff53be9bd0aaa0ffc50d91a6d0f19bc6996f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha285e1392b1e3de538eed49e6fc81e983a03997ec9f33cfe034e7dcf1e72ccdf1fea97d42dd475321215f9fbdd06281b274cad9a5b8496ff24320b00f422be9d0590c57708c4a1af711f09072f54b69e670c4c91f0ad50f78eb0b1b04a30a14aa76b2a11870a2f442ff5931f693ad60a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99d3476969278eafa15164d9cd7424e08287efaebfa912e01659633d7f04e02dfa9a7ede3cd8f2cb1cb474011361aca8aee2f9af127a2e3eb32355b10079597d66cb6516f2e4c1be92a0430151211a602e3f3b898747500ec85ed1e2dbed24d9c36b9f266c0288c6f483b8f6b5b4282c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cf7915bd59f85eea1b888a8dbc6d7ccf7834ddd6bf87b0c186516b6a29e3a396d881fbc998f163c7b7c911ceda49bf6a853f673a8cb76c9803962e121f641bd4636d1cf51cd9a6c2fc70dd108029f3a6b7a79e484e9a2a92bb2b60bb148c8d3271319a3eb02e0f9e65f20798c4bc6e15;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf593e98575ff87dc4bd8c926b91a211ba8cfa6e022a513a400745011e5f1a2053e18b9853ba8b641f38a31a23a950f6e2ffb1628a81994237fe2a6613e5edc22af0500a57e492795a26bbbea5ee8d9df871a82634318e9bcbd839bb95d26cd8abaab385434ad85ec9a666996b081337c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9df7acd5ffb227c2eb96d2af4b3fa2ce893339f553d7b84a5e851045ad6cee59b29342e0d4ecfe138043cbe89f00d946b711f2a56679bb6973f9e6098dda44bb999b5a7656a07ddfcce2b132d14d520d2e61244aaa473abdc45d1074a382d1161c4a3d6ff65fd7b0e75e28fd428be19e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eed1609b617a47839ad85ddad8d83b578825af8402f94038ca298e1816cd1f9bd36a36c7a24bed3a52a505f3e3297a56f32f9d1ea996f936194affcd6eacbd541c1d61fae4e6c2ea2311769236ecd79548a5218b846b4fbc74dd74dc9017ee4e53cb2111aa8361e6a7ab6433ca25110e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2e6d3582005707257437addbe9d631913255383eea82d79098ed9554c732691d35abe6b591299d2fd85ac05af919655978868a2b6bca63f223e99e41c58b35ee3728718879474880f715b29b9205022a88edafb9a70279778c2163b4d7b5a753a3bd66db2348f65ee7c08ec8ca6eaec4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90882724bae3cd26616155fc799677977d13bd9e14c3aa79c88944fff3b3cf92b690062e0dc38680c9db9ef962ce49aacceb450a284c54d6e79cce657e03c030b777ac730fc750e7c74c4f1e72f3413822264b598e9f151e32ccb6e7bb04f0583f1f7369022fe58c2c9cc8df046838d35;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf416cd773ca1a98298fc179740959845399b72cc963c7b79d9f1e82bb76bbc3820681f662b1d20c14fb604162a144de101536e14ca8e6025d9cdbe7e35bb669bbd7ffa2ff5dfd98750643c52d00e60671d92a3d7789cd38ff9302c0ddf689e1599960cd8879a5053406b1376b6c217f29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dac09d6b96e3d946a0062175309a918556f6856d5530c5fd368e92e47708519cf64e4d18d9b73a73b8009731aba792bbca6d4ed3c4dd87ffbfb6ef92ddc84a3c3cc20dde79be7d0fa5e2ee3a06d7b67f07ebcc0fb2ec77f4aeb5e3a6745a45b94c7009730d755cd7823627c77e4cfd7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb9abcd0a73db170ef7ee60c4ee3f2dcf20975854f2b6a8b025668455bfacd4231bdaa321da623708fb9905c3b251bd2be1dc127dcdae5f1b884d2233565522ee8a60ec3e7965e9eb585f1349783b852cc7ba95974bd3fab0dd6b5cc2d551f5fa36a4f96e3ffd88500a45558d9733773f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35fda1e20308dfa9676d2c3860fcfa891791c0ff0d07f58e8230d7c56485f0ef6840424af61eba09c96e4c8d8092e8dfff0579700d9c5cdf1156b04ef8db762505ac2f93e53fe27c3c3c4b20e880dc9adbfa44dd52e55f2f1f1f61e4ec0ed6f0acec4b4664451f76ba5c799076cca200b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcb50fc63bf2a24e46ceffe313cf2d3bab324c9232e7746f34f7f9afa50d270864fcdc828eed95eb67206eb55b0ed6e919495253169d767352a2b4fde1fa10db7be6ec0c9e16f7aaefbb0f323fbd7b15f42a197c4041bfed43cdfdbba6f8e54fd59aea46674f5ba8fb792078f37ca545f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he034657ccf6a2e6302ef3f949f407750b4e43a25ea85d4e959ef3cb7267f2b92b1bc9abef656a8253941d359341a54ea9b22e60d8af61a76605e38d1bb26cce474d29fe0bbc273e478117fab4b8f2d0554781b81be892921f5524f9cef6cd590c6d1797a0da1ebfa38b838786e975d57d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f0257426379f3dbb089533fe05e8568ad8f8690ed122874c5694cb3935d4c1c42f08867e04270a90edc506c116acdd2b2ee7cd55aaf123240a7006cd90e6676b7ffcd3956f655f845afbdae65007a5378532906cabf1d29855d3a1535a65f0bc5526b5aa768619c5aeffb6e7d0d20210;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27da944a6e4011bee276397825bcab1a8dc1771d7ef6c7ba92c9657d4278084c270b2ae03f427e4d00309dcf4cb2a2e4a1c155639d54671b53c429bcab3d2b792a48f90f2cee136ad307f1262bfec103026591f9b94d88623fc0d874c3835dfb85adfbb791e1fa3fde3cacb74ebf660d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60ad9a83760d84e573c843cb1af221aef8a660af747129329cf89ddc519bf2d29048a646c63caa1ad6a4015d11d8f731c9a38a9610ad408fc639bad0ce5007fd04a62492f71e0c89a78de395d432524518c4930f6fb1a9cfedf437cd2ff01d6c28796e13f784fef3113f0902d96734c9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17998ee4041ff9eb1c123174a92c6ee710a11a7e4f1fd091b36a7af56abba55accb3d95438ce539fc5b686a73741d5e74fe39e84e9079b02f94209b91045f04f34cd0940fb0e0e08d9dcd28dd368a9a5f2de0ede1c6da22ab173e238f525377d3c6de3fc16e711f19e53916b9be42d53f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b6fa412b8be0db8fbb240cfc86f8b98ec56a6bc2a3ed6e2819ce6abd175021ef98d9ffa85671d0e151db204869786d1d126c9922f596e80a4fc61e03a3bd8ee816231b561cf1bbf6942d4bd32b8e9daa0d9d93ead1a2a5c36b02941783d5dbc1c0cfb5b0fdb93a776d75f58a1f9b7bd5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83a53d7c1f2b1b382f3e0ca94044312b67d152fd9af03a4b971a37e520fd52809ec40279c0df2521142da7dff77395af14dfb0e6611dfb68f3615dd8dfe337aa117290d94b4415a1078413a8102d01030b0cab4ff5510f695603cab1ae8b6851e5f438b728f0ace572f3aad6977713e0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h503ab0172671aed1dcd267f9813aba6cb435c4a49eb5328c1574433607307a71a9cecb177301c81bd3552a78f1cc4732f8c8bfbda924dcfe4c68abbed83da6ebd9baba471d3d9abec20babd54f4701dcf9b99539604fc9271aee787c286ed50acbc55c2cf776394e41217cf88de4ea7c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12cf9179c21927aee1568d14561ca88bc5ac3e89a59bb277a786b3b73edf82d75d2805d90497e0ba73e4cf22df8b15b04abe4c36ac0d5fbddcc2e4230621040ec1928a94f0d3af0d66f62d4978fab75772901aed4bbf49e2de0cb8bf7cbdda869b61d87f235b80b7d6cd28465b48c412f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7361afd179f33ab1e369c62ce10b198efdb8c909f6551d495d068515d0bacd5e6a32320ec001780e486a588fbef558c54671679864364a9169f842f49addf39dbbf25766b2b68e5b834b630a73bfdf7ba7237f6b8f2d71bf9245828c21d587d9ed92504463aeb574c4811c9562d9567a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7daef483eea94ea43bf70373adefeb43e7ae43991496afddc1e2a1d1846e7a216a4300a708e77f5566cc8bc18803b62086618f00ce56a5124f304b3f7ec5fe3323e38e463da3fa3958fe254735176ae921eb05fdf10760f218f16d4da98f50eb0e5f2e960d474ba0d8427f78ca863978;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h166e20dacc1b5b2df7eaa81fafa3e74e855150cfa9836cd30012708788999595168f5e12753f4155e91d6e1303734fa79f81dcb88485ffb18a865a6eb766172f0d4f959b472567015d1acceaa3c03f456b7b2d8af7fb54095fe5364f2dfd5a0f59aad2641569c282666ce9194d08343e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h836a53954a49e4c42bbefcc884ee2db462ec913215f3b9ec3ac4f1f0853ba07a028c71d12c4f4c8763300e81a3083314454750526ad25827ce26feb44cdf45f199018758fcfe8a21180c7419154fab95e92bf059a20953e18e905aba7e101f11d535b529487fc89eafebac19f40180d37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56adaefbfbbaabf41fd22374bb5ab3cea6989d0cb48407bf39f482bf3cc27519f9d18497f50f9fd12531ce8fe20f1c035f9bbfb5c64baf6d480b4df3d7293e21e935775fbc2d30c65d256cd990b1153b9d7dc1c310997bd1a6a605d677efb57e5ca4f412c57828cfb07662d61db6d4b96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c6658a38fcb571edc27bebe905200debf43f688fae8a3e723ff08b7e0e3f60e85b8a3f60ce4bc63861e5241c3ff3b05308de73ffcfceadbed54254cdff0a2f264b7a15e34421f2794bcf129babb99586afd54608b1e716a53f63a7b713bc6b0fa9f81585a78145bae8a26e10f7c6a4ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3ab1171b37d8106e9daf7ad91d4fb2b17aae251dceb5bd32088b2ddcaddf87b5f99c0c63454785ad0b2c39a44f50ee668ad8bf8e4c08c5a2055a82a469cee3684c3a7624ef86345d6f37775ba177d7335d77fe9bccf1a32a502b5dac25520e2f8f56b0f481e38dd95b0e09c562660d2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cd584d51b29605173890dbe201ee907610bf30c40332a4016c94c46dc9a60b2d569a387958a9c9c2a0bdf0f94c094c16094a412b1e2238ab3ef3ff668d953cc015491c5cf64f5f267086dd5e82521bff78f5e73dcda6ff99b757b29cbd6537ff7a356de403a82afc7a530e675103a547;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55ea6b8ac28ead4b6d1856a1aff86cfa75fa29d53bd549c0fdf837b9aac47ad8de1a2f0f8a9ee8bbb465f1037f3cf2b82d7d26b87ad992811412e64074721086b2cda813c774233f22ec930d9331dc295741c9b9f7293975ff86389c05a9b49f9511182f7ddd6f4e4cf9a42de064cbf6b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb789ed670873a8e1823de12c90522b73b5629e603841d369e27a7dab1cba456e57076d7edf7ef0d0840614cb97a81d877a2503b72249e2496b0b8e6123c5756ab0818083d1dc5b1b02fb78a9bd0bd3cae9dc1387cfa97162ebd66a25419e97957f812782b139caa71d366d3bedad9b386;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbedc13a6a1dba25d4ce0b6d110d32a2aad136edbc585646d6a7a9d585b62cdba91f9af3fdbead3e053ba56761aa7b1ae2ed28a78c989893922b605a187586c206a4886930087a2e860b8064ab26ac7b74e6a158584e4eabb5ab94fb76ed77c5223e02bb298537dfd4e32216092e0c27e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hace520d9758dde4bb061af500499a390790b34ce69c4a94ac6e359e9f0e684e4bdb8e9fafaaeed2b394070e9b883ea48e811e81af4028ecd08913eaa349ee1a1e97500c5420c87c19de5aa12e4bde4d009bd3bd0f6da1acecb9721f3d6b832a70676a794a56c0bea05805cd767c1b543c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b707b6acf1af08e2871775d01fac9825e8cd367f162237a30499b491a25a3ae312857195c3015c2721185e54e58743e06d0bcb8a05eb7f080a1201c8fad00fe82ed3398d65df5cd359551305209226eafafed79e0aa6f3715a563c7092e6004730ccadaf7c334fb2c7ed5d5d772e384e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcba7e835ca8c689257c871bf595ca96293dc1c90776415a5250ec655983df43ef13ffd6f246ff999e193c17b9bdf69fa5a0e1e3aa8f0b4b95e4b0d09aeacbfde6da51f234b14e6c33cfad04e66d3816972aab8f3f04498826a0d4581fe0a04f2e92a50d7018d6acebbe0f91ee7246c0c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbb1021da8c05d8beb1cadacfe626f07eae15dc780633e899a9a3659a88c34eba08b095819d132dae273a942cb48b2e7fc6b435e2a212694fcaff5c0135341feac553c5fe1e509091dd04a65f5aa85408fd9488f573ab7c861051117e5aa4ecb847bd05d8ad29bb933478ab5d4f3b89cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4163f8ba32119b74c8d640c736838fc8287cc9b5f1b3345ad4f7b3e7af841ec639f68f88832ee3ab8b3fbf2fc83c62e2a1363f19351365722089873894f5a35b8423b6d08038193066efcde30508d283492334595acb6d770832135fe8633c2a6ea3682cc8b4639da6d006ed40ac315d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89c5f24ec616c5dc496d49ad7d50fa5fa8ad507bf8cd8f66badf2376623df3ff528e8f1ce226a95384fc04733a1cf39c704a14005d39723094a286186fc7bb34f6e9e59b6276f5772e03f5a8e2d601c428f6c0a59aad6b0d49854b3ea4059ac4b5497a6b31fbcfd2c00a632624e018262;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8efcc12bd88bf7ff26fbdc7b94947e28dcc57ed02e3e02ca93cd5f93b0aa8438dece4fcbb0201579a7330f4479914e61e4f073d6c8ee88301d945538c3feaec1c81d824cf080efc8f2b7fc7c9efa66b2d06236d03b2e35c707533b94ca80b3b7958722080d8200fc38fb7c9acfdcf5ff6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e08b4c8e4738191ed7e78d6a14c67b064bcf759ffa770bc1c6aab67b2674664df27f46a95bd537dfc3ec17c8a0c9a0d84158839f7fd541503b494586a8177c3d66c2d646108c381243c709877825de4ce2b9547b2318c6c094d8cfaa72d98ac4b6de0c5b4e43f67ee7ebe4e24a63814e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he091a09437d9e66dc02147c6ee62b5eb7c1c4bcbe95092983594006a32746fc335954405944e45d0e1f7bc85689bc743a2108e6b63cf7194fb67d263628b0d2ae27b4e1c9bfd1d9e45783b771227f7931f4a629a35dc9a1cfb4e35de8bc9711bd6d39e57082abaf84732d2522c0843c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe2e51ab4837b2ae3e8ac7ab0c8ed0c9e63e7152495f24cbb1066ae6a2f21e7659220a9ccb72b82cfaf8e3bf185729472c2c743c9acc81d30c525b8de1bb90e95fa141ab8f2aabb72dbfccc353839de89d23804329d44f30527733541fae11903d3d9a1fd740da2ab20e5cc3b27601580;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1e5e76ddf8b94327ab1642818d2d7b4f8256aa7d09bcaf365c54ce74416f22d3b8589f443f5b0e28ba0fc03d8d8ca475514019b837489d2efe92c1f4a9d9d90f57e446d6c6b3d3f388a9f9e074e5a499906a99f527b8333fd68f811dfb960db0539276058a4bd6be607645c8fa7a678e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51b98f0eb2a620d5e90cf608644a93a99c7f3dd730b509ed79df2b8ae03c533c10a2c4c09e190c19cde2c94f703067bf953123ed575f6d4283f89fee45a1852139318c36b705540cc7fa7285bbb92c143070bfbed38cc7c59cc81ea834909ec4178a322ee48d441be7beb828c59be2587;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafcaf2cdd02b02b7e2c8889b43d743377f12109f7214a2ebf91a01e310a234f135dead542966797d8857d164a277e7d3379d1272a26119e5316a8b1919ad8bc1fc9e7695eb97ad89f1327a6dba0a5ff407f96e028abe03cab3fda6eb3e6321b2fcbdcc88823dfba959d6f26b722f4656b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3384ccc2ab97d4a22bdaa5924554755f48a5da65c473dfac1efeae7fb5850de6951d58e070ed2b77ba4bded742d476ad8797bd07a9997f20f953e7f804e2ce66acbfdffa5ecb069d1f6ca2a410cf85c712457f6d5a77d506bf4f70a9ba863cafbb042ae714c6d4175e9b5131138de30ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he75cd064c558b2b7cfb3a6a38824e446bd8028e3292c31e1e43f75e25a1c025c89a416b897c12dbdeb46c29687384b4e3c0b2c84b54eff96be1cbf773229ed0c80b945e2dfccd45a190d7e1bde12114435c9d9b0c868939c1bb71e95e92b491dc5854397fd34e699f6999a75196f23168;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4bbcb05032e431a7af9e7601d64bda1c53bf68a233a34735b14722124097e47059388540d8022e88f4fecb8dd094e390a35ab6de83485ded5ecabb803fbf400382ca91133350356cf254b8e14a750d1d951fac247afa934e2d6c1402ad494a0e44436331fafb3b546273cb785a1f3f2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c8c7512a1927cd7402c7121cc7963628a8c2412ecffc3c395738b7f6e905df63d30eea8685f376925df47a5089561cc29ae5399fde46248b5332bf5e50cb0795f5ee35ed73c547dfad1e9a16decce4e7147ea4d3f7ed7798d94de9c8f366762f6efb334c83d2c1a21b45d45a59f76881;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bf6f250e25481c2c6956d48ba6ac7625f470af4a4434e32b64966880aca7dc562c55a5a11864e866f486c8d4c91226e1d286ad1dc7c8c31b1d0e8f36ad78a07d9aaabca7c1aa86ad6f38d42be466aa169114516861e77414a837dca45276ca59da32f2925064ebc743b3df722242f219;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfae5f47437cd94b6ad1b0aa598f33ac994e4628d3b9ecf32817696336215f4300be087eefe566f334055c92fbb7c93bebaafc11338e6cc2c75001af887eb05f9cafde23b809df12d8dc759ab1d869381000045cef06496042940e9cb6c85252b6bb0b04b1c3006b02c93e56276be60be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he162c44d78c0cf99c5faeb53d157ae642db228a3d781c5dbc3d2a8d0e873ec9c674a3b27b188da36b63effbb4cc9ebb91ee07748bd83a5b38015b5b7ac9056ccc5ef7fbdf6ee27c3ab7c826784e6425f511da01c15640bb65dc74e840cdecf2cc4a27a26e1b154f69a2dbea219053e5c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e5a59e965ac63490c008cc96c61f037e39bd954827fc76bea7146f84360efeaf188cb97213a2ecc0f70f9af099232e16f7a4e5ddbc75d5a5d86cd3236498eb32f36e6e512ea7d93b7a5081a72deae8c02bddb6e724f1a5b25b4f1248463eda599f1db1edc3ffd8aad51acac23bc2f91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dde7fe529f0eadb47a4ee6c2875b1b0a54bcc2c5f5843e9482ef66833aad59bf1287437ba95a6475a1c6c7a7495c04e2db87a93983c00730194e946d3324afa2baae692ba1eb25f339693163c23a77137b710cdedbf872c0753995f0097e18acd9a2d46bf67cf11c8a02ed8139659828;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcfe50dc1cde5ea0335ad3f63dcdae2c390297b580e4db81f73797e753a90a313376b80853c5661cdbb336187ec648f0a508ccf7db97710bb360d1a63b2bed5cd36b4c2d8176df434e28e925f7a7edb2f953332981e5f45a1a01da17a54f619000586016b4309d653e747287561975ce9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e803dade1c6385de5cbc71ef35d8be53ef38c2d116bc093e31e60f7d670cef78d0aee7c7db4c1d139f33b90e1ea66a87a158c72f3631c040c65e06c4c4aa68045c70b371fcb79b93a88214600fbbd461b0b7e7c4780e56e798fdbfc65b9eb4a9be3a3232998f307cd88b9ecf6760b32c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6d9a1282b224422f4246e890754766a1823d80c0543e166bdbce3a89bc706c6b9043cf634484234655006e961a30a440ccb0748be49901e63bff5846f7b1f8a58a9c3a255c6eb20b4b908cf0867ac67b40a79118e2ea4d3a1c09bc32c622ae0b64d4ca5bd73718364164a9816eb9ec31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd614e46a557519a4513f6921fd10ead547222304800c107d12ac32bc0120a99bde81e98f9f2db99d2a60aff8fc1b2a6d0a53838b1692123396326e577499d7e27f556c780cf4206893f9f6e813a79a2352540ec55c34732932e9b6cf5b4b421661caa31ba58e11f31d6ca3f92be63c18d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4707aac943cd89642c4eae05fe3fae20fca73c71b244b0181c370937663667679752c728e89da55972cfce92fc749ab58243fc1bce2a86cabf574a45de65556707b93c1d885a19e57657a21600a17747ac394193205845009b799c806d9566d4e5717ab637c35b56636b973d790abc5bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd64e1b70f7bead5ac587209e8a7a2ab01b8f2b306478eabc3d7b3958123a136ed46ca162199ae16b5b2d846e566aa9d7f715fa23f8fd70b98c961874d4e8effa53c94d8114685870144b2cae003e17e10c21c1fdbe642e3cebaa88f6ecd013884960d661be13037fd4c7f0c74483dc6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfef444854ad4ac6793765803dd2e50c838ae2d9c2f9fc435c6535cccfa8af44cc20bbef59fa69061dfcc79fabec22bb4a751b5e8317b0a41429af3cf60c9515135e03e5a1c65a3114657ede648a23f552120f5ecc155e4d958623b0e46870f060e0dd4f1b80c0a9fad09796f401487e6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33a0470eb4bf019c254c28c4d23a19293cc2b25f71ced07665adf5f3ec56787ec334268b36c3df24eb6386e6e6f27c6b0c0735c3a9d5fb91c1f72bf826402423f4aff041ddc01d95cc2a2206f302151f110ba2a472dcf00da79c02e52031a551695f9caa831c26b25966d459c649568c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5605918664b74b4a5c2a99d94f6328a8cbf04ebcea42eb51daf97dd4e949dafc758bd148345520b5889aa2d71be673b30dc65b2dc8bc9bc64a5e16c92bb0945a4fb9968490551931a645f6e4b2b2760290be6246b33a6b93b8630cfee30fc303c568ed05b24ae73488858b2bc0b032e23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8a97d8da955b958e80a9f36047a618753c8caa7c574307c6e8108cc4980437d55ee66ba5bd391291afa878b9e194f1a1c4ca7aa4334b1fa18bc22f6ffd701ecb7f50ff3361353ddc05b73ffe72966eff95cd29bea69f7110f7c3b1e89b32924854f13868681c5dd98c5ac27656664a45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9487bce2e0b15ac71bdaeb0dd43a8bbb9802045361f76520a1f1eef44500e57629d48bb1cb99378b3ff7725b44a523a37ab591986a4eabeb3ff017487b4790ef17959af4bc5fee7b0a0608653ab8166770f990ea6413bf0fa357a795e6aa455f0fa0d4ecc9c23d0b19ceb6adb35912da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e6e1998daf0c547a253675cc2bb4c7c466c942ff337bd5c70806e8fdd1ff4fafa14e02fa667e52c7c61fa3b3e3559707a5c5587af43f1bc42b0c9383f635c9e6dcf36e9d3928eeb798ab0fb1689a4b381edac059d1aa42fe3dba1377eebcac2012aed1ac0f9e1b6a7d8880135dde3e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44cdac59168e51333e26cc01b993664421ee520fa83e31f03e87613e6df37cffbb743335b2ee7b75a0fa712629ffe8f6588dc397268529c535cc226b8ca8d593918932dbdd6bff7d4421cef2038b689c50ffab1a6450f2968923fa7c37c7229d80706b2ef40cc357f7673897394d623c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ddfc2701349c585f24b3e6b71790a7e1433c3cc957e7c22fc946af86a5f72228cf789aa8947d930a86d1b186a25f793028446fae2cf5c8a20fb3c0629f75ef74b6c9ba935c46e125c5b186b1094261daabde4f6864e3566628a3bb39b81ae0ec98741206b3dd956a3a7d085a2dc1b02d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f62c7937a5fde688b66fc9cbb608046b2786b43a863997429ed20e4b8c10bd0bbbceb11ad05d1d1d115bb88187de7fc5ef065890798aa15fa5ea9b9add2df45bc870ce585dfe6561171067eaab96aa0ad351ec043ec929a243460de1f02bc489c4ceefd7273ed07b1cb145b5a379c6a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94f913cc691a600e0f407b984bd6a3c06e606e6b3869848b97ec68801b14c97d6093d0cebe8b655f6a6757fc53b7de9d989992290cc12495be0021356046d5df90bc68e2fd8eca892e2b52649c87c28e0b1041c8743bbbfc36c079829b7bd65003b65bb0cef5af709278eeb7bd997f547;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26934e607b4d2bd47a23e85555e5b01975cbb794c11bc4bcf5c2ccaf55d773da14668b5c07ce68c80ae3863fc35b1eb5c25a2a4acb67d7c0f1fde41744ce44b45fe6a506680e083b36ef9f4f49694b187a86303fa0aeeca4edd1448e4c6fc99e83bb4ff1dd6b80e5472b88af7cffdbf1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb22b04a3c91df44b1ce0e49c5a823c545984a7311a8f0096421af762b6ab1c46c8441fcfce94c147afafb53c5d5d628f21b7fbcb291fc4531b5cd11755471b78c5e2cbcc91fe2d33b69e8b9f76defa3af6ce1739e05034baea5201ab8605c214d134a12f967756eed52bda39b619789bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3795e26d4146824b01bad8bc08f84875d1d56c76bbfe26029eecd4efc72ccc6f1aa3576903490f174a08c36e7efa23bca1cb07317aad879b1e6b24b344d57682535e0b3d87a259001bf9d4dfa47b5c534474266de9482df37579758c7472d98e8d2d5bb70d0b73eafa6f2d29bb7d97163;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e4e28167927e5f3a943f1087095db9d1b7b517ec4328181d9d612ca5434a59c3675dcf53f7b0697f07b43fd080a2f172f53b1708df4ed8c1d7387d742a3e6fba96a779628b8354ab61a17f19ae23ac05f9115a9c997f69f68dee75fe1de728dac32f67f2ad0c694776b229a263132f3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3a6e9f556f1a91a63cb1766f025afc4f71f968253581c2801bd851f99896a74342d64500a2f19637d7acdd06e13a43ff29cdb466acb5ad39fa8febb2a1c4ec3d7fa4667b29d68ebee1b4d7b6f9ddc6f2c044da8d475613dc94f59add08ffe559ff6e29c78f0f0d182da9dee8e735264d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h248be63f86c7409f3b3fd293abd957024a89b85094f5cc4d873c09b4dcb17c3e66a1efe20366a107f20ffb374d0e42c591f2ceb5b62e9a6373d7839244078b1818b404f64e18a28089b28efb907a7c5466466018003cdd9de709906c77ec700d219753df91c2e2fe981272d817e63477a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b73ad209e1ccd17237d302ce91c3aadac8c1422f8b85180453637849e69f8d18533a710cb094a4f1019fd3c059f14b79747ed66b88b7f1be0a016a0696450c4105ff0c3cc843c8abc5b45c72e56a39ef88bc2d94c2fe66d5dcc54940764503d3b427906b2c8949306180d7a0eea09896;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h596f73cb5ee37b3bc275d74da95cc9986b5ea29c4fd05e69fcdef9361c995eb505132336a9be37f0c8c94dc138815a13c8c74b27e25ec2d747fc9a7fa72f46f1f2eab51b5e208be75bc4e917c09a5ed8fdb04145a2c65c521c11ab7c079bb016f506416dc0acecf77b9ef7ee61904fc5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60fa53e1b345426834af4282e761aa717565a54d13a0b8e2439ddf3afb3be9185569f7d5255f5a40756e95a773edfca94975e5c2bfdf8f0df6e6847a8e1396e22209844740eda176c53875ea67f6ea54925425cc22f452c27fc2fc4d471bb60ee1526f153dc15ab12eae403aade048a74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h512c999f42ee23334ce0cb37636ba58596eb5f2df3dc5cc95b2488d093bb19d214ff02de78fa91bd855f00c4cb152621462ec3a9e25b2058a72b8c2665ce07f73dd6c1ea790b7cd34370a75118b1930b87eb179ac46ae0f9759d891fa097bfca5c702e1a0be61cdd3441ab8747b874772;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7949cadaf99c060131f9aaf7777e3ba66858d65d1a6d25b1d28e88d4dbb00f09aaa10bee7d2b6ec6f208b2b76618f4f455a6f408c4868b0a4d316ba07253fa383ac16f6e80672d0ec18ceeb0e47b797d5e19a085e745c6513604aa306b0d9733772a7670dbd6993da6dc8adf9190fc8f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73908725b83a8a43a8f8619e5d662f41843503f6a91e1deb4679ce3cff160a2b4d3c72511369ca9963253f34296b6dc65a6265915005cdaced3252a7c58828fa8678b59d237870fc7e74b881c7e4b25d0aa45bdc8b0cd63e019c9e2369d7369c3c23b6a22edf60984da27e2abe44a56a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ebb79130a4ccd28afa5f6447ddc0bb504c9df9cb2935b539756765ea73f9c9f91bc3432a724b82c415879752bc4af2c8c7269724ae7c705cde3880fb9922eda5c0aacedc524bade3715718dcaba08281b24db3b9e349883c074fb3b883b901a31cd99a2994c7ecff55fbdd73d7d687e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6efa45c45c6c8cdb73d1c586033d319a40984d2db2344cc92b58b75dbd378efc22452fdf35ac9b63ae60333b9ebed0d033b2c0294a50c34ff52eef75b319a016ae947323c3a914146c7f049dbcd46a15ffce651520ab9b0f00598312bfd77cb9e9dd39e3a5581f3ef5efca6477caabe2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1747331b259142e3e3eb2e97500ad0b8347b426626b079ea81dad3b50b9593a50b4283d5939cb4635f22d23df25f965a1ed146515b6dd40439564539045e42a7bfe7d828fa85a668b2c33eabea8465dc8532c3cc15c96c5f954570010bfd3a76447c0670444f6104605373e914b0c8926;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50b21cf0c744cdbed749def7692159c920de1697f38f98a98a0f38079ebefb57c491a6956638a9911587acd5218c57c22caa822689fa2f815484886d9af05015e130470c267dbeb6f4585e3913c655e6a6673512ba72932a6c717d751f198acf672f2e5f51cd7e7b725a5bbf942668f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h593c10b3fbde633f26fb9f345a56cbf58401c4064cd2616e7172aebfe6d53aa98b503566a11d2015876b167b3f01c861f832c8d8b8a263f9c7e071ac9d55e5c0e58110a576c0176f05ed876e97315367f765c870136ad41553dc9619c04b5928c6df5c27e95531a6d1225aeec17cf8f22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff0c83b0f6a15fd88624ae394627b9704b837d88bb7e91ef7b769f89c84eb15c3c7551b8900d1715dd0909bca6c69c41752f79255e228da75b25514c202f18a7e90c735beeb6acc1b6ba9c3b43001f7847ec0624fc5ef5c5c86cb45ccd06b802f2f7a5718597e149461d222bc7f1d1143;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac122e9820dd13cc58dc9caacc515b4d62d42b4e5e047024e7f3bc7f32f2318bcac9efc94925b2d8c830050f834752818665aae9a18bfa83d0404d0867f9195c80377b26b31d9afa641243711a9a369aa73a575c8be9687584ebd57ee58c98586696d2e8228e32b2916a37f7c96a0c31d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4125356ea0d812eb9e934602148ab7de3761d519dd4e886d8e31b71670d5bb30ffab6c1a5d378fb9c788d65b06ac276da291517d43ec3a38667e0b0a386b6c491934176c7bb2fdeb1f986544f47bc69d770b5ed8612e6d9ae0ad8f7e0dbe1b92307186eac6faac1e42796723b55ae43d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96fc1ff2777039cb74610da5c80e39e8ab07cb5ed41461725326309d9d9d8b9b4aafb2f32bda63e6932e7e4495f2e0a9493e4b63667315b61bc9cb2b9f4a9853025c22444b83a4e3db6264b17f0efa21d7b74894eda5a38592f5fce8a6d40cd324780d539befe26cb38f81f35ee3cde70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2de1acb7aa4458e4361e8069f78bc0929d8509c9d9ff96d5ed19897d2cb22c663cf1de60bb54950bee59bb2da1445645e6cb920ad163056002aad94326028d961db2822b4bc065b810354c19fc0cdeefb8de29eac5bb00d5509f31d3aafbc304af8d1f2ead6065ff4dcd955b1bff4864e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd2c9c4757c1ee8bf146d70d639484ca63f9486582d7e25e73a051b469a6a9ec893f7699d2591240f3909f06af6660b855aa40e04aa2bd5039691735cbfe2cf50908f50f2b93d5e02c803f4607fc849148c17942bc97bcf83198364aa6e966eccaf5b1ff5eede86ee0ae56d6a524c0782;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h807d6b37cd33cdf9732477aa7ecd1de923afaf7b2b8ed170f49b32295c0dab6c09c74606257e2df843f764635a82693fa11609ea4ae7a22b4b7b61f1664485ad57930f7baed73ca5fa7615e57ef7e65187363c136b4def0994e3676eaab2949d5b9c07adbc71e674688ec11cbe55b9a2f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8975d2782742e6fdf27505620cabff828398c544638810e493487b2d8a6119161be251e3bb09d28636d6fcb1cded1b4ea26f4c3176fa46bf0c0af1bd4dcbb1a909473e0c1196eb80677632baf78a9b79315a962b8b2a71e969edb6487743d88eb10e3b0a8230b23386ea8c40328c33e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6a360d1ff79838ae1ad4dd0f8ee7f1c093a9f111d03285779941b5d04dfbcd7a8370ba4b568af7791da92d0191cbee108c136f859f98bdbac61e0aac6d927c1e883e4bd03c29ece1276999f73a692c3591551d68239a127bf7f8af9a0ffa071a38171303966b138bf05484fb14f6511;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ba24d3598e2eb369325e78aecb9bba614675b3d7fc777bca88e7026829ffc4bb3b9f07f4b80c83dbaaac2dfc918fc03ac5fd79598796f3b8496cb971fc85d2402023f3a5ee5b0b1aa33cf5c7f12cdc6ed6a8ead7a675d49ea882117f14ed09458a69440cafc68590ac018be1ddfe5483;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5723cf42473c8a88d4d00a1cd7f2fdf018d257de2c620233ea4c916056f74796da4461dd8a7865636b257afa3b65c991a0cb5df79c9fe49f5d329a20304f9e7b5b02f5309b00b96489b1f1bc358db4619ad1880a5f9f9948c5686e1611c28c5670a9dc48ee12fa1d243e611fa2786fba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77cf54e378415b45440096b8548bb15a1c93fe02d07e5f84afc1083bff4043cba9d56d90a3793c0bcdae8ec0e3d0df71b58586472c3810d9a9906717fc12e7462ce5685acfe22619c9a89befc6d4ee57dd8cc834b0c6d1125421a529f9224b72e6334ea5792f2531f4c1e2f631923355f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb24b2f1e50d9330f34b7125ee2e253dea6f8647d8bb3ae85ff9a3dcfe3bf6597ea0022b14cc7d25feb1f6cf5a4dcf9521c019534fa9971d8a224d95b1703d1d2fb0d0c5316cf95403e01cf30954e719a477e9e414fdc4c3dfd439ee14010f786fbec2221b0a476bae04dadbb47b87a43;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf823572f612ae0fce748067555e611553e793586a38d7c774c7fb09546de367ab459c2320f72be51a29b31114d80d2886eb820358f431251d02757d3616a13004bd3f985b9081f5422db7c78a1bd8d629b06948ea095cae5b51acf6d0a68451a2c51bf06e884428f92bd3e2d1ca4dc7fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h232479b6e4e36b89ec94e0d5847524981516455e08dfd45a9bd2253cebf43be2bf609d24370fb84e6110d7192745402c980845c072e525542f79cd452436c4b7b22271151ba8c179edbd29505c3c59a2effdfef2395e3ab0937c9749024b52981fa56d6938ce1af097329b1724e0a0d7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf86e1b5fbfcef9c2dfbb50a562409f7941e21ce65f52ab04dbdb1111c1912ad74c3edd767b6111e08a6ea8e3cf819d16a49c3bf6fa318106ac6206d1db166852923c7781b96c67b50c52cee74a5824770bec29a4480b9ad633886bb1936182931a279f41fe4dd29c28df3548d8915aa88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8ee97a14292929e8e8b4fa3dbdd5f453d1cb8efc8866f192f6118336ea2334e75b85ab39c5cadc8ac6c3dad8cdf297404285413be24f4a54faefed92bc44a7785bf181e173ae087171abc4a82737bf25cee645f63b0efe314d6c172282ff6eece18eb1337099587ccd2a714f907d6cba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha306780f852728e674921373c366e191bc2c3ea6db17bc60b8407f5bedac0da7fc2b299fc7a179482f97a5d88b3fe2d67b20cedb553db412f8f905a93b665dd52f4fd62eae940de3820a12508f4702424fea7220e49d7932100f15e67474c047561e1e90bb65b3f69d0327e77d9203242;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2eb5bac246c27ce06548c5b9e65b1d355797b5c2a4f194b68ea1a5c98b16998c02ee70ebb7126cee86d09124584f82bc5ae4e75636aa7eee594928b0242483959753fffd55edba6c708bac83c86590531215041674de3cd392632e17e223a702f86c1796f3e2d6d96fa860d35110bce36;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h761791bbf85409d9bfa08793fee46abe2fd8f4e55f3312039c8a2a5572f67296a420846bc767b8ca13b0d30d3779770ff6abff41c19486621f05d2a9bc246a8c5cb58db78be1e4ee7f926e55c43e1daf58b376b02c90b623a742e80e3af6199fbd110e679689da020ddee24b5182172da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54545c2601c3b7916b04c69aa74b592728f758232361357fa7311eedaf23436a38abdd829a969050301798dd188ae245bc0c43591529a88914da67f4effd7de756faa1a6e9726620feede59baf72afa0fe315d24ecc1e0072034517604cb22ba7ca2fa68f887af7739df2c4abefc99218;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9d369fd5af8fc0c3633a3f66292e6c5cc04526e282f7f25367a12f218f043451ca7bd4c0f9438f2798e6f1bd3dc0cae0138c9d379da94fad4d7583d53a97519a945437a4332d141d33efc680e0f4da39e7114f5d3687b4b956a19af90523c8ecae08b21bfc8576784dce37b29cbeac12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e1924aefd50728eec069b9903438ac5a2137fd9e059423811774305d0ec833efa8260e8f73c4514578c63f9a9ee87fb68869173c704514337f9d822ddd6a4d892f609c7480578a63242f111bd8236fb7ce3daf1d402aa68c8d622028b693854d3f8087d4a42edc9967b4039ed2d8f823;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b9349f9e1b3c47837d9a2ab2b82b3f8d282bccbcd62982dad2dc683263b07b24ecb54af4b5294a837bbb605bf079b2c88725df0f44ead7bd1afa9477ccda012b07d86b24955013b06136910ea07827f6d7b5b0e93fb0e2a972c0e6686fac7ca184c96d2e268a4521d6088b980fa8ebd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d6405a1cf47b52d8b8fc9474e88e012fd7a70abc573f36bb1345348652c2773c4ad474d5c636cd0afb8df87833e8e726fcd28e23ddfc7e105fe73c4b4e8b75ad6f2c765e679b2a3d4bf9bc7966e2f76e96dcd3d8367a60cd63cae593d236b74b6da4b1c9694cf2f9f14d5514b07d04ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26748410eb769c63aff8d8ca9347a559fe20333cabf9b57d10be534b3cee23a21d590b742b6b95742332faba64a701b44c88e9f6f8f4f03f8d69421d2f92fa97b9c0c9e61bec3b61ec1661c726dca8ff430c912a443cc63de1422b7776ae72d6890e71e55e3d94a9af03dde5c59d6e9f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd28a606f0f1903f3376816e75ea3ac595ac3c3ddf080a892d0ec85d1dff006d6b96c3702923a935cc55ee4841e513eb11a6f3f862aabab92d99c323d9f440e0579d8be183de6961a7bd438d2e6b9ffc086f8b9e764ed4880cb79934d59a3d8963a1555d2bbe550c05b53c645f601bfdf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9b16eb0ddd05d2ff0ac512651e1414395e5aedf00a4c0929b66a2ef9c3cabbb822ec88bc9fc590e862880170df8b6a1f29bc553d1d24b22df8a2c20d16ebe25f2839a22f73443d9d4026a73b18ed0238812674f14710f5e93be5034936cde59ba57ad4c75a0d6ddd909ded5e48a1becc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4684dce99642d720d499155d0c1f746cd7821e2a2b102dd0fae1b7890dc4342278e827c83acfc8edac4bd0206ba8333d3d3674eec4165630571145a2ab43b43a52602ab4ee04ba2dcba7b4c0ac05b8b51c4aeff7a238e91e8ea9ab2b579e23dd74e8cc3fe926e0c2b3e7b688c0d71e080;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfac9c6470bb1c19f84d8fdae2e2b25bdf03c7aa2fcbde702dcfe608d8625818f33a8fe5bd251f320aad0ada08402558a10663e47af1caa9fc6a938535d8edd01f70a98bb62ebc733b12311de18f5d89456a335d41a1f8824c3534bdfbba0a6f0e82a71837fc3a7de48f8582926dcda06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f29cf32990059c710588d2fbd59c51918c0329e68e1adcecdb42f3a2b3c88d95c60530ec187635b72af2ca045df607e841796a764fc5eacad1f7bdde841043b46f2e5eaac6445ee72697c9b9b515c12702097f4b517449c1368b5ff712e164b6a53110e645336c5bfc9f296ecdf44f4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h835dcf57c6846202e20cd6d250d13c1693277b903104fd33f106ca444140373eeed8c2264ed111c7e9cbc233e7f9e02a514e4cc975a1b29cbf750a93bc13b86bf50976713c3e2f1181440c423ee70218d8f72288102ff5efe248d4a33f76e838c9e6eaa79e65170c2685d9c2469c0f8b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha893f20d06bc6350ac9d21077f0edd362b84c46a7644b0276a9fc4dc83a62639c5d5100a18128aea1cd5bb6f8d3f8ca9f7c3a0672bdb5f0599b1e0487510d4182846ffd660a22be4021baf8e8aa2efc7771379acd8edb5825b438782de6f38f44a4748a2a3bb03c8d56e0cad52bf744fa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea71bd6c39f4ec4f2f5af3322bb5e15155ec973ab2c58c89c78acd545b4f9e406b5fc392d610883e7428a8aa65c4158afdb1a75761db3c679762ed3a76a25470ed3aa36657f5555889c2bf72eb4c2434165b7b9b46866de71086c67ca671c9b2adf7e9d1a7d8bc22ce79eb775a273a058;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haccc04b8bf5336f043133a972d942da9a4b6693ecd598cceeb09a55ec6bc8c156726c9be694c33d536326c818793aac0543d015bc488fa14782c6586d3b13e3a72bb946d0d0771451255c271db323893531edce563688cfafed44a26dad4872673dde4eff872ee0211fd0500b9f488b64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2067a42d8a68f624daf3876e4728ddfc9fce91d6f0348d813c1f8eb2df0ee63b935a110d3640642abe4c5da08f07e83635c9fa549d3ae7c60adb2e6a79a2031d0705086c6b907f00998a29049960aeb2ffc0cde00f673fd7c6af33927111352b705344f8eacbed5ccf1adccb9d3a06b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a2db63eee8585db34509bc94d946b925edaa140aabf54554a541519860a1ea1e65cb08e65c2a47be7c8fb55fc31f190474717bd8739d8cdade3b5456555c40889eb783bfca5fd3e0313ffadd3fa342c584d21cebd39246dd195e653d601dceba345c7d353ebbffd7d2d95818c2561b78;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17a8ce334b8f88c8bbab05c6e554f09781f2ca3c71619a5d8976ed9358be48ee533b6dc252e109f240c6822f20d3a599f4d0ae6ba2e1af30190d6c45a70efe1b0b3b5bad77d87abc48cbe03e3d515628cb3f403d93b12af9a80354fbaa049737079bbadb6fa65e76b81f33dd65f17bff9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23badf321f31a2b9846bf754918b8be5caa58a2d83fbba3a24684fb3a2253bf9a68ba9d56c8c38815c7cdee97464bbccd7f053875392eef0e3921a1eab038eac8a36339db21c01f11946da444b6753e42c14b5d0458b3579047450f61f1777023da375b8319c848817240544e3022c81b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24cc196448135544b3442732550eeb220ec155cc19d477611081cb36f2115e2fa0c9f7931028fa2fe8101b17ef7140510408641a5b37771429a750e75d8ff241105a1d5897b8ba06fb8f38f9659b269d8611b75939ba4d843d9d608d801aa87801848adfec06686aea79c25de9d4d3c1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d9a9d66d46d4540529d95863841bc52bcabf65534498fc7c3cb38aee338e6cdf23db2b52c85eb1df33318e8542f024aa44b5939b0025fd03fba55d702f4d0a34aba32afbe67de14612ecb555d6b0774ca9d27a22a3e928c28c4fa3971991e7186788075744e066a6fdae67b06d546d45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d23defb7af5df2a1db8b3c0efbacd4370f8db1dcedb9602b2162b872f45eec5f5f7b0224839a1f14347b187c30bdd729820ca9f52aa25095525f0a00917331ed63116b2cb8bf4e6a90b02f16e6ebdd419559e3cad0b54b9e4f21dac742e1b2e17bf3ebb4e267fe1b4fed7f6871d3a62e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd18dbfb4a4c1ac73f55a7b02df18086460cce895955f59aa56aefec9d231fc26cd63a8bed786028cba23a9abf2d803bdb258a41841629307c4b503b13ff85f620828135a07d2b216bc92b576ac55bed6348978ae053dfda0ffa55c7a174624a7438777dd23a76348bce370b81d1e3333b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h381768db0e559e763efb0808e638a6c35f7a64260b558d946167dbd7fbd7bddff4052c98b17828cc696fea3ef2df50152009cfaa429a6e6d48809ead004ed65ada939b4cfb2d0719a19ae7717879681fe3c34aad0406164ab61bc726c6cca938e9b6500ad89d9370c15d4c7f5801578e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc597e77ee757575772744f405d1ff960d378d809e1fef35d515ab6fcd5f5313aef97646fe892fa8de16da9259988139841f65e53fbcfb03184ca5cfc999b4906029b90cd36f6d7a675bb647dcdd3a44284d3db22a5c8ba9b661cb1f33c7abe080e370e2877f8174a5ca18b12d34d2bdc7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74e44570b3ca22dadee0e0f6aec25086b84a12e1f0d07a23065054b9f2df9d5d662685dcf09bda6056d6587ec8f7d7d21b85b45426efda273a2966e763364c1d2046278a953953ced2ee83ad050a1ca7f177e8eb147a274b815a3dfcd954c6eefe80f19c6eed8ef6358909f7bfa5d1ee2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a7fa387852ee677585542a63e04e07fce3fb11d6892b1bdd6d45969d7d72fece246ba7975d12eb61f5bcb5b524d233da3a857eca3cd7f58daba49ca0de5399ceb1cd9479570dd132de418c7476e7fb7c261ff3311709c206e242d28e9392e048d86a3c4e7767daa315d7923c418b6be3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7179a0e1a3ca50751053af1ad6915cec7da11b7ed6f564d5e2292a0f68ff151e9c3c7d713a01d29203f3b908a0d6477a97d165d9047afdbd19c2feacc90d27525fd2b37dff5930200e328e58228feb90329d8ce2c2ce34fa3be3ede595eaad15400315137948e07e2e5ce4e134f70ca2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5e5d4bf665baa1a1839ccc5cd4bdb9c7f8d0b185558d7e0f5576182f22ac0ece9b21eb0cc3f0db7f7125c5dab5e33d6f031137590ca2daccb8120b5042eccf48a13cb7e5c3880c04494a87227198a00e3bf4e135de65addf7df98c5e9a8de947a0dd3ef139b245fd68061c8ffa9f02f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7da98c01fcf4c82b5d30188b0e3cbb78946ae91d90be4cf8f40fb602d02fd1480afcd6dcc6e90778b5b83d0ec2316192c283f07c4d14f86644f44eb4e06c005e731202fdaf765591bc0f94f58d6b314fb0aca962f84e70348135b84f70b3476644b4ceeac7a999c53c9c88fb084ef775;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4973db5c46b0d592e050e6e336ddced48ddb72316d5745b047bff0651b84c66427bd4acb386f5b034d476d5515907b9e0ff60b9b0f2cca1a91ccc194f39ddfb79045bb828559746d380b58b79a8db468343b1348e7aa98520059f1f59863738eb75d38125b013b249ea3b0cafbdfc2cc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e33aa9201a2e0690d21dd77f81264beb3cca6cc1aaf6f7e7c4a8ca7f5693e95a48438cad177610230e85215a5dd85a8f535b796fbb3f282fc8c2f6a9db17c7e2a5d770cf4eab5285e827e15bcecbe244374861a390158fadc026a0f2fa0419b330f647e2598ee63e40529541b8103389;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed7521f9f47f1b5a9950ed31fa46e2451405e53f005b29134c31960ebbff39a12d50358ea4125324609f1be430a6351a56d12f0c5da001105c9b3d40fde70401f8c743239590ab5bfd4402f39ba897e03017a9d3ee62271c43ed1bf6e2be0afcac62484b5de5fd137df4a6079564ddd11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9930e8b403e7d9a643abc9fc13c2a4c7e581c86958ef06a5ffa119f10e7aa2135843aeb905a6609645344768e474740f1b183f8a79696e2247fb95ad7bd923b8ed47f2ad9146a498c282fef37f79161da8cc9ec13af0452d0682c5959015b437243d43304de9396c0ffecbb1ec8ad93bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdeaeaa04a1fa772c47a31aa3f583fd332cf3c8b093e8d0050d63808c28531d171268acc1e79b9f663409b0d0caa77d2a242411a8e74947184d1813a861ed011f4b206f834cb7c011966eff660ee3fcc0e5942b29f92e7f109a390d4a19ea761b81b6218b9c2184beace3d8dfa85e9063;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74b05fde51c8c793d8d756f7f01ec3a2ec1f5de449e3760772f468fc32403ca5887d1e329b5c4bfef5d0150877a8125e2f1f252c1e5d576c228e32e3b631193ee2838fb624a69a180fabb20be7c33606bb4be99d65c6e277b02510a4f4c6efcd82044cca4e97b9151e966772398dd7e3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15269e4eea436c3dbc2a19f677d6d3f0afa0f376007739934e1bd7d4f25aedfae87f41206a8c324bdbb427719d3c1ff1097f186c7f7dadfa18ba3c013220a6c1045b7504f5424c3fac1c436c15cb6b84fa4324457940773616a03440bb5169f93732f8a40bc7c2324cb4a0c751196a79d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h280b3812f728f958da59b01c66ff5e591d9c228fcacbc559271abeb08e9fbc0b8befc7dfe4a799adeb491e7a5e4193229bb958b42c8b69cda197c6f1787d008bb514652d6c0495364da2a75c8ffc54aef579ec431028bb99328183fadbcf4131b835604ee977fe47141a28845c326fece;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7f325980c101a0cf4b2fc6791ae99b3d2c1125879c49acbf2fd71448d597484b017f98cbbf5e17e43d8a840e06e2f13a1bb8fdc0061ebd1804b5b0514ab86c2eddf97e1c280bf3fa8987ce55fbb22ac791c47bd661caafe90a01fb8cab9087b6b61c70797f64b4166a6342ee86b87c05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b5048670f3c96fd616796bb8ccfd4511136a1c00ce860244e90382bf45d8c1a709ecdbe014e7eed9657606c862cc66b0f09fc8830b295ceb4a0b214aebb2c407122ed3e6d423827d100584bfd4763e6b40a730b25d5d30252e67379e36f540a29249eeeb07cf6effb702c150629ceded;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6e6aea291303e7d2f3daa724b4a31e2f95b9e3ed0ced805df2fa6ae918056781b1bd12ca6148cd0f3cc86a919790d2263571897e38cfe1d1f746bcb7b2320f77d311e4c4589efbf04813c9411fa2b161912e5b83b485798deb09def0b4ad61ca1b37d24be46a9dd3082bdf6516020f7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h204dae34fbfb7720470409ca9541cce3f9e5fba509b55bf7a5e9d369eedbe4ac42e4980bf17b1c7d64e04b1754a387f9d61789e8d74e502867cd95675376029b8995c453f78618be0ff833d6bbe353dccca3c5e987f7185660b6b824950b354f2e48356318464d96a40f7d5684a49034c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e970f54f59c455043078fa5b374fd1adfe247285e204e566ea103339fdfd099181bf23688dc90673b4d7842164eb28770db05dc6aa319296499b354ce49ad61fd309adab6cad81a166d411b1ad4ab5e060cfbaf4de3cb4fdaa0b3e80546e4bf086224f70e0bf3e22fbe1dd540fe3df36;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8615ff46af82e5570864a1a6e715244d9aa0e9936125cb4d0de8c7cd0d3608a4aa4af4e788bde64c20e6d939174cf7650e9cfb2d60c773f85e810923c351aaaad5a7da229464e84861c479449728324464a384d446e9bab250f3b22ff0ec1983a5d36f37afac145974c21727d791901d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hded5c7e52ee6972dfb448e5fab77f7f7ad07e952f38d8c831f014d8ae8be7d5e171547408947e75e0d64689b128f5c9ff15a7af9e3751357f3909ff556f7115997ea0e3b6abb44d5dc6bfc2452515fd7f47938f74a6a508732c096bb95edd4d71e6d0d8d48a9e22c643fcac81928b640a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0b7b5a1a01707ea0c21b3dea864c5783d556658dfa26bab0d4c9f72410d0abf70ba23610e94528450763e9198814422647b5074e7d6c45b39fb2eee9f4dde05a3358145e2614585e1a14b7abd43335e226ea3089416c291ced2c1f58a4d678018c273f0d83d622d173c93939f2e8b34d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd255e5006f9f91a1163de91ebddd64a3916cb971f0a414e11f42ae3976d185af65fdc967c8c9aba140889cc2cdd51241bbb78f0a7856d8c244ef6112beb7da9783507d3cca5e64a60a8246b32a54adf0c2f085d60d396a100a00e24b61b3aea4b9d14f58aa61360457b32e4c4b37a0fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bde4660962f57677504731c5fac0a10746cd01543bec3e27f8c2edbfc50bc5fe9d83c950f77a6d45694051083a5db72269581c8e0fb6206aa08225f53458fafe72f6379677b5780e2efa7f81dcc695bb1431606a8b6eb01d879037d30a05c228c80c57c0f4cc8bbd681743e5a5c32969;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8974a79943b2a0a304394abaee6d424157cffb390c7fc56482bb83f7eab1b188da363c15ec379f2bcf2bbd5061f2da58b702f604d5df14e7f895dfec9df38705641b328ec643ea5b27d591051762a498c4a6b7ff9bbb78c89900c977074602fde64187706923392646eee981bdb7b301;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d8511c3cf06595ab4fe2885b576e6d50a170ce84fb59d13ec115406c6fbab7b23e0373ca4ec4225ee225b3c823c41330c7e05b7634cfc274f07a29df3c4b82e2c4e6bd779eb32f092a3f3b1e602bac7b6322575cfabb7b1d227a2fb0cf30a686474436a11dd9cbb3d1556034155e01c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a504f3883b33fac79052eebbccad538cd2ef44ad84be494c515c0207b66691d21087da1c2413e4989fcc3f303e9af5cece0293c2c6ad0016a4fbdbbeb9007bd7b9d5a91f8ec7e3d1f6aec200177be1bf3256365581b78c013d7b824e64352313f681fafa300671504b10c2dbfa992e6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he17f3587da1fd861fde92cbbb7d04dec4da6ccd687c213e0b7f4aadae86bc902d29d9daf58359cde298886bd26b08a98b9a8b75772b0d1f3c0546eaef7ce0188ba186a9cd6f450c9086f665a9696ae5d8d10d22494d054b0dea8e5ae14eef67617cba70dd57be2177a73fd5cecf1a3c79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84ed616d49e9784973b40cc4fef33eb50cac693b927c280b177a6d5fdbe8945dccb62aec0e2577c3a07b6410d6eeefb81a8339ee0720f42843138678e98368c0549201ef4c1fcda8785a12fe52c06e55535d0b7e605463491ac084b68929013c0c7478cb50cb2c91258715af2f1d7359a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab01d9ee6e84599127529dfee04d8cf10ec2c509c720c6c9755876a82751b8f1ef86eaf69f1b8c57a00b51decd06b24e8efc6f147b01322ea4d7956c974360fa1839e6b21867b7f45abfdc3a2bad311fa4d40754e44940c845207fb5df211c77e4cc137fb6f8283ed50da6e61fe2d0b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb213f2c865807f23d0d34146f645512005444218bfa17d5942cc4b0bb1ae0e79eacc96036aba1e6aebb9e04983313c9b7c04d19478a7cf8b21190a3deb0fc4ea6e735bb26b61672b5f5c0297516c2900012e9b06e46ef2b8153f50c92585f677ff037e5a675dfbced8633d7bf7b5ec7ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc41f6204c27ffc8f4b8129531a54d0f76d027e67d5a6b1ad0914f8085bc2a466b445acefc29b32ab30bed02f8ac16efbd9e4b85afe718924aaab546476920fa0a118f661dd4327002a01333dd834f830f55f2423e9707adf90557bcd6377799de05c76e3c48913726186da6e3ce8bcb27;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f8ba5c60e2cc5e18ccb50e4edd8b6abaf8603cd78220d3746cc8534860f1eb87f64b5193035ce875480d66bb81ee05564e103a457d18de430203865342295e7de13f9108b5362c165c1d6406ddba48348469e2f19c2872cf1b8d429b5ca50b846e6cfb955c11b05a657c34a7d8649b61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb09c2eb0f531b7043afc9dce0dd5e3297e4417126476868dbab0c98c49283e4ae5186e24c1a34602b92f830119adb0cec74297997dbdd443d72ecde4f5a407772fa68a4d7245d90749984bd3cdd346fccd4634b8ee6ba1b30fb7d8c55b850853c7f8eafc135d7ca6cd7bdbe5e1a34b67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb09bd00ef44a48fc02d8c3039108805e2113f63360eb28d4c1f21464e17385a7bb86e260010fb049662388a2b7222599b4375435fbce86ef0f99e681f1e517a412d2bfc505583232a57158faef5c798792d47545eb39d200c8bba794cfb42c3b44f52cba7f85bd26fb66ccfdf1756f297;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44ac40f2377574130d71c20fbb2358858b0a72c44b9524d1623e20b13a7b8d2dae2480b8e56d917f5826147e9d8653d4fae17ffb8fb8c4736361d1ff625a64e339d59bed5af23cad347d7cdd440b184530efa92b47f49c6305dd24ff466b84be36040bcd977223dee10ffeca1af87737b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82dee3534fc33960bf7d721c8e7240824093c82ef3aa23f0ea30fe041a155553ddbbe59ed72bc0e09c8473770af4f3bd1ec8285502f427b7d8153e4b1f7575489659944f024aa828620cdca481047d56054d4b61757f204f485d315d8ea6ff1bd3ea649ab3918cff305c79d6c312f2338;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf829db13349427c718c536a2b60afa4fc5f0a9119126ae0b6298248d47a45c17bb758b97bd9a4e275db6ab3a0abc1cf51aca9033e7fcbef4f7f9b7c69263d3746a35c432235fc19fb29d3c0b1a08907c316f482da1bc4f68d7debf9824823f6dd0568bff1b316bab224d6a6c90c86ecd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebbaa077e737159e943619026670aaaf44e0161a49b65cef231d2029a1b16320a64a002d705e8f40a8f13bc86663c98dbdc8fb87c4e46a786ccd7c635845d11ac0bf64377d151ca3f8acf1d66a7a565d29b7d13ddf5f74d1ba9b297bb7dcb0ac2e31405d07c2206da59617c6c19266e41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae7b276c204e62fdfced660cee7a1a8a383c2c5a07058210e5cee05786c0b88463c3831168788a15915175b4c350fec4b74331ffd4624ca8005731f1067df4b1afca7818a4ff6f4feea0b58e4d790764319b6b503ba670d05b8579d5da54cbb691a4d9b0d19d384ba910ef232d89e5d3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf284d7174f872fd43681e2151659ef8dfcde31e9bec471689b02486a99deebcc6ab1633021e9811bcd89aa514b444b603b3624c09664dd79544b2b74dba3fa0eb244948ebaa7da4bf9ac319d46c84c31230ad26e414c95c664e7bc88a1c1cc89d506ae524ecf960e776674f65bf429bb1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d0e8384a3acfd0aee436dff2b0ea0eeb6c77d3f7a03adad6e9c6dd42f3ab9796aa4b2d8ddc64bbb982ec87484968a39676d5387379d232f2d255badc69d144f8c6fc94983ce8f06389f4536ef081e44039f732f807b3a76c5c8599d8d5e0f8cb2ea5e3c3214c63408bf963dd7df0c061;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h130cb422490468390e6d88325acc123ca056d3b3baad94a20841657b9dda2c622366c40824d1b4e78ad69c2821044ca62a35a94c96acceb90616a19ecf3d12118e86a3816193253f2add5d7ff5e5736b13fb00537c4d4fe490ebd8dd95eb6ecc4f62f52159266085fe5591b65eaa77ebb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef52c8eab18ca7f41477bd75586e62ab615f601495d1b56b1ce22b702ec7f16d99e6b6e564dbb61c2ccd9aadbee98d58c0986a3e3ab3ca7cea51f8c6b5f812993fe0adec6fd18ead6dd5e85df55a7a19c91ce4257e99a0cd5fac91ba047eae5d46c34af19eb7f5656fa4612a647f75a38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e4169dece5fbaf612cbaa54975252e632bda209bbaf3bb56f2729c8751c677172f57ea43b8766894f6de2dae6fd95c8494684ec3cdbf0079db1f21693a93700ae6863675b633c90c464f10760eb5d80fbb5dad8dc495b73bba4da9c4a4330863f4e3f7070b03f2bb060959c8d0e21699;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1479a826fb3d864a6bf36b7bcd47f4859f2b0c2d2283c41b27138d95d5a05bb8292d54335746df24332ea7bd22dd2f37255330b5bf887c756815572d2b5d2afe82d6beb2765a3093ffb2b1645d974c244d18549ff9c7c4fc44d57c708d389c37ebecac1b20326e68a3226e2395056278e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccf4d83276be75b00ad78ee5586cdafd24908b91df293ab7cb62a3a07be9db3ab026755352b4deafedaa922050a12fe2225d689cf59efb1cbef20d16965378914bfcc179f30421a618b9d9e6298b0259c2869226ecfe7532f3a9c8303f7762c0c2f77546196725690c3bc1926fc19ef44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h898668c1763049f976defcf30060062258ea87602543a7d8f85251139bd1b1d6cd19227510cb7761c1681053d03d2302ece6bcc4062fd9d78bc209748bbd5bf8cf94bdb82225762f10f7d7abbaac12118c3449d27057bec12573082b737f8d54d8ed998d01688550cfbaae3f2e920792d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7d2a4ab72973925156bd55a2deaca30d77647661479921f70a6658de8e5c103dfa75bee1fe16b9fb3470bb7748eb9fbb7c05426015160faa910f1a870d5dac4e4cc9e3725be33abf03a0f4d4734a67433c7dc5d922088b2a224f09c0b6f9a59cbb8144a3da697a3812e0528d417c851f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a6ddbc53615fc63fb1a5252f58453c99de3cc9032fbd2bbba03cc484e8e3c034975532a9eb5490b828e9eb6497b028a8ccb3b0ada9bd75e7300b4ba74f765da5a46dcc243c21cb031ae0be125cdcffb9c3cbbb708645c409ef6e7bab8750395fb3c82091bb6597cadb940eb626914e77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba18049589029bfa646bffcb3337ad91bfb399b8735f44619a4fb0f9c90014ab6723dae057a1049c1c79a71751127e8a7ce99dddba6f8a2d978284e53fc4f75df09b1a82f84ef762f5535d67c05aa2bd5f5c1164aaf27420651af71845a6fca2b746524f0f38abc205b9bb010719e9af9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdda7d053f9391b1e66ab94543c7d771f8f17cc5cbd06728824935de07dd3a25a040bc9257f5c44caac3aa27cb4c69cac0f00fdb9180881cb645aea8eb5536e814c84d8ac7491c72c4934207124b7cbb8067fda2c925402bda500c56ede4718be3419d3de1be6d8def89e550f1aabe85c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha046159db3bff8c1d2bae1910945e1b39490eac39592df09ed96dd1d24aade1d6bfb90bb6458b69dd9ab46ae5e81fa708a31b84555106c73cea2b69d3b23a9e15cc61e5f7d9eb8bec9d663ddd6e7f3e930e6bb0596bd849650d870e556c8e7405a21985990c9a2b986ff71dbe63472be8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c7adc5210bca80a550a5d69199747abd25ef4ad6f48323cf4be1263b864dec9a9821805475514a35336f45f7faaef647339b346b06b904073608b445cf3eac30843651810c869a3bb8019a82413bca64dd53ec9d98fd1c084669d6e1ac70e37739a8bf29eba42f69f2dae172b3197e72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54cb9ae6cf9a44a91f6bd5a9f7ccf95a1a09d0241959033464790dd06d3a77922adbfbfe410bd8e6dd75cc9a0dfb0b910dda49e73318be9f676e98fd00bf65d3df8c9d16d23ce4bf08e48b81b06fa796b8791ee9897ffb43c2a36af6eb250664ebfe2ff5fc5c3992994c4fce19aee9294;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb72788d2eb732842b577eb61f772bac2cc6f9224a03b882c7044968bf3b3df6a2ef5aefe764aaaae28be3b62f8fa51f6d04239dcc02f455b2067cae1c54ae26ed5aa7d1bb3e4457b4e561e0ffc3ec44768ebc322bded376328bb3a773031a09881961928c602199c908d490afd140ef2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h540418970179ebb66f00e73c4fa72638218c8bc3a057823510c3ad4935e79dcd530041db7e2158678ece14dac555daaae5e4989744636d2905f07083be1299da3a2ffeda43f4de3eb473bb090f8db4e00c20510e8670df906e415745e60a718ce1c25f4e00bfcaa52a7e517e5c79038d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hace769621363b5a08d29379482ce78f39f5b9be2d5dad674c92fc21f68073da6b51abba81d2afd09d3c1baf3f16bcf1eed70cb95e9aa0f99daf408a5691bb75888774b06ff9902cb7597f3df1693aa6694aacad710cf5531a2ec92b5c20f458210271ab283aeb4f3b5bf9f073a9ccc91c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdbe4f61bc39d2f3e1d36fa6b38587b0045b835014916aad4efa9cc3ec2f35eefdb6d21ab62d94befaa1c53ba2b12232df6216122437b652d3401125cc8cd29d9578b93295c9d62f8e925863cd3fc8f2ef2b8df644702a9989cb18459165043a13b28aff707c45e8990fd3f07f4dbcf9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb98db9830278a891c0fe6bb62ca30ceb153c301b318ee4a8c85d59d38dccf4f7a0160df862118962cc511f399fb3f1fd13d27584f2d5a52e8afa0efd673943bc0f0b8f79e0a259e27dd73025ee069c9df427da6737f747b03008ea400ea51e0c41feaca48c12a51a88697e2c85d6a1345;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cf88a42adc150c34bbfd972657e22d36bf7a3422ca4e91942e0dadd0f6b858ac06ba3f27227227b9f7f68b18bade0d67f27f0ff14aea6d5226f4195f03aa6a009e6da88b109904fb0ab5963c29ad42e11d247b81ef248b97257de4279c621520bef33cfb91decfec43a1f49bf6f9fe98;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h256b345418db2d8ca8c40e3ee4caebd20506a55f131f17deacd992f5f90f2ba208f195cecf0e565549a83b16b595d0e3342d1aa56e44ff4ad458e91dfd59a0f0bc3d4b1db8740d8d56f1877bf066dc21a0ee80fafa9f44c447725b004b22189b93a7e3a6bfaf3b00cf46ea7ab3537da81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bb88d0671d6581f6ec34906724a4cce55e67f52d5b4e5369681603c36334d4f06c152d60bf745c25f2819224a2cbe9bb9cbf18df1cb16ed75825df91684c6f1c77c03506068512f90cb70bdc7b2f3eedc526edc826406c0d228e3a9ecaac03a95f10b9f7149e893f2ca8bc76f7963862;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28c8517d3fd206e4d8c7ca2fc03528b3ccde108307543cf47b4a63127a2ec1318f268c81dc844238709ec7aae1fbcd5e06ad5650872e4a398dfdaacb213db9535fa21d5f7368dbe3a970b79cac4764aaa64fbbaafd12eabaa6cf18742a1f583a92d5e1657476cf2a66898310f410472c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45f278c147cdc66415f18c017cca168af136361c813809323486fe9ad4ab99021a6b136aa2603f78de4674344311cd78d4499e9b87c614197cf61589a5facbda5f407076e3c9eaf246afa91cb26b56bc7a00233a3062b87363c38c99ee535c811843cab693b29219ecefa128b682399cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb964bf5ec5fa157e9ff510d768f8f1fb15879c48ab41bb74af9ed259f9932e5d456c37399b82637839701c360f283abcab0d17515f4e99422789ddd600665809fe2cc3d879a4425744b389f87989548a125b3b2fff4bebde80deacff690a6bac4b7a040784fe314df99a218e295bc6cc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4afd095d970793d7825fe31a8f448ef5ecd345d86bfaa237bae8f22c76e91d6192ebc65467c8a7ebe595c69d9d67a2cb32e4c7110a57289796305804d73e480f67affe5d30a5e0503b7eeb61fd229db3f832b2c4d2cfb1288c2f28b2ca95ca74065f6dd541196bdab70581d85528f215;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed48a6359e10b5fa505d922b899d71b89189fb54cfd5e94835d8e0f817fc455f354e01b4d8388d2871e63104bcb6a383e6d26fda0e31333f5401d85b34452eac1fdd06cd6e979b8076ca9613b140eeeedd53a506d2a38126083b92fbd114a2c83cd5746a31a5394a62e1fd2797da7ccc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h679a64368ddba48c857e39db83184f697a68ec9496d2dbce64da178043c6abc6b999ab3c37681377322a3ff7768bf34029140c087e64c57cd406051b98a0350909b593bf598badc65a907e8562cd39577df808621434c3b69e5857aa81ed03aef800759f20fe626207b1e1dbc530afbf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d5a782b40e26a5b2a715f64e8b998fb51339a1c2ddbe6e5e2665e6f159ce58944b391a4173b4cc113dd5186285f52804886e733742786b30bff1f4a8ea3bfaa8180c9c9b750e091db313118f7c0306a098361f5714c190628decdab0b9f6d13f8b887f82d71490187226063b8839bff0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeb44bba5123ea5ea014d910c3da42a01aa1dd400da4dc0b144dab8757e1fcf7c186b32e4f0e3382978cf9f9d06b0b462e5b43bcb13b6bb36ec0b53269a1c52ac12c9b8fa758d65659bc649684cc798dff2e4d8bfa4e97cf03fa11496d60b0d7012b7e933681621f7e192bf5c1e061c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dd42c6087be5a0238090100275fbc35be8e08f6b93f2c5707d3f6f47b982afb33ab5f2ea699f3c79cd7936f30f32737a5481183fca2e19a3338bf40161539b8a12281d53fca96baf482e0c4a111475542373c4871ef8edb55448c580e19c8fbe18949a63a2c120af181a1bf9c9fa589a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5a055f834ad93a9a000680f2c66b4b82abd1ab963061163007c782065fc6e29974ac0424ccd53ec230a00f449068115ca0a4056ae07fccaf42252350ec0cd3f7721d12918a7162902197d96deba45731e3cf4dedcc9f0ab819cc86208dd2c6e7a45934528c4ac16fdb4224269b69a9ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3ac8bb01461f58e091878cb4326ce32a2fd38d3c61f1363290b0395eb19f512ba8d466719b2fdbc6bb400c38d7134de96cb75b6441135bc87190132f9b3d80eeaaef3791130b08112bdd069c94a353004aae0fc6fede0773edd06524705a030153ed0de42abfa8d0e26438f99749eca1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5187a853917f8b599d689a907a695cefb71809b255fbec24d0e5f6dd94e0bd980a75dc9809c0e5145794648c95249ade5ca09a6573799eb02312bed10fc2d90a1e26d9b4cbbb2abbe649fb6677e327caa53e50770a22359821844ac800646dda2019b35932def50115b66220b89afc142;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h289b699e5feafd87a51564a1ef80a6f5c8fdcc56ea661261120d3d6784c3fb252ab1675a1f955ee60f475f1521fb50288ce2b7867b77eed8c73f27c45053b221a960ece4eed8d63ef19f6ed5f5a787678d97b928e46b18138c6f63055f92327b73ce9cce7360bfb60e5f0a6aa092b5a84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heab69720ae48de6afdb3981296b0c9f0b66c6be66878fb7ac89f88e955103d90660c96d4ae309285e00659da9e9e3569525d2f20fbca49571172870232933d9540ea403b7b61b5930b0235346bfcb27ac81eefacaf935a7b2d768520d64c890db8a861f97eb372b002c6d89bc13d4132b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f4febd0f1a5ca7a0e243607ec403eb6368e68a3aac788be518cf09bd9c95843c759ae08b0549dc881e860ca0130c47245f8e69d704768133d0ff3bb4ce0687231224e9410a958d2799223c83f20faa8b88d86d8278557fcc656c9459b2db9c4543d2b288601eb5392fa315359c636a77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35662b51581f95f340e3049aa4f0a9f2c1a37305a9220d74cb3cd780654a93e120f9c155c212d1b1ef91f82fe17ece4adaafe3bf596464a54eee09a9c3aa61b3f89eb5ba3493b4c907eb7d1c2d3c5569ce1b4ac2ef8c8b41c1991e227094e96c3d6e65e97e528083971d5799265ce65c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4e2e68fc93ef3b8abae0d822bd6168396b6084af0ed8a4e6503525f431541ed121b96141585d7f52f656228986e9eeaad84174ab069e70289f2f2775185e0ffa32a2f23d9b6d8164055e6ecda8b1dd3dbfa190252029144a0dd89a400ff474a79b0b468bfde61be787bea7db4d4125b2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e0875de771eb360308037fbeca46c21d31820497ae8e470d3081c58e759c1777c0753660e8e2239068aa7a3dc2b114b03ec1f26b2742debb269f29ed67aeab289da37f4b9fb70d74995c2591931c7b7421353f335fa6b302db6d72644a8071a42bf51a49f9796007eb5547426b0cde02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b3c7b15828a65664d54eaa52b00a10048da70832af3740a43f275b857753b443bbc066b39b0f3cc9576862d601e54138fac552939dcb4ba0932332f1c64d94a7c3f0b0906c8cc6fd7026ce1a74014d30a211b3f170e387032d587cedf09c07b285df68d84f62113b22bc415bd8be3f32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha35abb523f6a168b260e9abbe60edfeef7bf4a251eec29a244b7443467dab4fcffa2ac130a9a498ca6368dc3184958a3d5046135f3fbfccfae34e58990dd1aae2a7899fcaf01f9508130ade4c29d4077076e0eac09a95ecafa8cc548f2884892d3c62bc85126670826111eafc073ee80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc07d8a77411297c43360b3fa79f702f25eec7197ca60aeb5ebbf9a58f057c55f791918aeeea4449d2c35f4f8e5d4f54a37fc1881283414706d614a8022f0cf927953f580c97874a4647bf82da50fb35dc3a7eabfbb42378c4a898b18d121bd1ae0a05020671da4d1d0bbea3a469737411;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bc26b770b8270494f5e70ba04f288523aa601cafd6b8a77c5286424bf2cc2d2c62462a2977dac4f5cf4b02ed50e9cd032121a761547ac9bc3814fe6f476dba7dfcbce849e57dcadb11a989913e79501a0a90c6e27344345017a70ea7cbbd67f7e57b55a741f25a84110cd56c4dd53067;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25c757ec59106c60e1e7eac824617456625baee6dbc23ae98fa516edd2af59d34903b00635665c599fd99cad5f96ecfaa6ea947bf9a8fe0540ce82efaf70079719344e10a8b49a97935a9db147848ba6e896188656312be3f94e423df0ea44b8ad404547de1cfbed48e2a76c24af59205;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfff11324399ec98d89dbec47fd1e6a1abd435ba89de5f656d3b92151d9a993db2f81849df62471ff766119854de9207fd8fbe38a973b56a35073af6457a6b5054ec85f32b4d1aa40cbd8aab04cdf8c54a9ca6007b451af72cb040f9568626f2a4070391aff52adf8c30e2ed30dce83af;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h277477e6245900152451b6f9d3076a64260a12774c5e8b43fb89677540859c50fc7db446f30963fd51484c6ffa3899841bc05e3b360455136260741dc9aebf0cd2e458d18ba247347caedf109b10513cc643ca6c682a97c53692fb5a527f949378dd01e362ed0912ccac46e803652f091;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54609b2fecfe414f45d6785b443beba74d239c6717d028fc5bff430c33de88baa7275a1f073850885ce0003cb684d2be294e3b196dd8eff5cc1b482d4e4c35f79b0f547fbd8edb407386ccfb8d166373c570e17d82e429b744f028b0d25b20458519cf53cfae319b3722a6b2290501e43;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83ee027fdc2426137dd7ef411ca1d9b1fef105cca67333002bd42616bf291e4a1629317a27162ba5e28d30184a15e0da0dc5562c390b586575e0bb71ff87d69938482c26a6a21d25b46167fcf1f3b043942e06c68acb113a9159be80160f2460a8b545d13acad8b236eaa2a3a157a7e34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h623caa55533fe305a3c69b2fea08732768aff3843061aa27aff17262efa71bcccd3ea65fa465f12bba956a6ee4b0038e6f8ea3b95cc4e0ab3e4f558e4ed5d8be72e862ebd7bb44ba0b007261aeccbdddc5412c624183a100cf9c12e9bda52fe4edf7b6bd8bb08d226161049a8e47025cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f1e678ddbae7c9f473eb83968b968e1797254c5c0e9620fcc24a89323df7ef09f59c689ffc8b62451cb9d3930a5765136e8fc23076eb9a2619713c48a1b6599119c818a6c47d94d0a5d190741416a66e268690bba9008de831848b1f2603d8637d5c928816f7a8d5b70e7b5a47cc9a79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7363cc533d9e05719ca026ad6b2bd404a5bbcb0320a2c22920a0912dfb3bbf926c52efacc60009fd10dd5bd3dda3b3175c7d6d112e584e7579b77a853261ba47e79d17703469633df2d73e4064b94afa80da8b8bf5f7ed9d088b11151651059f23b453442f3ca61b47b051e83c3a2952;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fe90eb1c5e84bbc3bfb1bc746917ff39f62f814b221579e101b5fef81e8842bcea9e6343ce40628643d98faddcc6e5a33e56e18c2cba1b2fa9ecc74085be4a8f5c18df23b073409f494b5d1c783e0e34377b59a401a745c9075e307033adf87155ca37e24905de12e89a3d1cc96ac367;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fcadb96751187d996c45995c3bd7397cb3c15e49fec3728e565474b911c36e6bfcd6884437226f0e709e8dce407df4bc9e8c95b4d3210cd3973f9a598de07777a2280bfd7dcd328c317af4519a2e88b9134af9c890d7ef9e095eb1261d2635b3035d9500791b9942abb3218cdc150fd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5ed518301091b3f48f420e20cdb59797c84132fc5b865868017f817245b769559e9554ea73861f89bd9d85b00872e0cdcfe5aa8ba346b0402e0599c9a0e2d7421b9eb085d3e1544c0bd8236ae9a00ede894a13c576d35419eb226dd16095e5fb3ea9a0256cacd6ae8d31e8b6ea719906;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5884305f46afb8b766d2f1b03df3babf3c0f7f2b6b0e540c389c8f525bf4cad8681cc588673fa9debc0a33d80a04e3cee40506bb4bf0a7445b878532a1c89725dfb85bd40bb29a56c074ab48e949b8db89c018c69f5467fbd22310a18c55df4218d1911101ca4df16f0536cb27d53b22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32fa33302eb8bac6b5a5b2893e8d7730a295a92ce29455d2a63c284a0be295d244cbd572456bf2439a49723cb3b23ae59cc54bd90af2a866985c5f03f931da08be68048add293633479d294de019d79f99bfa03705400ae13f4204e3a466197a8ccbba05581da6b75e3630282a905127a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h871599e6248aaa930ff11f80d0672a78133f5732b8df438af16c46b8f1941c6ff6af07b26c3bb8b282f53b3751e800085c29b17394ef231ae6f9443f524763ce73c49a8632a52fce307fca3c1e41fe74d99e62e5ee20fa9a9d42cb77059f6cf43857253e48c81ef8fa9b3ce60ecdbca6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbef4f808c48dff598bbc5ca0ebc07df15a99c20aea47b256c3de971798025c356d9840a054aad777d54089b6f53945f2cbdda8e81da0241bfbd45375e48bdf36daab81aa862f15fedb67cd4c6812c59bb368740aace0a6f40425c62201f1ddb11c7fd8df014e4700558ef598046caa5bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3190c0d320d33d8f85a27c3f057e57bac36765d5c4ee8c9f8ca9d46ff73dd1a6e0d5ca8ab43ded0ee7ce742d9c44d3ed2c2c7c398163f2a0c5d14651dc02433c01958f00b27b544ec5364198a2dd8fd92efc77d11274e649552398c55338e2a7f8478be48d8ad46000b088b36b128963d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd407c17f86bea3790041f82fb3e98f35013c7e8d7d8dda6e14f48fa2e78384fe37ae1eccaa737bc17751c9b9e772970d210f4b7b413026f6a78dd31cd4fcd124f06f923c9cb022af33a37c9d71afff332485d26fe16a8953e7742723311af0d74c01b9eebd0b3f6bc28c263605f2619bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f2d2479d417c7932944238b16902bc39e10bf6d18ccba90078a3e519af60f9167de9c8bff04044ad17e015961bcf9dd041cc9546ac93fbbb53c8a3dc2bd6d4a158cd8b2a53d390baaf0639c039ed1d74aaafada55ad51830d3e074c9400097341a2b8167036e07421d48085c05abe49f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dc43480213d9dddcf40b580ce4c09712226f0a7fd0c17a1ed4658e4fbed24a63d6e947b937abddd079190be50eeda744f38a265690c1d0aa403b11b73b4695d68eaa6bd67ff74fcbae4c646c52b98c93b296273832607e239599d74a74346badb665eabbed2fd486f2da00d82a91f4df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41d524126ae22789e8527eb0cc4f5161092860ca1323a48dceaa70b309b19b1d4241b2ffb39561251c6a6211ec0286a21c5007700d8d8160d3581a73de635d5b248366e9d1095b05665f45e17991e8ad9536c624e513e1659752137ab43a63500b609486a00e93ea17afabe102eb01992;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h315b2321eba73544cf8c0e80324ab3fcebc526502b5ebc74d045314a241745a8f1923eb86049bad421ba18b698409fd17f07e1ccd0d2c4c96406c8940c556257e66f8709f337b072ddfa3b346ee721d713b86c04a350afaa924f1eb43dafaaff4087a772cbf4a9bbc061aed86b4f561d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe262629330231ce73dcfdcc97d9681c3cd8bed897587b2a507b184704a31456e59ab0afa2dd7acf99542cd491336e697c27ec8b502c62d1dbe3cc9582513e83020863c733b3fb09aeb1e0ef18d39dd78122b4e2f3de5e2f9d3574e4cb4a531bf42a777bf175e32aa9d54906055a79248;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a00d2185c346dd6c8c240f285dc21fcf3a40686233eaaaa771d5b618f37d6098e08ce318abec324ee5ff1765cdd5182b9fadcb91cd35f193045f874d151e1e5b3e8aef9a0d506ce2166fae6980a49184bfad5702c74e911c28b9c803018eb4d2d005853df26d0debb99c88f218e50748;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcab41723cc5fcd74439442192452980a8823d304aaab85a7df1989ed4a968100c8acf92c45c3a0246dab4a36c59484fc15b8cda3296c57c8964de8ee90fa9a13f889f70e9f595b2389acbf477a1f4db3c107e64e3ac427bc1eecd67ae2ae7a7c2051aa3ffca55fb1d677185a737d01f95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d0c4efa5ad29fe5a06ace9dd96806733a55042dd299fe1e7d22610961ff17464220c6f5d9c32b816d857b0a356df11cea0c9c7c6cca4bef3b276c83670fe9ddea4d8b777dc6c09d95209e5ca4090b712def7300abbe8629dc80f4f709f40f3c80271e49026920748f5a13514c55ba6ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae065c4f7dee85b6be1c5be172f7061db8049010dafc586cadaaf807a07c05f78b1583fde43a9fc7f3735b1a0467ae94cb51f46cad8cecff5a7b130b9490e2909347bc1e4f624d976d2b4acc3d9089dfea2d6e0d1a4ba05653c2589c89b5f4603d0118d54432501a354f28c6bb51eefe4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ee93a7b4ae574b41b215c47e3f35c87cd7abd2b6a28730d89860ad874cb3a7b574538e56766e207748d4a7da8b38e2ce70a27230c4404d7b978c884148c94c028c40c967882f932ad7330f15d3e96158c338a4068ef2aed797e44c3b05212245feaaefd3790bbae2259068564102b8da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h196a49f015f07307d43026a25715f506fb48974be6b7c7d969fd79d352bf29eded59152ea1748826f3df3b25e2197b20904823dcfb9463b9a8e4643928367773ba8c381b4b28d836c9e57b268ba4345a3bf1049790dd04d60ca0d0f704d414515a1efdd9a47e36aa80b4275bf217a5ba7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86d3256eff2374fd10126a7b86396dd0072c6c744a7fd722376984d805da7bcdaf86c7ecd3992ce0c96f7385db8800af68836d1d0f5bba5b198757d83372b0be12dfd97b9cb429bb4430e272c39badc05e5757125632f1752d09d5202ea7ba43de68faf8b36d1cefd3e6a33e5dfdc655e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1edbff9908ff33c6430a7c2be6d0593bc2006e13687b2939a3b3ce5d6da0c9a4ef3de77068e0561159b3306300d30eb8cde09cf308a610f41be27934bcccd3247fe93c49b577a1366585700104b6aefb36c6916e5a7c279a8f8af39e5fa66d61b003dea5507e99c737f2c2919df77720f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c852649aa5a48f723434ec7716f4326673abadb97156a8edb10cbba767243b48c2368eaffe1101f2ffe0236f5f46e60b2b216002791602906a67bb2aca62ba80bfbc01c0f4b575499333a8fc16640434416d0dc51981810bac6a19e1494c6fe972439ad82ed221595ca023d9ac0f1c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6625d2880d77e4aa04925693374ab8600f96c34eb1a07e4fde5661e6b8d5a0285934175fa383ab3547589a84518a9d9a00591e1f287af234e8d3a247e41a242f365770d81fd7d6594a7884c73ed3fa7a5d71b1e66b3a899f0069992befa864ac90f1dcfc6e73210564021cda11a331543;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h627c9f82a6e95746960962ec707c041157db7cb3ba55ad13438a846f4c992fb10a1cf4e311cbd69717a6df00d0a92d1187d605702c033a190a8935c4da5961699251c900fb3e988dd433eee5852dc07610b670467e3da137d99de81e0b0db53292a1c0a898a558c68b675ac2b90638453;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c30a7339fbb1568dec938a42dcb2a29ae9b68f3dcd551d4ee574a7896d70e1bab258e19449b4afd480c34aab56b8fea3836e9fa83f0b4006822ab941edc877360331f8b8a503182ce5314b2c02b8bf5cd1dba95823b1b15bad903127656e96957225f562c01f9f6a2c891ac354f03b42;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a1e22f06359ab23a1fcdb8b8ed24a7a2c7b8c31fe73dab13d6b1fc2c7c7b9bdab08b25382351cf047583e5ecc44bf7ca7b87161b03a20a013d5dc339f3080edfdab01fd9f49f67533e2dc9b70c66b0858577cc57a43672eb88f29e6255988b4cec4ce85c2f018971f9ab30b56dc417c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9f97b40d94207efa18ef2fd22abeb628efec4634c6cbde096ad9a8e8b029e82c0796ee30e1a3832bce90e3df40764a9eb3b6e3b12168a209ed17fd0793f47499409df433cd99eda0eda93050807e28d649ea268f743130eff2172ce4e6a05d64bceeb2cbfc2a8727260d7cb6e0a694c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28230532b7667c04527117855288c66868e4dbdc3e0244f7e90d79263cd9bcfd82b9a501d86a31af78174980f7704355a4411b14efc7d48f48af64449e3b9aa9eefe73bd88399e28b03cc14e5e41bb5422efa9acca6eee67fae0477dda46b61f5dc57d9171df14842b1968b8dde72d364;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51760aa0ae5355a49c3bc1b7084b07bcf3f7fd81f298599d097da32ec6fa0cf84b1afbf08ddc0ec256a5d6ab1086073ddd078920e93ba514f5f8f6761be40949f85dfb56c23ba0a1c6f01391f1408a1da137cc8e04d2a080588fb4f618fe3af8213f5aae3781aa021048b145a98a9c089;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6c874c6a5abeb2a2969426ac6d4401d18890da5c4f21239ca7ad7006fdfdd224b29c045cafce38e4a4b20f240975f72649152f848f762e62127b41ae94742af94c40978cc4c9b5d741ca8a89af3233cf25fe5c9677a011174725e83a47c4fc4fb2b46fe2fc209386463a852f25d59b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f60db0b240797b42a1683ce4f43cc28d37f73ac42131cab9a218a2c5012f83f4309c878afc00d1c9ed2e584cca46c8255cd287ba5913f4d38390479c5942d3c42d3b62ab5172218ac3c328726d6f7a65bc4f4e2a1e73c539634c792ef3d77f837635f7d5dc42470d9605f5e464fcadc4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbfaaf9428a8a510657a7a948522506f3366a4440cb8086001c5ae53995fe1b13b31476355aff785ec1a27cedb5a230814486a8f927c265fc3bc50ae21cd0a21be9d74b61ad1315631e5107db117c0bd3c04a2392f773e1e1f61f7499109f08139248f78c6af9b85adbce0a6fde22f517;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h305fe4d6add3c7eae97a06263b12bcfc833fbd917b59f972742d0b2e5600bdeb9320ca0166cb7314c4854a16b94f8b5f58749686f6b466a3e404a69f594685bcadb50af51e27ed7ba8b38045ec8ab03b44ec038e1aa7df1e274836654134f5b4333cc9663c386d8565a4a9f8b25c75016;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae3ad09889592d24b2719b975831878eadefe289f057ddab3258fe4f5175d06d8ee2f94687bc32e74c6d2a5a5ee34c0b567e4a9991cd98637d8f438e09c2e7e8734466231197f49fe4794cc0c8c1f0bc3c992819e86ae640c918b2fcbb87d9110176dd03d1003333cd384ad26af592ce3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5e1b40dd73baab8169dec5f9a3b60e6c3f18296371fc73134332de3a47a01231a8b9f44d100032c7d540f66cc7643d7e0c6715124833b426e2403f8becb404bf469147895c6da81e8800be94e36cbe97413f0a2e4b6b9ab0419f13b1669049dc293d4c37152e2998b6262763446d5ac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h116ad81c5ce83532204a0e1bef9f40e4b5b6c9992ebd8d6ace90a1abec8e3d91646beaf966c8086b9f48d0e2a591d0067e7bf4353872aca21a7a882a8961b081e8b48285cc87d91f6d4f5a01126b2855a92542257e458ec132b088f9db93b50249f95d0bdd17fbb01588f7ca98af38797;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc37a08102a00b7d98ec596ec8b7746f434b3bff0a8b507c60a7805a3da701df1e38cd8a34a34230bca9a598e7912b6daab16e3a7baebe0732af218ea899d107f69ee21fb0ab2ac9aca613778b4c45e53f01bf45c529cbc12bb15b731d8548dd785ae81c0b1015f2accc112197a0d2e219;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d39a47bcb43d75b52e9c5b47fa9fbfa94266d237d8fe2e7df5912b252b024990aac3a6da33738aaa70c1e36bcf7716373f4fac77f3c5ac28f6961e98bd1f1d71ba944ab9ba23d58bf6f8c0ba9c2cba370b96081b671bf26b1ef841430c0b2cde7d7ae854139d56cd0313195be3dfbca2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he85645765dfe115bbd08fa6a49f2adce9fe672e7ed55591e954a89c6ccb665a5c4e78e9f76192dcd2d9eb5cabc02c5e980bbdf00a34601aebddca250c7f6507184bd059f6e0c6392c89d1e938b1007bf0c4e03c3cbe1b3bd237ca3b794609601d464bfeabb7fdde591e9e49dafb1c78cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb1068e7cdd47085454e9c9765ec0594830d55d9c8b0ed5683aadd436ed397873977e7f1362b92e0bff5e84dfc2841607588567a7c7ec4f224e4382cb16f13d08ce0ef34d573b29e39999cc779ba24595fd9e58ecb4687035accddcf86a66e57d9076f270bb1e18bd78609f9cf50b559;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5bd2e52eb240e71f78ca8639edec3643ed4dfa572441d9e919aa5e158dc760caaf8e24375c8eb8866ea9407cad9b252e0f54043b8c024a4551899812ba42b12199ecbca5dba8c6ee897bc41069596c850fb7442b55d58471215a5829c6dddd84847ca1e798e4238db67ce7645f146be0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5709c36dd554ef48cf2bc771ec467380c49775ea4d7ede717c4c1f1f3510a58bc1609d14a111fde3b2811d98ec0d862a6305cc42e7abbbe31bbf98fa7afbd941f1c7068fd618427057a6f8883ba81f7a5f2ea8d6c061c69c08ac8c1a8a9d7edfef957317cfa4b3b2e409acf42fb6a366a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaf67755ac94765b2096356b9b8ae8cfb3e41e211a1c4e0763bc42e8b30ada2949a31c340142688b3468dc3b37bb5249e84da3fb9ac0426fbe8b3bb0f6302bec0eb5c7dc3e1f17c9250d64984c6387d77bc0da86e4036fa46cec15bd65982de5daef8be7c47d13209ff9310b211131d0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83348321fc10c2256521f47ecce00c19d1ac0332a9f2d187bea079218a8c96b036d5f63125295efded6cbfa8b3f8bf929817b8510c0bd69cdc55947da28803b624afaea6ae5ea442df88cd038653ac51b0d3a30e83211159f5eae82d2ce417b4b12ed04a90271ceb0dc479bdeb0dfdb2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1da30c68a4ab20ff63b4ae3ed440363a4b442c31c15652af9afe39db1c2befd33d101131ed816d99c30ea74083ccc4a2ec8582c2ed1840ca72d9be33406ce980d813be8e01edeb8eb8b2a933efa83bf145c1cb52cbc47eef9ccffaa9db0257577306f0859fa70e990fa740871159244f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4f2a16f0843f59441c210f562c252264f512000d395945359b4d4f5aecc9d0ea27fcb793e91a499072e72e6eafc27d26836bdf68835bfe5d19e9b638045c8bee16d687110c29b0834299463c23e8e11781258bf3df4109afaad52a654854ccb03ce166981b0d514a4fcac4ce12cc2dde;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac7b90dbb1493b24278c4066977e899f0bc73c4f3a53ad563897afb7ed73517a3aab9c8ccfbc590e67e3f232f1f5766831afb56067a5b3d3400075f7c83b893bb432e4e5d820595f0c3941dc99ffecde1f276ddc5f58f60c58d0f531ae4940968965a2068cf0dc8efa8cb10511325395a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fa857d3713352267e49aa4bcb6446e880b72444646421f86954b0732d2684998cc51f9b7707c73fa35e212b22329fd69f01bb2723561e252b5016db224f32552842b7620fcf552f0f0c27083e91c48b10a3fcc93315234ea1cea4f6fe70d47e56fa15d2ff479af9064eee6e058616353;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb1d5f6822c0e9890d4677916e78fd4b13a8dab2a77af4b49746c0709d582dd1a2222045ad96af0b5df125f863fd60d9f222259747fae6aec26aa47e4b396bf38847591095951d14efc7caa2b8b60d90759e555a8a9f3e0d4725660f9d97f01f09df7e5ad96d29726a12c5a2cc7bbc260;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc064eb53071a5b26bb4e698f4ebdaaf1ad4e6ef623398a64233ac3ab80e183e09ec3e593a3db1f432339054e1f637f73d9b142347b6b0894eb3ff80d9dbc836974e0d48baea58b6f3a26557deae2c2cb46cb421c66d07d805dd9ff35f821f8c41026a14cb63d3951c01c51a403646233e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f28dcefa6698bff522adaa46cec6b1aaadf6fba9654433dff0e9120deb31374b40c275d885cbd5c2a05ad2dceb3fad30f2e25da9a2634113b8f445426e67ff9ecc7887423ddddb8cdb86e071d390585850a3420a99acf8dc639867c510cef95c2db6da645ed8a7079bb79058e01c0248;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8a8acfbbe0dab6e9812e41dbb60ab130cf8e023fcb0df6cbdab2e048d112c2d3395fe0fcfe6854f167ce27d376b82eb5355ae5324cff9fae3c01ff4f2e5a96f6e88b8c3cfb2f987ce3f6a348569a15d643082243f0426af4ffce015044637762c13de222fe563a66f94ec7cf571df99d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h931b1f8af9909ee6b99d4691e893e6aec01f581852ca320d0a61b5024f1690af125112f007f3885ad51cbf9f266fd797ebe730e761f4d61b6b96f17e3ee61ae626b711180e1871431b1f4f4beae4f462b093748c6829c54f0edf28815db80ff3ca52e200538264e3d506eeea46bc6732f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h129b118deca7e0954b784069c5276dd506c57bdf1a51c6c6b23a51bdc88d01763737d40fc16c896c755415568360a12e1b022eb2933f5586cacfa0c4c792b00b9a4bc775e99c4feac2ed344bd4bed142c23cc96e26022b4ffe3f3bbd55634dcf27a2fb31f004b800b50b56c3a794f2d83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6e5472dcdef2e9546be9b3081dd7b22dd2136b81437981684a757d0219fe00983c725dbac438ebbbfd4f71f732f586e12f2de37cd8c1cc727c959017c949edc6ef2890ac2553dd8f9ef16695289e0e58ecc4f77764dec8d37f24f490e1ddad6ba4d2c518e839482f1ee2afc1f40919fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9beb06787c85e7fc5b12b49f538b07c54ebccff195fbfbedce4633a519bf36c5cb7ba4c4014a8655303e17bb633eaccdb40d1da14488f1c0c69a92366aaf0bfc9578951eb2c4fa67f7ac6114334ebf58e342457c60e97fd341233aa6f6d2834fe4346a4efa413dadd799e7c7bde3d847a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5b14bcabd512bbab4fe800bfa24c1db3f94d5346edcbea74c11125f7c60741d56531d69bc4f74233157fcb79d1d1d78764e2e2a8337d064852f489dafa490e946fb4d1f5dc02db58884d2785181d880519fa68c67c99ac7d894f483c6b45d94f88bea322705c70036a57a7d4f605554c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fa2aa3a53ea12e4290fe250e56b2e73f95a4ff0d0c5e3c13f3babe78b4e471f28c285eaf1866c6ef7ad152014a1bea37301fca87b59fc9fb4cc67024262830310502914779f7174aa3ca39787a684fee23343ca720f5bd28d91ced54251e8061f2efdca9f66793115a49fdab17d185c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27ac98e5b83e95a946eefc3a44a45f4b1b4547e0ac6d1d16ac217202e36a43c44e51f5fe7d1ac826129cd8734ef21128ecab5412101f633f4873f2c66d59aff01ae0f899a02f7d6499b56e4d9b97eb5a37a51b0aa6be7b47d897487292912d464e39c134e2e42c9f09cc77aa7afcfeca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h239e38d65d414b0c2a842d9f29d776da1922b2b4d2af388fd3c43a11e770c169b9efc35a981844a2a78b41a43c6ac59d1bf4f8a3d15ba87b70cb2d062f1c7e3557cac92446479c8c3ce537ccf84a9bb808aaf10260f0e95a29c6cb542fd3fd7485010f4b4d366f04d475d109dc0725500;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75a58e7427face5ccee793cbece0c64dc06b0ccc8e33ced35d76d81abaf3c5d14b904e84f49eb261b006622d104f8094bcbab70993ff74ceb94ac9547bbb48c5c380941adbbb5566ef539606227922a975baff03dd52e8e23c77e70dc7b4a7a12914c39e1795bef385b09f99ff7e71850;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b9dc218407e3f821f9d7fb0342b3c14acc03638d57c8c8a209939d74969d7bf62015e007320298d40f24326a8ed1325e45c0c7ba8bf126e8359856f92c6b0fc6ff6f8657073d18d060031cd2a8ee943e20ccf510556b44b5f650252c355b39ae57133858278e6768ac031308d3718427;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb303ddaea9de9e124b9f453f3b6b008e44177ac3f5fe1b46a306d9d7dbc487622ec9173d82781d19d7ff34939256cdbe5c873ffbd8e0550ab1a6b711e0cd5b2740e6b5d1b3c40b706e03b09f06b6a6c4ab336d1c74910c36c7adc73f24c1e720fce78b8b3720fad6c30968575a8f2c7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6323eb24477b3b439bdb9548f5fd85b07a2d8defabeb10a204dc63b62cb842781262e0995f2103dfbaa09fd3a615bc6dbfd9159da648f8c0d210f3b4479ccbe56ba73d5150ee0aabe98da18ca9fdf0907de9507f5d120d0de4689d20b01ee3504636a78883dabe14d84b36223a5464dda;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda9079c8c56177da64d461166cebe52c6c9b1f271b91953f420b99c40907c3aaa16dad11e3b9a8712e988f737ed877a6071582d1f8c83f7ee6f78d6953e96fe9407a82630c36ddb6a4230429f62427cc9762e96cbc97b5b61043ccddd03d1a459ed9149f6b9335a074cb732fa98167d3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb493cd50afa5c58c35b3cb8475e872db183d440d6efe310d5a209b95a3682704b1f162950349fa4273611881a9ce17e897701f76d114a2002f611280fc5d6d4f04254459f57617d0af5f5d672116525b9923ef6fb059522a8f803408745213a010c313b9ca8cad2025f1c56513509b4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99c54cdf79a1c8e1a6b699b35eb6d2be0cce3209fddd1d23139f28006f439e98ace0fe3893457075f8b1a8080dd10ec4d33c5ef95b7f3bf48b65ca5c551a3615f4d3579fbd053d1ac22df45d59a62921c5120c91ced183e4c686821a4c63a71b0e34656381087888432ccd5bc0b9afc9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ed86659f98c252d5625748b71a734faa35eb21f2870da137276f3940af042c3fa9d3fc70244b5b694844fa190e2614e719340bc09b8507b81d8e0830fb40ae11db325dda34b258c618303edbab2c7f71e524ff069aab714d8845ca6a24dba2fa5b2204f2fba8222176ccdc8f20f3d23a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31925450adf692d0ddf1e4754e1e39bf0f90e4987e4d41e04f76588f2bc166cea7cfa4af0906ca3c5a1f3c943256d1090ce96122084e32f4a60820c9f3d8a3a9aeda16aedcdf40b0ebc74c495ab97b4375aefaa5c785c506ab48179b4513bea1b2a05033d305388c437a77be8583d4b69;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h956bf0e3d6db8d18b3922a7ca2410fac6aeceaa0cabfa30dea8eaa30fd5a50efd09a1f12cb2881a00753ab4b5b2151a74de70a712e969e9db7a5413b9dcd06bd29ffa8cff4b4f59272079158425e6cd82435118f03c4c3f4b6a2d0e61e8bc7be9450ac84380d7b3df0d83dfc3aa12f28e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee3165a14f5efac3c18d34d351294ee9bf59c3b603b0d2e6b9e70c0c8c13fa450e2fffb62c3d1e00d9bc2b69039c3e831a74995c99788be9c91c28e73d5ff5cfd87cf7c0aa9733bc97b5e76b57d780d6bdb04c87da82bf74d874d00666c47fbdf8cd4c2686ae13c076e7a5c4d760ef6a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h513d7de6f9928599711975ed71c6e430e0e92c4b91bab1c3a63dcb6b91ca5627aa95552970b4ae330bc1754d7014fa59e562203a411f45ac325d9e109b3e4ef5c8e0b1a7651e817b865420bad2d102632b619f37b2db82207e178cfd844df3d6047899eab35efa49e6a2b715c76eff55f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72c29bff0afd3184a5f1c09493cfcbb160f9e33d6788bbfb6f40f61d871402d27687e807cbd1e923bd45e9c128b99371482e1fcb6e692319b87071dc8aec2d86213292921b873af249ba46d70fa1c1e305a7ac473099e9e87e997dd2cdce148ef05b6d8bfa1b639419724ed623d902917;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc6cbc5b92108e2fa2e286aad9001e9098a7506d87e5c1e2c163e23832ecc07ecf305961efab6e651734f4edd51022c0449d4b178b2650df5fa60cf4632b5d85f349040001bf2c98554cb2206d2788b1b0ce41f6b1307396d52a28b9a25966d2eef40dcf02f180be3cbec0f358dc397b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfedce1d5cda7867742bf0327235b3125ea3ba5ae0f5a70792b74184b1f496197cd89e0e70d6ec68f2f599436e7ef57df472841a357b5f38b7f38070b439a628cb80b6c88ee1087b42a2cb7028f8155568ea249bccc65bdbe05301978142bebdb9a0bfce2629232739238562074297a2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51c984c3ac353d69f94880bf5c949ef2d6c7f5d7ba4dc352055d5512170ec75d0b63142e8a39305d5b3053b78162fdfed7a887f6799386f7e2f70632c51a58b82ad503c4c01ccfab67f2e47e12b52cb6896527ff15423e5d0e873fd9d7dca9a009c70789b5f5520a3eee144dacbd91172;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae082afc6b1b638f2e22358b4e8021d5e5494144a8140d59e652cb1a01ace8c79809c4aa0f9b3be88af526a0884f561532ec7eed3a34884bc0f2cb17717654eeb252e25fef322ffbfd999b12cb311471c05ddb4403c6002f4f6037db106d2f72498f184912d7d7049283386874b82721;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecd59a71f222785c5e33da04304ed32c2e1b498b4b6677d9d82f4e4ed4312936e1f169d590f10ce972804b26201ead3e022de4cfaa82d7e23d982aa7d338c45b3ff1e30a4c6504246b92fc23e87c8220f59b22f88561dff5d65954c99841383c9c2d318a8fe34707e2af3083c5cf0c9dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bef10e7c2bfb7f5f2267e2c8165e88a4aebcccabcc5ae3190ff143be6e9719b289f275713f97310331b062ac281d7af96eedc21da516a4b528826718a6b626b3345c2ee87b0f7391a8bced550b086ffd4b9c9ef975421354e9277eb380c067c0991281c65f4712b3cdd60acd584389c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf97d7f2afff2db16dab183c4a21fd46049152f655a7c71bc5c5ae1c95b7857df863efc401df8d9942c3d840498e9bc168e0cb0642bf3aa3f000ab13e1703e413ab7fc0907fcbb4053bf491bb4d49c66bb2a0b2386b3155d87d496e965860daeeb8ecc7a577a0559cdb093a8d886d990fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90c3f28aedf66dc030739286dd17b1fe124c15c788790cfa000cbd2c00530a15c87c800530d964ee9a6678477b2c74d0af67505aef0f8663fb3a9b3febc9d5d7dc939d3a81a8bec8cc8c960db63d977ea25cc6789115006083071628a6eb69b6c2356e66399d088d1decebbc1f13ed569;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ee2b363fc73951ca4662e4d2ba8be11db0db97da91859494ace70ac11d3ee6af2dbb8c129345a8dfc4e9c4f30768b3e64e20346a5ee35aa6e7c6ac01b40a3a340cb813202ac254f8cc14900ec46e41226f6fb9954434b00ac8c27294ae30af83e8a78f05e415907c2ce05e35659dc956;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4cf274b633a881a3a42bcb033967dd0a9f2a36d4cdc309d5be354c7b8a0cdd35cd75c54ce444ef1cbcaeec53e850563c735c7384e7449122db3e1e58d6b9e44b11431ec26f8d75fd4466cc6afa97688bad38124fea23978373ba351cbc9346920c81f1fb4d1032ed952229c61c36e3b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c212aeee39269163fd6a5f32e24b9a96d362e5b1b4f1139dd0a57772c61f227f98fab1ccee5d8e71657ecdc5eefe2432141db3cc2f0cc4e0d9b788e645243e8dc1876e0d819ac97530f3fd359580e039f14a11be20d735e9db4dda806df6b2ed10dbb7903f6776618f15e445fdd774be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81a807b59b369f7c1cf560a175baf54e716351342c20d542331c0d6a880445b734521024babf30b26dfbc2c70542c67bbd4047d1c2cdbc971bef2594dac5823f4270fdfe0091ae48c5c7cb73ff6e5615ce047ac278accb7c121ac6c3da7981a03c5a778faf4aa4becacbec2416340c63c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h364b61245c7b095fceb817491329785411a438ff16a542caf97556b70596c49886f8766f37bcea1902d8dfd4e34919e4077670415e3cbe3e338cc659800ddb15d62fbc6e23858b7fc3b42539b7dda53e5aef6e08f2bbcadae5902ef4e7496166452b473c0db29915949e146cb5ee17b38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64fc754f94d1fb9c86d75339c116d5ca8db32b3380cafc94b249f3a8ba2410b7806362e3652b38f297f8be6a2dcaedd284b3eac2bc2354c09900e7b86fd3ef932bb7468bef4d53410dea508e3570a61234e45642487d65e1fa43f123c984e25a0c5d197bac16c729e831ba2f14bc1bdd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h544f4ee89a5990b7f06eeb7ee47f63bf1be9b9a9ef5394b099e6889b5e1ed559aa87b4c22a41aaab0427a0be8718cfe9525b616e0e05fc354252d643caee7a6968c5744f35ff982610fbce72a75954c8c585460163832731a68c02e2279db28a89a76317b2b3dad50c0e4957c336a160c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb351d0ebaa3db29508b0ee9cf31bf6ad5ac2822b366b534a9b738fba161797f53acca63e0c67054931ec79bf3836405967b25836837c8484c65ac9525106aa73160c098b2fb65b49f5f4718cbf59fd13547ef9b61d14046f7083f697eb62674026ab2c81f736b538f1bb385229d460e3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h924b8ae5f336c83d1cc121012913aba5cf355a4b8b5ff4161b7732a82e76261bfc85a98903b19947e011d11b352c1cdb04a2dd697df075f3e1152304eeefd0ba81b93654dc6c37620c0d8b2c1df28f14e2477b1e334640a25b984c66afeae2f2fa61fc9d0e961458ed28036fd90aabff4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ffa91bde456f8908efb26152302db3b8e9ee30f556176560691ce1766111786703c11f9b34fe2201d83fbbee4a19bb6a2cb6aec877d8e307a32542d451c4bf63759e42e7ebac1ce63c012522853ff36f32d2fb70ca1bb41df18dd8df80d171620843064d7d91731818d5cfbebdbe2f83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f36336214bc73f4f5dec7d8d60ac7f35bb95825770e0be25b048356202748cb8cbe9ce586dca97b54f6039ea2ecd843742f58e510109e889209458e4fde6de6bf3a39cf1453be3857892f59207fb28a5ccdac252388ecaa4b33f454cd5a8b9e14d7350dc0c2411fb8f0b5399732e3bbf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb33e1f11cf87e55dfbdfe02237d6587f0bb1bd331c3ff6811dabfe56d82851e6d7c9af6759c34e206c0f2ec77fbab96d8adc171d2774dc8763bb4243ef98d7ca7e7dbec35f6689091471e3088fa1e6e9ac3fe7c8b1db37e53aa7f90cfd7380408b18865e0345af9d1766b5200d50d70ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2970f2e55fff333734279bd2c539cff77e2272d50ba07cccb4d634b9e04b57a00b5084ab1e30074f9d6f57c64e83444b6ddbe4eec2cdc97b7df1146dd868d7e8bcd396558875cd2a0433cfea58c80424947974cdce618decaae829fa17072f1b28f7de8da50e0445c6879956b5aa3768b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76fcbb5ca7d10392ed4a194c57c8418b1dff7c5b5eceeca489cccf821a63423e6cc7f122786fb7827954687c7b4dba54bd0f8098a1231a4044fb49bdb434fe6f56ca9d0b6450773ef12ef0fb1efa5fee72293eadcb1e0c7858e34f0ce49e91ad43ccce938c5e95b36ef5b5cdf6dd4f33c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb82f177fb121959416819c4da779df51d2626758d0a87efca527505b7f63f1f47ceea0399efe9afafd4d52fdda9c3acf1fb6c15f2ba660858aae7786d38e6a547c4d657da87b8dc12256d87b7fa525ce6edfce634f52c633134c896d27b71fdb2e61f8f6e3853a580b6f356270396dfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79f149db8bd0b2e79b00bd92d70f5bbeb0501ae62fe403881ab72eaf6cefa9356d7c43e5fbbcd15265ded92ee1a9d9fb079afe1182ade25e36d622174031cfeeba97908e16678d935939a18600a62e9261434153c3348d6e1e72caf8df963ec3afa85bba5e1b1f8133bbd29b21787b0ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6ac94e58f76bed931a385c47adc885c1158aee1ab593caab84a1ae86a646e4073722a102272b0586cf7b749c5e7cb8a6e9f62146d91173f4a1c8f315954e4369d9865fbe3dbe74dc9aef4604b5fb311d9f42008eb92563d48663f31c5a608f65f57e213185d2adb05de1cdeca047d44a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h239ff872ae00e3186595123cdfffd672d3a6999f0eb1ba6b1853dd1d849806b9522e10c22223b56fe9b6c1d049ed556b121e8fb3b289009c5aec5e2acc3d5a488e3c077eee2eb150ab556d1a47ef9ed3a72e4a1e9b4bfd20bc19a4ee53776713c2c51c775a425c641a43e1bf23951aac8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ef22f6eb002013517062a8f4e757a868527aed9cfed2aa1ec56d13ef7c3137f48cc2b6487e1d64ce1c73d8757f5cc5b2129f5edd68a69d491bd50d19481351393a654362bdd65958c2c1cb470b8aebfcefaaf194f93ccb4313b4b92c1c11bd1e59308f87c497ba7239d4101fe115ddd5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5788f9b8172de6080b50b090a6190561231bd5caaa77d48110d2027fa85ae1821203a87f5538b6c5627822fef675876c80c9897146d30f93c769deb0ebc5d7e01811f46886b8a348a4df730d2f3c4d3a149425b9c66043fe9db84258d03e9092e21dd97348ab5f1c42a13a9beb6204311;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18c6afbd7e19fad5a817dea83a64bc7449a19218140f465f8605247e4926a51e6be5983939512b119669a12298f3c1c6a0d9c614a9ed6543e8ff5b5ab2112153ad8e09a53fc106cfd54b675724358267750a43abcf0d9af2e8227b31c3f1f792eaa905259742426b06554136f988e7bdb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6cf6ee8f2f9f27486ce22d7676b68e54f58ba10e6ae8c83d16b5d37dd3b84b2817056cbf32a189ac38a629421ea2052fa3c7320a17e808daf588f93e74ed51b5bcf9381ba8c5745e0b5b2e973f3a51002961151555ae992b5e39443b84e6d0031509e2361ac64c2f787af52f9929f267;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h757d2f517c1b5e57ffa8a601f55ad50496aeb6c929b117c900378ebb42864ec3f857cb7ca3d243df863865a57bf6f6aee5da10a40801496ec77f39321f788f140d2c1b643c651d376c508c1a61a1c160b2486becdec47705d730c6c16b5da810e74ea272c08408afbed088167b44cbdd0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3ad13fb2341827f3e16357b764f83db5e3eec2bb3d828100980c31074cdb89bbefb37a5a807b49f88a87f9837370766f689d48fe781166f58d47e2aa0f6a25a43adfa0f0a75e7b3880ede2b214126ac1d1c6bcddc1de5e4cf6a8a13acf99063d822c2076551694d67c6ff28534a06a1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18c7859dfd2980c98861a45c81f0f95b74dfb77aec55d46d264c3007b7df8e412c7e25a793786ba2c5a2a27d60fbf0eb70d8d16a379c9da870ddeb0090d8ad3218972bf0d6618ecc359befb1f31177e6d0c986da3e2ca14161d2a33aa4e438591f9956c86577c845b06d8a46f4abed66e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h826fe3210cbbfa359ef46fa2855c45861969438b940531cf11605cbff3003ee64da26e08da1ab643a1b95ffb4f13845ef664fde80d29ace5c2440ef21b3f2bee9b032708b177696958e04ae8d1882ece4a6ddf6287dd4fe8e7773671d1ac6d3747b278dfca35b1f1650ce704c28aa6090;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc8cb93c55098bde080a6275745660fe5716ca6ec6e26c30d5039f69e69a91f1db9394a6b7ed1c6a39cdaadafdbfc603fe01595a38ee7689a6e7d786f9411d66220faf83def842431ea5a508389afa77e91e77336d2d215384e5684a9849e094cf72be27867afd1fd3c0c14199ed04691;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65ff9a8583671d1e70dc72a8875658390ccc649645d6babc25a7ae9e373c5207aeb91241a94cce2d76cb598df9b60bb465a14e474a20b11ff97feb221ed2a750ec488fae8108893c6eac111b7d8393c5228551b31ad095d833f9a63cf89f20178d57dd62dac1fa20c7d3141e79f0255b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4d4ddcd02594216c4e79faeaae7413445e275b5846f6a4927fe3182de68610070229bbbbbeb461acc4057fc8eb0d3ce01f031ac7a4c554bfbb86fb0cd700bc997bf043adfc071f7125f12d05fc65502176660b78d88a0d8c96e4bf4637700cf0a718bea831a6ed3edaa7aa52106e89bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3c94e3fba36691a5b0bfa9876234f3ddbd7aa23a94e6c8de7fa79049e604e43784667c7896e198c710140917a4d4afb693b9c262234b95d8e2e2d7a3db0cc6fd8e781ce3c3e8585b70350a55bdab884036361b52d30b6b32c2986bb9457c5413f41e198ef1e4a8755b47578183f90744;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3cb8a34894031b0c9071af1ad19af9da804bad177d395b01a582f3f7af811d33d862839c63ce2be5f600603cb42f8a7496cb63986a57dbddbbaf94e9c3b63a7249ede8fa12a180e491402ae603a98621df2f80a15f474cff2aa003871280a05193cf993a8642c1401ee2e5a433679d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd19bcd3d728fd5d70927a34a3cda2a82db2d49f28e4fa91421baf5603417e1b91f0c66e039c69dc806243a37286844919affadb346ae424dd8df673bd056c8788a848a1a1265f4a06c964beb61b38081e3be577e609f5b8fccd62e08ec3f942f902ee9d941ec120a77614059074243719;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21b4c6356c43150c6c1889ea27b70dad3e1ab0979f1e5b1c2bba91f54fa6d493e8ee25054c48684fd668f29eab3b8deee8622d796671333b6372b7e12616e979a7213eaf91b815de291fa77f9c0e354e4392fad359541591734c28c463419ae5a405ca34c7bce353719c250fe1c9ca445;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d041aa6173e90c735f259fedab883d647e60ca53dfc91d2e08cd7f6cb7b9b43390ef25efdba504e2f2a1d63416ca4d55a908d0f85efcc6f1c16d65a55b71baff4db4b14e686ab425b214d937e9216ec30cbd7ae4b8ac712a796254e4205a4ba95f7bcf0052ba1c7abf56159d589335c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaa9f41f867198ea7437935a4ec95443993dcc32095614acd4afda4176c209af3bebc573c5ad58cb68f591e20063c2b16eae826452aaa630d7f8f3515a9726de84df4f190bb7d702683154fdce7eed7f4620e8aa645631c06e562d0e50018c19855c7c95c653a3e2d255f9c1b6e4b0663;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c7e23783969e5cdfb0ac909a425fe3683a9e220fdf458df576ff004a24c1d32ea21449c0ab0ee374cec6bec56d6f2fd1ab1a552a43e1b72b6c336900a201eaed8c14fb283670c1f44e8bbf0dd6e01c2695f7d9f3f48bfe9fe4cff95d882b57ad1cf0f149b794cfb6cddac4bee20daee8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd136373d6ab5145c340c8a8ead8b1b6eb7399ba8a0b069c8f6c04da6dc191ef5611dc9937971185e5f06c5823b296e545e4f1d514104366fd4ed374ba9897e5c0a58605203ac078b4ca333b62bd6c58230ef264f0f0d4d5cc53f4774af6cef125613ec574cfe7a730040229a34c779;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1114988905d3ff0baeaa1d1734249b0c8a589871a83609d57773fcd7c16e6577a47a47caa8ca06d62ccfc5f427df3a1cc59232a8f59452c522b2104d1398428ec97ba6a8e363f7f4eace1eac860f4dcb7a7ff6c5c116d0e75ed285aa03e6497a7e2336f37bdaea3cba3d8ca079c23359d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4921507dc34fe5dccb39f71f217e98c2e9b12884aef4d98931890323d192fc0c32ca5a8fa85d14afc03acc42f318beaff7e30b1cd0277410cb2e1cbaab7df8712c916de75db1f848ba74fc3291745349027db2f0cba5e55c9b2efe351b15005a22a125cf6e5604d441e48afe51182e823;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cde592e15faf8ba33340a48414e90f7873bdc047dffa29d0bd6178cdd5856c8f874529c96555e762768fb2c54df7f63a8b278602e4e66e41a0bbbdf1d139c7cf15b87a720ecb0bc82e670ed371ad04321be2221091386bd4556dea1eeb30e00260b75bef8908d7474396bd8d6f5bfdac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbad636a7727b6d79f93ea900322184683d94a12bdff40cfcb93d688d7d9396f15cf2a5385eaa71b50cccc16e0870b3eea11aa327de40d4ff88d4ca81e55bccf24459341ad18473f92dd12776f6cbb32b946e673888cd86af9b7eab79f05ae63901d3985a6d7deab8f5f72d62b9072d44c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f71b78498a63b9fdf7d65ac01eeb17cc8e30e4350dcf072bc31e1c8c5c16e6ad1de1e8b666e20d79540493e7859974320b61e6e527c5ed9870d1232d382add9403d858315f2be9c80cbded158e6f414ad0183847a2f430b1254a34f4f75abf215044284b35c8d949b62f57e27781a642;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41c224c97d29f205591f937cbd3fe7d7d205e31c89f8e1428fe89e22ebe48160ae31a0434e0cba1aad97f70fff2a9127f8fc24397d2ed9469bd4fe02e2b52513ee7ffdd8711e1d56ed0888c8796b8877c3123c89b8589db30b9e95ad881b878ee016983003289d52722e6b577cd524ead;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha72faeca5bd1e62d304cc04418c526b669a55bb00c9c5c3ae6410eaaaf5bd7451069e7e33580ff7fd31855d1dbab40b78a07d241a123329fff9691f15a8e9c6e46656867e06805b5d9f1836dcf2ac1714e31947ee64f81b739d3dbf27557af06777ab20e65b9a7835223fa89935d46aba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h976c19cbd693545c98d7527b205df42a234f8662f6f74ec3175477af516fc2acf5d3a18456dc1b1883701afb0ce7ea614d436f056864609d8f251feb08b695fa4aadff1e24c6f09bce66b1479fc1dc44f4eff4aba395f7aa85b283fee55eb3d4c4b6e5c8920f8ea48620ea716fb9b5864;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4a3c78cbcc181180c03c5136a78f72c868287f7675180330089ac46a981e6c94e80386995109ef93a77cbdcf58f4e386e873b046a43f0da5d1a846d20f5b8aead4b94b2340b76f55246df6a2974e18a4be28247ede93ff4197042241d8f8fc70223cd943ae0231f197b7baec7ed7e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8e883fe80baea6653b345933538922a53edf0f25fce5add8b48ce7a95394d17b4f2b81b701e3128994c727ac9e78f2ab57ebf2ecb10e867990659e35a9517b9e9ee0f3a92b8267b2159527f6a8464758169d2f4ffa0ab95cc3afea84a972dca646d7e40e842841033f9262ac5dc06b40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c5b2a072121dd201dcea4243015ca957e6cc99839fa3676a746afb10b730c777b796d5191025ea932d3d5bf8b9fbef30f3f2be05a717acd7418b22853a62949ea5e73ac321113e93000e60e31f5c2d53ff7cbc53477c4df29553afd43465aec2ca046cd65a4f8ee408cc07fa6d6d5d6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h770dbdf079b6e7dddf605b3a7acc7dac15b6cc2d65b2c9dfdf5d5bd77b0c21815e353bc5f5c4c4cdf7295691efbf9ab3df6935dda506bf7f06a3983ab1da7751987926131494d5007e4b4ce7ca590b525ce923fb765f02bbf1c998fd05dcfd31322b6b2ef98826d0d19b21366e7001300;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h119def8f65467f1ab6410f510b48a1a3526b450cdd6fbf67671ad7cb750809c58acbcf5c638a524a7fd912f953f0206342f9b9ce7438e93e2b984ee5f386ff3bf1b1fdf72798134a82e59e1612e12419e1888657d8b3dcabfc516a5acbff7319805282e0fb2457f39d9e82e37e50f657f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3870415b8bfdbadb5523064396967c719740fe2d604321f7518e4617c109864f5c6e902f962f6e1d19e8506bd6101270ba45676d207be4bba8d7cfc4c3fba2097d483bc9642fe508b8f94eb189386e84e5dec48509835d2947024b324ec5ab4b6c8bf1b0fd7d3eaadf58e3d101b6a42c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2214db9cd8261d78be4fb1d074532ddb3372a8d1540e70dda070e61648378916878c429a13dbae79d502cd76d68aadc7052473da193b3e6b2fca7295e3b9b7ee54de7cb0d282874321913f6dff03b62f112919a8cc720eea9cf600d47a7a6681fb89e9fd8970552841f7cbf895b0c4372;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbeeb08bc6b6c9c79a13b4b367bcacebaa2c950647031b7b9b552f64395af7dbd618cdac6820bf80c53c00801e33e74270c834ddd5ed95851abfee312227144cdbc2e5448adddb9cc28c1fa44e7b63f13a27be2f76fc5194c4f9cd6a2a81aa521221c594bdfedab58ef4a8f9e726b3e63a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1b2c2520f0caae2236fd1bd0620cdf898318616394216c63ed6aac0bebbe5ced687f7e30add3782e1c0cd5a1e84e8d435069776be382dc8e27d0c939c47f1220e76aaa5f263eb6026637a6697f12e02cc7b9dde889940dc47a3487a29dc051b9662c53a7bbb4fd13cc04305c84041abb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b1f3afea7dd0e53b0780893e9a4aeb3dadb17b0ff0a7575d08f9f356733d56d8b4fa2755cfe7164029edb133481b57dd07054f11e033663026b453ef69c61ca0c52602b3e2284891740d875ee368c8305d16546c4231177373a1d57e7df156fa4466a2ddf0a9916faa81e01d4fd96fc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9337b5c4629a16b8b81958f06a8ec9afd7f25913a95559969a55972c79848e0a2265f295b453b7ebe6cc97ebfe0296c13f6063478d159a3d1c31557c4d0cca4eab6dbfd25476fca726a09bb132919bfb07621824128aa75f2c1b9620b8c738bfe75dd110ebf4b0f6b805576f3e961cd65;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f881d33ab8dd483592c11cdc5ed8a7ad64231724187212e8ff6927a42d39cd9e70dd0944d4e02cf049c13383314c9acaced00a7cf24f4cea4e1f7ef68be6fe3b687c8ec613e0779e9dcb2d54d734bb985880451f021c2d9fdea35393abbc6b506d9d6d1579723d0eaddddc7972a8ff5c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h305318cc2f36e42c15105228efa27fbb46fd49f9b74e23a7bcd97012b371cd72ed299161a8a4a6c7e9a6451c9493bcf2e76cb1d683a315076285d948a7693f1808b591c2da1cf4946e3a8b9bd194a2063c960f90cc0ecdc4fe495fbb888fb8867ab43b42259dd7d8ed51289df5ed14d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55000de9f756682243c0be90280e9952bcc9855038fdf5939e50e4be8b86fb6cc4a8b79a6c231b4d970184de8ae4d8a5dfde5deb899fc50ca5e144ec078c1c0060256a753e19ae52f797e5fa09f37e3c0384a03bc8ed55343248a53205c6ddc477532951597bd924e370ec5eacc5e132e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a52a32a76151799dfe5abc4b5e525106edf217df6dd45720bef98e4f20593712214a47537cc70070b16183c912002accd84e88f3a6b51bde8cabbee97747be4382fc95e9719979c99099d1c6d0682623d3d3760d039f90bf9102b55252baf98538181a540685ffd9831272c6f5a2d2b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1dc6669723ac3c3a006f80cdb18c1ad297089d63277f7624463a02aa88acdaa32bfad4d3a88353ae3f1fdc1946d359686fcacac8f2981902e354d8959bc489c02bb48ee1d7898d5bc40f46b1fc0cb789f136ae26a18de78c911cc57be1887dd521d2e15786cd91ca4227dea93413e62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53232d35a26ac80185b7f7018ed733cb87836c168f4a2ae5e4a53d43511e27b866cc0dd32c4669777a0b09ce5fef2e7c21db302d45d0c90137e7023e887d00757fad8fa8ecf24391af96edf95919a46cde14fbdb7d181014fa059e08f96b50749a9d6b09433427b8f5a3b94c15a96a65f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ac49246ca75ab0a1ed2cff904a4790d33b2e4b4226adf088e272e13e4782c8a0961c961ce7c16de24fe7172ea0fd22097ed71f184569ca2c2905cc12450c0c5fea910bac1cabe2729ca4bf3fa668b079d51e1cba40b91bc05daad60dd64c5f43f9d70bed23959ae9e7adad9b82cc5c8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6073a52719a661ec0ca65b63eaf34a7e3b6a76e860555d444900001d9eca5544f718ebda745f694637541c288afbb3f4dbe80c1edffee1f954a9ef7ae4351fff0c156e30d515344b87bf34e8fca34a436c4455a6d59bf47004d973df63316cd811de5e9b5112391f7cbde05ab521e8679;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha030082c32acd012cd818852bd32ac81f1f35fac6a5121b4e7389895c5840a86dceb819b8c51923ee943dd7950939b24c9db7dd9cd24324cfc395e5bde03ce1f8f3218d4109a20b452a46c9be2ec01d855fc57af5391f115b199b5189e80ede2fdd472676d6cfc9dac4fa35d47bb66302;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6bf67d70eef2de537cdaa9810e306462830bddbf36c951dacb4bf40b5675268fc63250ed77d610da99698714b7cfcaba095fd887f078546b5928e9d33466f42c95c5ea927b48c76f1799be5230095ccc7801b86cd6a93ed7ca4f850199e68085cb527636b052a4c6084898a666f6151;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c2990fad194eb298704941527ccbac5d28825c85f24b07abb976cadf856f89f46c5ee386c25e854cf20c0c59d045fde90fcab07181fa2a5678f894690974bd5423439136014cb811a16b4780280c5689158d6bae69d8d63c0e12ee9361b5888473e16cb215826c8a4d15f1582944f1af;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf831648c36a9b508a4a01c58fae53397ce93ab88995640d86d2b5fadad5bc81b99523753d779568c3ddcf7bd92203daf743b56d413e6cf4485d08c3247cad44234980a40b80a1f283638a6feca609092355ca462632d05abc1b240a56dbe19466728ae82114474efc2983455c6319376;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb99244ae434349f165f71bd7cffaf73d2f1dbdbf42c8d97ffa0fe379aa7790a8b6a3f3d9ce045d0d7d04875c2c7ee111fb5583ac7e6028ddd10a642629268d9ee19f762e728ee6353aff668b5c3398ea025b63aa59632a687ddcffaa41c2275a078e2e487487468d3aecf5139361bce2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68a1f9316970cb36c899baea3368c5a8e7367a559ed3f362d424d43fa5dce01409c9cf2d2b95a3fb3a98fc20d009fd879371a63659ae55df7422564d04f25b51e2873d97c9b5091dafbe1170564213a992b79d0c30af917356a0fd180aab34aa018d4a31d7a65803661be6c45973c3314;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82926820ad6c13b6932e761879a92ab3b961e31a86aafe390249fa97bde9de4cd854933a862d18af14e223328f1ef44063e4271ed45104daebec2decbcc74c19ab5a984fdfb5748d3a0b93cba428503a11327444122b8b0d143757dcaf07b32e53846e37381aa6cc63e66dfbaf1540242;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f47958940f2da39c0fa07a5fd7a6bab39d9922139bc3194ebb773fcf833d55e39de61f7caa98a63365b35097a39a859e8f671143f8757d0b42c5769a9d52c93ea75578c8573d5b3c25ba0476103bf34c954d4d524738e581204db8df97a617bcd60a7953663db3cc46b4c106dc54cb84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4c507c9d9684e327f30b465721f59dd92f50f19114940e0c7ae07f3bc6ccbbe8609ccb792210e0a54fe062f4b595d004ac8302b47a2747e55907b6c72bbae1fdc82d3cd7850ec4575eebf549cb6c0757036e81c53ccc8db79c20d99d4bf09b854f59e577676fd2f3a7e2dcd7d03c4368;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1cbffc5dd4046c392176ba43f9e31a8aa7448cf21391b95e512ca8210e76faa607a7921ddc183c131d71fb614606e6a5a1149c9e39dd774498b680b23df0970dc62bea4c499ac7f4344f3950aebcae86e5dad4af471adf1baf55cac9bee941258c9b97133c7267c750d8d777ca1cb76f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d70724567d659d0f1635a6f69ad0effdca1b8a82d934570165e6ac90499d1e571d1381ab438a3a9310ab72efd6cb184480f4ab6139ee0813d3db71e742b648864a717cf7f281e1d9434b9750ae4d819cfec11fa5a36f3e87ec6fa5ad92f034483fd680a290a91d87913df9153f32200d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42449ee2a82e070900e4e94122d680afe7bd7f1f26ca84fd71ebeb66ba814f61a8773d311cff4bd5a470650fd0fa33ae55db5b85417d87214a6b97fd3506f1763f0f654f5742a57713449d4560c4e879ec2d48c518358a9d146e619bc9cf66b7697c07bbdb43f3972a8a1a9407ae733ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82cb16d7f787d1c1881ec5db58dacf4a474f69e4fca82b59767a7097bcabdce38d94618f3250189d0dd6be5793a0ae511b4397b58b657dfb1735ba084eef1655466a548620148f5e53bfaefffe77c411829698cea2e4d7ceb1d2c9daec0b192dcb89d133097d9ae9d1749cc4529683131;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5ce20cf18b3249a2340247d4195ecfb56e735c3a8f90c68496be61bd115dd0f7484bf1c7775620f979a213d2ca2aaf10130b825ba7bc0a86dc1adba498a481909aba5a392d7eaab0550dbf006a4db249b6eaa3dc345ebb58c35bfb01fae01322bd95b74379154146066a03321cf41084;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bdf13cbabb861dcfcd0d76c08a06316698efe7603ab7fbe6dd5fe0d49582556f8461a72fad6bc28da9fcd75ad68ff2d26fa37db88cdd17edd567cef3b622c3b7ed73307fb01111dc02958b2bd7568313c738d0f313b2203951449b595d1069f62456934106e0e376b526cdb5138a45cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h102a7647950ab0ff646ea1a38a16d5332abbc23b6daa12dd4e26538de07196f2767e1970e6f9a18282dbca2ba24eab02a6618d46dc2a3e67385b99f2f764573a571fd251aed40041c8c67e3e912a8bd1c1e364bb8daab4a1fabfe38829e784c11d5699cf3b23b0f99d6d2042d148bf48c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h309c2bc157bf7317bba7064a2ccba44242edda07153f086ba4e88e66714c34f8a8951714b553fe49f294fd2a49c57dd55cfe922097244b48ecdfaca8f4a8a1484bec153f2065ab68c2190aff822e60d777dc976a0bc3ff0cb27b951c6a6ded56e48da99e778733ad0539decc7f3c9b700;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc418086cd02512a80a458f44e5856dc09e065061a2030638754418745b6de0a51c0200a6490466fb52796e52dec08922b6cfb17d1d191a09678d109e3d8dd2d7d66c4e017864b34b0000e07d0f0f3c37f4a535297bd8a7ca4b117f661712eb3a84dd21413d7f8b456677bc7c2a0ee85e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h793429b94e5e761c43eb037df48fddb17418cae394abb5cb2654b6c2df82988cdc5308e69221ce61bba25cd5dfbd33d39bdb366802bf728f57f70f50fcfee0c0765eb0afc5331387d91ed34a4254d684052d81e4085267c3d2f966c7bff26db454992bbfd65296863daa66d0881c541d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b1a8247575735f278444b785f8b97b3198673c9fc7cf1d4aa7ed3d39577485ad0e160365fea869bb6624954a5713ed5152bb310a2c9d742dd8af0c39b906d40d2d63cf41ee49782d750055974bad55dff482c7b504ab466437885635cdd715ba6d9d81ea743587512682a5d34d223061;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59a44fbcfc72ab0379d4343130b57522700d0b6ea8f5eb89a56d02cc49367883c226d13356cb7a0fbaace13dc2ea22b4245556e54c06851515b5fca09f3aee2ba54763b872ebdab07f74848db2fad2c815f1514250a629eb5a9c7b199065cfd489c8ac2c4a840caea3043f6558208c335;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb993b007dafe54cc9f1cb000903ac0f93dbfe7294e075730cd8c405f7550381094620b171f9fe4b0df02a6c683ac555f6a8171f546999c262150ccf9074a0e94c35e22c7010ac031e9fbd87090d66d7cc6b25a53ebc9ad64176eae2436600b63e0dfe0d6d97f98c3cfc679d06529a9fe0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a5bae0bcd855b057539ffa534dfcd448df45c8df1042da62c5baa751833418db5a1271b7f74bf03ec124ea4395a047d1f075235c4ac36a99358118a4c5d01671ff117717c1f5f5327a3a3284ffcff20e52108f3d3b8dbddd3c45dceb24fe32b604918c17ea0ae36706e813c257f4dc2f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7752c495ff37965f9720e93af2f33c7188935a7d5b62b39d176fbe3009143810aadb22a7d3f494133fb354edd51f7b4260bee1dbd2e077e19a639e5a586aa853ddab7f5f2add93d2075bb1b9869e6b17c6f7bc0a4cca6f86ef7edbc520fa8ab6998998da4db40640e81dd79710813ced3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c397c0fb73ab7b152bc6fc40166a333c4a5813c88ab15982050f90610d01abb61673367f0f792bb41ad62afa37ca88141d3da88ee3e01b75a07d2541fb868ac1cdf9cdd7b578685e1620133543c19faa215f07ccf0e1a161f9a836d919bc0049c0e005ebe7fd69c87b803d97b534aa73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7cc42c7be75153a51eef346c10986736e61bb7a1e5a8b818565c3247c58f42b509fc2866914a2d281e00865643d75e8f0d0ad64d63e61db71d3b9caeec64d233299fc5498983437a430f981942f7f7abf4dd26cd14e594cc39b92defc062ee3930e77b788846bb7849272eae37f648a33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79a507c94cba9eab8a310f86578d6d13e48861043a0eee343e80229a9a31e26fc08c6c286b63b060bc5fd26ff2a1208b424f764001b09367cc590317ec4380d175334d470006262227cbf4a672e2c3f683e186a242b3d64bad0a59a7df8ee4ec50dce563c72d3858968808f962867a679;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h184072dd94c37f0f682784759da0ec93757f0036ee0bff4b2b223cb1f00811e7494ec37a90b02ab883c923116c003b023b2fc57bd7b2f13b8ea34aa5fb95617aa2f42f1156d0976dabbd0766c908d582944fc3f17a735135fa0c4a6d9aaef5007dc90fe68adf4e48c4882c7ac0170ca7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ab0bb69205d6a1fbf01162b424d16081654b1fe1722169421a698d97e4522dfcf436a7861cb7987fcd6652b9da119962178f55933e0326408f376b1e986974862a18d287f7bbeab5d4cae2f61a2378520f69693a7d65fe43ea6304f9d4363fbfb7b1cb3b7f5d32c612b5574594f8c32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30568507796f1c37b3fb3e3948153eca970c4a84b11541ad1bee2e504964a2104dc46acd552cd4203d7e3579948a58e6cdbbef4e065e58607b064fc42afe6b405148a278862beaa24eaf418b0f06803f62b5b6ec6d4333487468d8f5ce56819d7325cbbb0599cd8eb5d32050b77b0b890;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b1cdace708b6ab065b38d0bf0e8360620fdf5ecf203f819a99c06c72c042503fbfcb9f1b558dd7259e9520b71dcad683867e9da917e9221dd4f455a31c09d40459b16953a07ed56e465a2a93b55d5f6960a388a84fac85482edaa5257b827b05a7ddd65d9e0d9e0c88e18a6fe5623317;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86889b11271ac43009282ab14ebdab58d6e143b813120b8fb5d6cba7adae291669ecb25ec12fe98a9c74e5fdb5944e1b8ce3b0994a03ab74293b716d48fb917685b65c8f47b7a068d2de3f357ac6d8a148299294305b651772f34f54d0106ecc5a42c380dd089e90e5785befd46cdf0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4cad1cdf4f245d77e151cf68f5ccf049b1a2e51164453126717488fd97e942d89cdb6ebe977a8d79bdf39e90d71cee6941525b5b7743e30274c4663c445d775ea165d24adacce4af602658199684b54e82cedbbd4192223b970cfb58bc2393bc2df3d27751f9dbe5f0679ef0eda5c9f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3123358e20968b3d8db42632bf94378ce166933c8464cd35b0ac9a7eedb24bc0283fd1e83f4c5b2175c4e21164b348bd2f168bd6993095ace86740c7fd9aa8c42925863d564423cd5b4317e96bc4900a6c42138b814d894c03858f6c0a6453d93fbc127e03f0a6dc1388e8a5880a3b776;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde020f32da9496f3db03bde8200902652bc33a66f0f5236a4b87181ecee36214e0062562e2984afeff82a70816f09d506f8bd3bdc287f5f44daeed28065f72d9ca3a867cab87edb754ffd90093e0d01962de4984af10ad2462fd2182f1b2ac2c96eb01a3d7bf5149ac2751e6a9f802a1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he61af2fd061f308bd36efec208c30273567cea9644cdda77d2ab590c690fa471d95aa7d2d4e7f8762c37bb2b055756106b70e8a94f7f8b156f8e2d4f9052dda375365e5a6d3fe0844e30c48e495fb4486a8f658f56e7e89ef4162ed69923228a075383ed16003d3bf8824197c5c0cf239;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha213785921735b73694937f65a1f1cd4c053e6637e0ec85de5223143781fa61e698223d4b3460ba8235527add3e0cb6307f91782cf2b4243364472857a7550fb900e99fcdd6286ee3d29244f346a5824c9a75ef0c8be7d62c9708ccc59f6bfe5045f874754956a3295334b82700efd244;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8dad80335c9fc6774889143fdafac0292ebaeb556a98e47a76132e79c287cd8eef78b0ede390c48b11d4ce4f7d995e5951778128538070a3d70ae267b6191cb2d48df35bfb04fb833bf41bea7e376e48d0a96f6f56b20d8db1c069962a0a470a410e5bdbfa26ca3fd47a12fc1510a26d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a264ff455cf35e7bf27071ab250985881d8f932041d74e7984ed1edf99b1637ece74c0b8d453dd42f694b69b38a305c1561f15fb992a57a73ab194ef62f564bce34c191ef6259da96be97a260358c9aab9b807363bf70db72046ae51250379b38a9c6115bbe55049503696fc3a737a75;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f115a985f29cb448e9fe80f3640622c1cfc216a41dd2115478021f654afc57b68e51a0d7a2f8301a08c817a119c7ede6b92f5185d0a80f50f4fd4a0e6b2f75f3363adb86c6b2b321f154685b8a206b1bf7dc1841186efbc0c33ddb48fed905d33c9b3b56ec46f479ab13f64dba689848;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7569485d3d6ebfed675762598697817fd346448d9aaed444f403d057d302cb7b28b5427eab3c396e2014afd5aab1ba5cc2abd1f890b65216f480ad31354143ba01d35a30b91266c59a0e563208f5bbd1134a428399a2a7f919d92a036daea66748a50a05c1933251f8254a17e9ae2b54;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h186e2b8302c61bcdb8357508de9f5868577757b96b746cd9ef099e13d8f69aea5625746503b2cd7098ead4e26598f454c3c17ee180cf77c48618b4466ecc7f0860fb0414cbddbe109401c85602f143dc210d05d6fdc55cb879479e1307207c9c77f10655b736a2f04ca85259719935cad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3642423cffc40c92afb8a05b118be9135c2068907ad6227d72fd9839fa257c48b9c40020355dda97ba340b7def115f5a5770ca1002a2fa397997b2f69f8b5f169242c00717a991fbf56ebbeefda337c3c32377c2ba90cc2be16bf13e1223a31f3bf10853f1ba8caaa37d1dd86922dfc92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83c71814503640407bc50cc85fb173a7f3b7960c34bf1f69e3c306a9ce4260e4adefbf4119bcc1cdbd9a6bf1ec89202603b9a7ca82f070146f9546c4afb354001312111e49469e5605b08f3b0231c14a2f11ef3d190479fd0ab4999825e93c900b81a6138de317b28df535425be0490a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56ac5b3228f17782e2d59f699f8da5407f6510d5313ad3f276947095f80780db2541400fc01110ac985aaf0d6ff9d1e4f2d4960969db54e03ad71e3a344db85a3ccae030d34c6ab9eb2db5f7f9e589f7131fb64b53126f99875afdd6db703f3b9acd690e4d00176b71ecdef3c8d24cefb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72531b3e397ff2b402a45cba6510491744de6e1f2293cd966e4b738467f3e2c43d80f2ac428eb55df661f91a0371e594c97150194317d00665aec362a4c6f64df8e8dc74248e18986156a3a0a9e94e404f782a7053611c871e72d8d1357aa487cf13b3635a5b1f1b44d63afa90d4b8688;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7047273dc672444eac0f2457fd778db26192503fad11812bbcf307838840e7fc06fa4434985f80fd80dd0b157478992cbf7d09e30d20db3517197328242a511e3dbf7bf113ccaaea95ed30612ce48c5a8f083b8261da6cf844d769f8b16b8b1e5f385e736eb7f6ec1c6328836b94529ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9406da68a609c8b185eea55f343339d210f46f97fdcb93e149745329a69ae5050dd129effb29d13e07ef2adb65c081aeeb5a1cee26acd90898a6ee15f869e9b3759490814e523b911316c883b6736cd0be05eec4c939093b11d66907717028d44be311bfc121b502372ab6ed5549c222b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72de4cddfec6210b408c83319a1f49c0e39b2a8b7b902384145e4abcf3798c19dc68860c8dfb51f8a3fd3592ec67571b47ad58e13301d989a60d1c0500e50db2a6edc19808db5560bc4288eb4e655fb5fb2c0361422930d5504118f92b37c98d3f3f8b99be16dcfd0507dca2742b1e28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72c13c295d7fc2a539bbbc07ee4aed63797a7cedcf968185bf411fec85ef681984696cf987d9d8bed908d25c802feff7c06c4a774410900746db81827f98ed7ef1e4271ad83d78aecbb799fff543b03405f855325dbd41fbdcaed412383031024d4498580fb47f61e8e4fb4814873c42f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa259cacdd27c7f73a764834441051e1ca73dce0589c15f6b40fc16721036024f269d03d99a6adfcc270bf9e8adc0a484022617e8672e7ce432a423397c58915e12d358dd749484ae613455b73cef09f61ee0ced879b0c1b5baf70bb3f779b6f4ae827d740e41934cff48c55fce43529;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h512b438a8bf5fd9594d8dfe8de3618b7f0e504552dd99812b0e5048e7df8f68da47ccf5cdffc28773b8a5945626663f6dc51cc6abdb68c445c0564a99a69d76867bc5e9bbc30a23580c9e0c4995f3a16612750bacc4cc91d5a1b94b09932c576741a886fab65f7e21eaec0e5576bc961d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3db1dbeb72db745f8996618882d757001e783cb1e61ce3e513e85b088f91b569133f7f11ebccd918e76775654afa8ed88a16662550096eb605555edeba61fdccdd0739835c3473007610e6e0452b778834a790413256a878304fbf1f0c2ea2be3babda5b99c6f554570d6f85be53a4f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52f7e6dbe546a85a823b350ae7b06f63cb26ba89f1492bac4207f9b810c779f8f6bc54b68e1699114b6f8fd188e160041317e7a83a08cf1587e3f1f1db908f86cbf0d361a313a4ccb9809c2eff1a4f1888b6b4fe66f037088351bbc44b25e1b85acdb268aa2a5e7a233fa0d9041e8b8ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb20f1521fe55b8fea75f71a9033b232a23decffcf786c3024bbc0f0871127774fdb18891fd6d123ce92da31c5c2a5b94bb7480094b280f2cf3bde6ea30e421314d354e5a18dfc99b2bba15d5f26802906fdcf5fc2b0b55c29d0b7ed44f05d4a923f6c1b5b84e64d0cd5c86ef5fb6ff9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1145b73b054df6595b7cd6aac7c0c9181e06c0e6fafc1b683ee937db5855bea0a3283e73394abed4d497f082180b69b424e2088aa7606e1e08f618ae8f867b3d7d3318b5146a8c7f4bf53a1b6e3901f14962262e56800a1ab2f8a53bbcf457b67a12a3f791055d45efc49b5124bf7442;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h635ea39d27212f58b607d4d14d1758c391077fc15edbbd3a56ea1d5f774d1bed57bcb21512c71ea5b098e3bbb6bcb2a7e1e78caba6982117fe383470abb663c60953405dd8a632d207b4d23cb309f386c1fc114aa5481a490dc08d739cbd5c03461e4f5108650a7d8769e1eaf212206aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha19637de57344595117674c31299a4f943253f404b4d920f4565d5c2afa144e79b1fd9820aabb5372d83fe843f3759e5360eb3cb81d0458f81aa2a46e49e3548dedf1e07f789911477348349bc6538298b478f8fc15113bfec3367813ddd11c05ea5d8b64b001c0ffa67e40bd1017155b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2efa98c7741da206ce4f9aab70984a29211d2dcc1fd42d4d2b2186e47e9080b3be5f858257f0056ac3911a5847b1ddc2ea45a5be8717a44401e86dc8257d33bd97bb21181b13a2d78dde69f9ae550f1b66f84953e000a7de9368331b9c0f8cce89b03accc94fe5a89f7fccd405c379cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba62b2f223cab0b6c230f786950b78761a55e397cc457b6aaba52f593a63e2b2105ef31b9bb73bc133ffa79f53e2023fdee4fe5cb609658b05bd1efe45dbf37341e099ea067c0154bdcacb68e4c356ca16ddbd05342ee78579308b14d213be8ea302d8eb71d10118d2c61a2239ceb9ff3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h582bf696bd514a6cf363218dac5e01b9f53f7ecd18bac99d24960ed6715c1042cfeacf20e918dc158f70462cf6a79c4996f79a038d72f7b52a9288943a9d83b99513309bbebed45718dfb8f1ed72ec722cbacddf8e540d8889fd737962ac254b1996b317a53cdd62e1bc930bb00e01d94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h747b6691665879bf557425e003d15d43cfb5fbde649b649f38110e680ef80701c6936050188183cd73fd684c841576e8584ae605713b73a467607119602864cb85d99947521b6c7481cfdebe750f7f30d19c22789fca25a17f0a951c04ba96dac209603e26be7d196e524a7d8e4fc4e6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1f8d59157f9b9afa900ffac0dc9be077532d87ce95308aca6f472e2c5b2793b251dc54672e5c6f7549e33ba74b97224c907929ddb10b002bd04746a3f081cf49fca05a74f66b7a2dcc3efa59189eb3c784591361e1dd7d1a35742c9214c1cb5a570fc224fb24b7ef272061f0f337f5ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31e811f993162df32f126fc39836ee745b29a86da0db70d7074ee5259488db799d5d5b3e851a3940deb340cb89e0f27fadf3405b144ca68360b1ffe9d80be15e0daaa38100a915e90994d5a39d552368c1a08e08f63fc45ccec50fe73d938d668f97a712e28f381c92f8f62eafb02a907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc74759d835241ba28ac24fb432f31c64766dcb7f102f5ba9bda95371ac59245082a101445a22d594a9330648ddd3af97acbd8312144b4af482e374134c1f3ac770df08a034dbdf47a7b50c2eb90a1aaa3830c9a69389ea80a2196ff4cb0acc49066b1f97521f29211d5919521c3f96902;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a051db2852ed60e57656b94bc6c7a87a29ded66702a578291b3f425033cb9527c2fdfeb17961b1935591014b0b1109ad643b0a67232613f5134934e796bfb131bc949ba0e4dc93f126af98965993f80c1bca85bbc4a6650395bcd39e7a2d15a8c0a725342851c0169f1bf77d58d679df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fbb61240459603b55144d885aee604e60258c5aab68c1e90d00a5f78271959dfa3b8cf38f8d396d0d22531b114e26b748711d66caad6bc04944c766edcd4608d0c17c9c1ad3b1042215f46710551e47626c1f306ce32e55dfba04d5e7ed819b8eead93160e692cf0acbdff55d128ca5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e22cd1dbaf96a8e696ac5a524ee0a2ffc4c63b3525caa1b43d890efae818992bfd19fd5af79aab1f934808b678e07991b47ff0f570015d6b9043064a7697808771500818b1892586b3f0e7a85280a0a8ff374400a767372a423787525899bd4d8679d63db649ead96f2db5febeb2cdd1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb09254222df216edce9e8b2cc293e80fe7fa6567e487a9cbbec4fb33eb3ca570473e7fc7837e812b80e9bcfad3357994cd894db3ae6bf8fd42609f4a1516d0066cd7b9326e94364fd49c13d28e44abc91e77f37b63f01f786e990046b3fe0d4db80d5d77d4e96021c9f7c5ba9931bbfb6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1000b4fc21e02679dc98d1f4da095b9c8c4228242e91d05c10647db0998ef81fdf22d86cb224d0e8c11569584ec2921b63cc1c10937ee03c3c5a1a0cbb98137f8eedce3dee8fe7f49a79bb7037aa5eef64edc6280587c180c6bbe39408effcde83d059682c2c0f323a8530e397cf1fbfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdca65ea381d96658d7d8fbc23e91c595d8f344c73eb78df5804d6b87e557da7c3100427fb01b166f356f0d56c52a7563d3c6d209306d6f67c28458dd60b3f4f1beec694ba9d31b6bd647ccfa333634b750350005ebaa000a561a17ad05584282b8d8007e099d62d3ddd6ef8ce9c762b00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacf62bcee5c751585e1d2b357b6f45f465d562f8d146fd372b5c3d3310e6dcd43180b37fb61fe6f05b6b26faf847456374afeff539bb95c57e7d8d3c510d4f433f9955e3f413fb9997b478ccc97f0de5776f19864a3b6570b1a9cda7b019e7805e65f4eed9fd2205df3e6cf1e4cac1439;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d950892d0136b7d0c56c08238ccd0cdb5a5567481cd71f35bd47869d08f2d70b326e481248f4be0a430b7039f0b60ff6ef22c66506075b4be3b26ec87e72c34cc806429db41015f92b66abb402dfe5f476ec63bdb90676e0426c02d8a67a3674b0cb5d030dde85bc8038710e0c4c7b1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c551ff70f387be1ef27b536e20ca232dd1b218cbae899538dfd9e88409c2d3e685ecaab3914012a0dd321b2fa0fb03a1e1fd8157a4fc6a538400cc2cbcd155053a4778e9e60abce1d876ce4df228cd54dffeda4035a6fb962bfd0ac3895212879426f62f9cc1f502a1fee80cf96fdda0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2384ac5e3f4986041d87e1d316f1c44ea5d18453c7e7080da995788e4b7ca5f344a59a793f648b61e43ceb1925fbfd6c62194c8044671edf1494290b5e6d581c6611231be947f088450b57e623eb0b2a7f00ffc88d4c1fb33571b84a68ac86fb94afb235b25244cf4e3f9904f170b500e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95e85efef63987de7126b1b27e1121f832d0b290b6e5103a0f19272952c83a77d909f00e6d8b90d9d2743f49e219c8a6ba73aff5587bd8fd703216b3dba4f471fadeef802f6977e73a9b3053cf0e1609f32fa5839ffa55a45a36476b77e5b9424ccd11ae433f23c194485d22652f05b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c7b2a16cf309dbb681a42184dbfebd095a8225ad7f5a7314f2cb31f946a7e6d3b4bf84d72d06491edab4ad944b6758a343b66efdac17f505f19e672d356dea06d292ee516a61ea09b5a4572062a0731f84ce300d8d1c235da5caed5476c8facdb2facae65e65ddbe1f8c1cbb9bb6b968;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedc1f9f627202f305ecfa19da57df5d8988a6d5a99ccb6857937330ae32d63535e33b5fb5a512f17de97ac8c1b238478de9d58541d5f837bbd294dc57d8127a8f3f2232186d8e801a66f3ef01b07f7f8021b2c31e7639b71707343ad3507cd2dc9bd603ffbf261b56d98a08b2da4a54e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e0e977bd4981be213e2cca4134be12c5d3995c1ad981bec41116a8b6e190a9158194a3a8f990447ddbf64bd93226018a59fb19783b450dc347f7ef6a486e63cdd4917979c92db2c4e4c8d8c832096a787308e1a69ec2e87ed5541b519bf83a85390764200659c3e061ab9b5f435e01de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9f8defe60e9b16901caceb6ff0175558cb4552ca8106bae8aa15c4d9c8540e1f45ec3c2d8694fe65c8d4e529bafa705f60fc6f8c96c54dfec7850235e571cc236808b72717010e018c8961c37a10178cba15e03330183c6d09d2fe6e6020dd9ad7053f3e650e16abe1023695aba52c60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f4e16d2aceb355e189d77f3232f24c9aee13742924e340154f8b999728647ca9bd95f1576773b9e1d77891bb726f81ecffff4d0bbf12ff767a96c7d7142729f497cfc711e22f5faafa7d8473a22828559ff6902356802387f3ab7303e990e239294a70be83ee495406a89dc4db58c02f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h599c38fea82a2b8fdb314b6b8ce02f090eeaaee4a3010a991e3656941f4947abb59bfc6f73200ce75563e4b39e01dab91741a1f0637a5e3186881d0f6cd5f6f2b69391cb749713a1b3cf603486ffab10ae75f1b24f24c00ad4911155c056839310932ffc24c1d8cab4867ccb05a2aee72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6207e2388154042078427ca38804e3c02d1a715ab3e9825a28527f04fca5ce12aafb95a718bfe7743282291b521cb9aec42da41b62c4651edf4dabde9ff24c74dde36f9c29059633aa669dbabc71e2410dc85a8de9cf600c4cd29ae16db5204d51acbe759d0b42bd726cc0576e957dbf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54ca983bad8da1a1421b6261405eab8f4203a370bb0cb84200863aeae85a1c73727cb1f65c4f8cf6c597bab75ba107413a83b76520f9bb07a21883d3a4627fe663507e6fda12dafd44d67dddb4722af78547d28d7068ca8a464aab293589316e3cc95804f1086da224b261ebd61b8d421;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he61423c396ceb1e6751d98f1129837fb77bb8623b57dd70eee76ce60ffc97c577d256440621f08ea5aa84504a34136afa1b229d0d54af375e17fdd30078455a8d372957ba0c075010bfc06a34742fd621883d4dfad4b4a268462999e67dd5454dd1a1a31d235fdd437b2a8c992021ab35;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bd89e959bf1c2e3fe1c060aeacda68195a709a5b1b4da40c7a80532450d9202e8d2c6605b897a44e4c6562a87012b75df18c4ce737c3ab7122e680bcf309497a43d1ad0e0baaded67098bdacbb38573b94adddc8897a1e768394d3e4121340232ffa31a301fb132bf0640492f9053394;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9393200441da57b05f64a51bd7b3ba1d824de5583e0b6f89db19cbc5c4450a29485f713a56081e254dcd672107d5dabb7624f9a4b4a493d62bd0cdf8cfb0b6cdc6905af3e96ab2b23268b78275fa73925bcf2dea95bc3a58f3fd95bf47cb47c7cb78241a41d34ff3812b178246f2c0c62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69b5b068e5d5c18fe90edffc97b0ea02c2239959965c33589e4f705da39d6ace2b79c347b987bd757107e536bbe501291e2ec98f0844caa9891e5111855ad9d993972aba7f6f7b0337aeaddaf0ac575f4fb14bceb61320b720e1fecc97590c9c6c7465ee3ede45877ffcf69a1d8710d9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcecdb102f3275d174e9a293305edab6f0e5dc94e925c4b18703f71aeb64f7bbe30a434a7cf8498f26064f2580fec9266047bdb81a2feb617189c3bb6b5f7ec0e2e2b0b75bc3d8ed82343db489ecc2a7f4f84fbc6ebfd4a2bba73607a84f4bed811566f3f91ecd80e35970da726b98a50a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1efca670090eae865bda3a069ce88e826e31a0298735e016b877104112cce57a7082f2b751b0f4628befeffe9968074fe2b2861af2de6a23ec2bc5f74a86f1d4547db886cb1508d55245cc6e781820926f9becb31e305178ecc0ef06365ceb50d7004a6cb3e27f2a77c22f929a0de842d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4d91d770b14695c8c769e7fe4c417a546f4a830e5d41d301bea3c8a92bf6a716b4239bdfb4f20ad0f8075d724cfaad29e95f417b2681aa33557bd63d1bc0017b8149efb84094953bb2478f17e35b77c650ab4b913b9ac76a803dc91b385b279976ea7a1c8d2ecd4600bb6437e1f410c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5654e1530f11ea8db53b869491fb6403692707074ef6d5679c90d662afc095f89657f9caccd4835022801bcfef2a6fe7ee08b418ba08ba0392fa7e3255c526dc59085883689e7d91d2bf4dbfc336629e633260e9bc871a323c78ab38e9054ab4615ccb831a1b025d4d3025a3c5726ff6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6e4a3c593f889f2015e839c047081bbc9a62f4faed6f0c154a158299afc7439bef79098e2927f015af0a6c3eb6e2a20c3f239720ab1615e03a2c81a85308eceef2e426e39cbcfc4177f6df3fc14b6d12edd3bac21425935a0304a975cf42eaa9ad76c437369eddee77ae17297c03a543;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd09c69f5cdefc94d974fcea48532bfdf10e19841a4f35158be0c206947496510afc29f28c0c27dee3fd5faf9b74bf11108031050b5d1856fc5cb37269867f34f3464d4e9e1678d3c2903e95a10f0c66f69e43f9290c771a11bbd39d7ba7168120efcb662455a8d9972f2cbc8deffa0267;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbdacab8ab06da6dc8a3d73a11b13ec88242846102e0c5e5a680b694026aa2a32405603dc47815a3c9533acebf196a4907a4f741bb5d918a52dfe6e2abb00abb0a9007237229eb4a7032cd42d3a9844bbe013d2dd639b48fca0ff4c904e84a081c39566b915c32d59c25b9f5b1f0328d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10f2f46ddab27b040c2575fe18129645dad29b9ea29371381da308c7f4e3e89b2744670373a97032313f4b8603109253ccfa9d19fa7501e52796140a331ec7fc7d12e31870679ca5caf076234c4414d1137c4e77dec2fa07b328fe942394d9c795e262d5689eedbee0abea4a0f41f1d3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h512713b1d9da6441edc16a2fb737fd636bae19993c2f549a6e9731c37ee91f1c0bb1bd7a28eb8b6bdf56b4974623c2ff7d6ab8eedadc296f92068f6907b12439d18ab7d781eef7bf6b3dfc0682d2c79b8258ef659be0fb888f2e15c05523473e08394ef6f6a5b68ef7d549a9985e14d4c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd74069a6c1ec899eccea2aadcb9221fe5b506103b9c65c0c6a23569ae402d247796c79a4b7814d2ed995fc3437a460f189d33f19c2de907a3eb8e5b9b5e2bc7360b91dc5cfd64d2124477e10b8eda8a36d34c345e86763ca34bbfb8258daf4a73b3444e3e5fec6373d2ea229a7c9c9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26579938a27d9f3f6f797ecde1fe29193dd610da97f902ff646feaa80d00a73381f66211c6fd8ff7f11f1ac8252639b3011fa3b63bc6c3a311eeda2d5f6029e533a7e618453471f6341e5ca816d8a8054f8e26d84de26a05d32bc8c4fcd6c0e7d5ff3df848ebc398a62e85396e87a975a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67a7633e71edb8d36bab6701565d6074f1268e708d3dab7b169e6dc05d8e0d818a6dc0108fbe0b60122290468bd6d6021da63842c3ce910096b16e4283c5523b6a584b93ef0d0a58c1b0aac51d14af8a2c9a4601dc20e9affb2119f1002d86e5c56dc10b2045d2f48d57f64ba266a38d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59ad67acb8931a7ff1b6126fb775286da8854785e111491efbf34b0c43a9f8c7e6277fc06e4359086d1c61e3a61a67ce3805285e778ccc1a104a0d61f57dd30bcadb853825804e97679193031960b70430955d530ee3bc76fb356d15adb26b39880b9da397abb4267a0a315a855e71521;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bb1d0cfcf82e63895156ac4beed3560bf0a3a0c6d81a609e3e49c9a57f83232676d550b2ed76e200851844402644678c87662d1368016924ccbd93ffd964b5f6b25762c80787036c1f1e2c69e44633977fdac48e2f65d10eaac45769dc908affb64e9f0c458348d0199bc879f87f5de3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e142e8f54087700d92d546e7a9f41342bf37b94444d944334e8d6a511e2482b4b3a75b4c5cc3303b66df3575179e13c435ae92fc9f70425f5eeda53423ad86a6926d2ff2c15876835abcc5938302f97c81b88cb78e8a62c3849d9101b90a840a79f54744be32e20e1e630626c92504fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habc4f6390e37e4c9e1e597a46ea8d0863ca40dc7a9a4a24fc33f3916b43b0bc16c239b74b70b23f52d35db716239c83d43d79c9e1cbced2aecf3f11aab15740a701b0d4290a1f43116761d1adc37293071ac76dedaa03c96fddac83ad592dd2459dfa7b73ead76c52966b85ed8d1afe19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6bb030b8cd75bd5d3143441829d0da49d4bc2c09eaaa3aaddabee023ee29fabe1a0dda89444f676a440edd468e2cdcec7d66e1b39df9f140f1a483ad68c69b8200339541f462095c3a098744477443e99d554ca8d87ac2cb75f22946c7c7ed9a5d3ef34bf77e2e1145a8a9a205d51585;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8db33dc481ee19ee472d2bba58bc4546c15eb5112e8a853180058dc9b7570e1b35604d28e04f2890e9c79ac604429eeb78abab9e6465fc18e679cf20406ce3e85b03996b0b429c0d70ba440a29460338ca05ed5147282bbdcd3f996f66b02bd83e9a9e002f81fbd25b3b6724972de2162;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96f8d0716791581195ec4423241b2c850de39c045a59dfc79eee1a812f02f179a037df237eeef8b89b247a75d4ecf80a490a285446445a573fe9279415495deecef1835a87412682931363b4ce0febea94c85608a92a4bb3067f83f758a4c8ebceab204534545e686ced66ea20ffbaaeb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32317b474dbe5170f63a3d6a1cd16256e4aa15bcf0a72fd4cb9b83e3d183f008c55572c15b061dc54ecd2a247a8899111e16cafce78d23b64287bcfe362140b400ba564bc17271915bddc047d95a429f81a6d8a2c675a276e2686149e6ea8e297dccb9e06d6ae38888d689033ff5ca78e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc77b1ef37367dd23f320d6397331649a6979fbf76fd6f97d8c2bf7c03bb77f25545603c2b7363e1f7bf3254d97c862a8a89eace2c9ae93624c3938964720bb37f74ebf02ee7723006477da606ef5c8d82b241b26ef6750cdc3f40ed5e5117e08c291bed42f140a604448c10cbb3a9a30a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf32e6446758e2a9fb79de3e63c29df460f5064f1d1dd900de6eabaac1d1aaa95caab98b2f5718a6e5be76db3eaad30ec0a5ccd2785b13033955c4ba392648472763c867c43a4ef5a5c7e337a446fa91715955d1b2dd5b5203cf0fa918fdf193c428b4dd0b2cead6e253414ed5aa2f0e05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a829ae1cf5dabb7df9d0e6d4851420801feca575e8811a073bfb0d283a4d3ad4a5d46cf9e43cdb869bea1f5ba1054dce02d57c442dd4df0721d1259ba2ff003b4984c27598f3db42bad7654df04b5629f4ec681cb885af47b2bc2d066bc0d2d0f9f4ae36490e2e3251a1711c2cac11d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc32d98be4ad37cd3edc61d008b7c08cb0e5090a6da231bb48c2d29bd206fbc94a9a38973175a8301d7de2a9a40307e4cd1bb60987249893afa7c4f929b74985c495e20b0d3ade6a588f1a4c0507e0effb571da6ffce75c11f24462c308f4b89b51d9ea0b15bab5952c267c7cdfb462626;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h316697fbccb10dd821997b07ae531a36e84774909c862a6301bfadd2e0eacb47a93c655296abafe50309ebdd679a8e71270dae12a7eb7045fcbe7bfd13237439bb53205ae8ff6bfbdacf3147ed72a245143399bb7ef9e115ff29afdd6b5b5f84e673f412fe77859a973c3cb92e96776bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5af22b6c4cf3cc649743de34d141fd6f1c8583251c19fb373784964418338e4ed6b9436b2dc05a6e6790700bc9b1fb6aad49876b7a689cb264fba914aae6e81575c5d223d328423e5f19815319d8c2a326059fccf770d545256e4dc49a8ac22e5206345c55dc36b6ba1f6d149b8fce870;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31a92ca4660bc862ae7d86a3c81793dd3bde3135454cb41405f2e716e4b086255040cbe6c65035849dc60cd30a9fe4e53e785e05d19be588c55a0b6c105458cab9fdffb6e7674118c38e67e5de8c2dcdba49aca60caac22c6c94b35bb8ab59bc7a3fab180bfe60976ce05447fe43be7e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7535f9de3749b8bce9758bc2da961ecc4e102cf9cd69609b5b101c06d05bfb6bef77801ffcc018b1f528508c27fbfdb793a7cb024f414bc6372e82f53e190ca2deff5a8b7f2baa7ae6b7f98c57131297ab33e4f6ca6c1a0064c84b3804f43229e53963201cd73540a27967f14188ebf35;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc5e522f9805763064d71ffd6579b964abafa60e4925e2dd63856e2d67d695da75bee6f5e72b507efdabc98ead6b484ca038f8355aeb70e98823eb0563ba29570aff0422123a2b22a4b4abc2216e5b5ccc67c0b4e8ac65ba83dd6a766be26d5daf86fd9e830edac8e27c09921ddc61bae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h645a9441238fce01eabf6a8dcd3c1c49f9664a5060106af64e7d8f0f69e83e8e85b1fb52b30e4631cbc682bbb650e36992619b3f43e228c273e871cba173ffb907c4acd01295e4f91bed02eb4a2a5f740f6e5d26c0ae4839cd479de0bd9f6048dd1aa7d179390d1c11725576f76486cd0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc3ad04a4623c6fd6d28cc64ee0840519b93ed0a101e100c1bf60a369833ca35880a77501a6736aca2ed8929fd25633fb6b43c43d43860029401062a1b98472bcc14ba2652032944e1f2146e4ee64e767598da62e7251cedbf450c450a478be0c5245d711a144b073852edafad2db701a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd920287cc022946e88b5d9ed7d9246e3d2f03ca21d5fece319dd91c7499d9b57a2ca1347ae6ca457256669763464e08b5dcfa1cacc2dd47229e6388a99e03c9d7786d26be59f2024c2d43ee8bda256bdd450fd2a8afe2e3c762156c511774484a81c8c31ef16912f4888ca5dbf909ad1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68a92c558f7b5db82b829039f694a5071b1b06269adf55fc000646fcc6374dfb0fc805fa8d62b7af6c84d60316e247706825c93a5a6103aaae4cb845b926341a9bf620186c4669e804106ae60a4517ccb45b76de374fb5d330a821a76bde2268bdd0ed2e0c8f34ed874da52e113fbc146;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68e6b22fa30671590bbcdf05c21ac3e526fccfde55cc9d799cbe3ccf7bd399a773f6c4383c6864ddf376481ccdb5d42b5b4ee4d55e6d9fed0a553d7cd7ea1410afb4b5a79f83671f9b82d6f6105bf030dfd0a0f05304b6a4ea8451db039e20c92926a89607fdafb2b4ea232e0e30463bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab728969da876797f3fc74ce451b2e4cd3215c13622072945858bf29c372f680af0971e8103caf8a9947b2d7212a2f47623c8e01ddbed18122f860ef74edb872d14681ab5094c439865274c66d679daf77e503e33ed13c1d950727c8354f87ba350d7f84cad8572ee94e1e9126b8aa426;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb383daa8e8dc048302e5b14be768989c8df0d6bcd23a688ef93eaca18b1e2904a2b5ea331a9bcaae25fae4824005cd3caf94bdb8e6df4a973e35aca94fee36bf9200092d86432cd4d0f2e1903b7d3db65880c7d0d04e13eb676d731ca116d7ee0267636e9e9a6b3d54c59bfb10dc869b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f5e60f452239a782b9c7925fa195922b3ab2dfbc4cd5404f836a914e04eb47aac18178c4b32e6f6142f92d1fc631ad1437b0f31dc9c3cef75609765426f43ba18e871b5433a0a645273ead8bf5cafc35017b7803d968458fa1b68e1b39dfe406551a746da639d3e72421e79bda0a6bc5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb55451822896dd1d7df97e9663376ef533ccafe95fea34c240b7eef1a0eec62ed6cd3a3ae61b2cad5c3db8ca468d688a94bddb9b8e04637128856c9fcee17a84a0686c84a45245059255b894380893b89862d7593a65b1a13002141c8c5923789a98b02897389559fb8e6322f4f3b6bb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86629db65c0f79beb120fc78f7fac99f945d23bcb213a67088fa49a8ee1d7997ecf0098fa37fbebadce410cf6cfe21e0ce54ca6ee9868e3f4646f0e8f8ddd7aec530517d2451559ea2d674985e26402cf16873c7310c5d090c137ab02c1f7fb6d3da715632d15fc3502f6e1e07ce3a11b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8207f84aadba1bea608f466fe8e6e1fbf47cae696e6ba00c7f6792bc597ad1761875ba0f41a0561ccef60e4f832f159828bf09d6974619fbfcea47f90f7b82288de0f59bc02ac8d8dc58dfb14415cfb413895f3852c3d449781fd064fb1e88f1780608a71f4890842996e27a440a2a00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83b3758985103e629711e771cce51df5c5aae7372efcc28c149cc25efd09f0850d9e232be86059da867463fa194dabf8bea65b83b4bb1d3dd1c30729b9731ca4c5f20ef008eccfc6b1104327750ecd1f618cd6f567eab702d172c6a73bfc3769f95ef97544b8e5f50cfba7491b978135c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5028b8131b47b9d133355149e661a82838b0b04c7b2c6f413700a6156581e27e3a5d916b8c8d018a73feb93614a84b1d397b747ca4cff28cdbf2715b2de78738584bdf691ecf576c5ab21a073a4dbd70e4e19a3365c1900b1558cc1b7b35ed899fca546e3043cae5eb9893e7e6c7e6c03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5688b0acd2ff1886e402f41d4a07503043ff83a8073394c0faf5c26718f8cb61f9c11d8c991f5d0151e8f0d27cc14440ab48f3e29a46adcd6090c96cb502246775fd5293edb7e61b559ab1d38f0c380a59f19b1bf05a22883442908748319ea09ac177071a69991b912559a3f28996f3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd59e1f7fc27f298832ae092dd98f03a827b122f647af9a2edb05f962a9d62c11aa65e4b5620533662681fbec0fbeaabb5e72921b101f37cb2187640d58135cea021d18024996d07a8ccfedc77fb664c2402fbd169658c8fd084821ef06d2fc1e0c6f932ba2aea3eaa12a78a26cdc4e07;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42ada810dc2b4114ce011459800b00734097933f91f88a6c1ad9e640b161f6f084776f60a2b7f4014066f0bc76630806ff254b0692a1e17d494bc5a670c9095f2fe87768c088bd9e5db8ac06b073f8d9e3cb0d5474a8f5160ba599386213c78e2400f616b3a3d1c0617882595f6943958;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7832a96fe9046574083e78d7c05fa0c42917585b89480d4ae000ffec1a84c38098234f6e8d89bd12b6238842e89c24f8a1a7dbc2fd3e12c31383b074494fc7909837477f2014324c0227dfb45988240f049e281f4a1407983e2bc5343ad799491c1cac80b3a7f670061a084af1c2cfe73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4119f0d7987930208275040fe9cd86a193fa02e181542e40029fdee935ac80e6cd59ad8898b9c6a973cab88a4d035165c2fa6e3186811c257a4288ea4861646ac575ca04bef2b094cb3e720bcb3a1819bdbf6a1fd7c80bc462c0bd12f634d07190a1088fb1d3f8e83ed8e6712de34a157;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaf28cbf2337c4341a37a1cdd3cb138af6455c71d1a81b50902b4e510518962839e121496b0b83ec152db60474be26f3cab076c011e6f6c4023cd81e5f409c4d5d41748057dcd88204ff242702938d3ed2d5d6106431a827a35ba067838c9d5321aa5df48847e42ab718258b72e9704a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbea61e16bc0e960205d1a23c35c302d2cb194263f3234022e8eed5f4abdfaa971a402a89ffe04021024c4916e43a77b17d75cc762f4ebf23940f04f038c16c27de0f646cd547a3d9bd15cfd6e204c7dbb0e806e3f2656e506c97169f37602fa8f625fa78b625d1c4b1daac777db3120fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7a7e354204fe6780b3dbc25c0a871bf7eb2c1cc04854d2631a6e566558fe8120d39b879a25fc81b97df87ee0adef4de639261c697db49fc964fbaa1154eb227c3a233bb109d9f014c787b14475d3f06e9985b653aa236e4419f3dc24a9e2d6c3d449acc0f1d0c68ce2096729dcb86463;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34032d01b44c7822db438a1775dcecfe1809b62c998c42924c226ac50f40db4e1a88ea2a01a49064cfed45acb3b045f9e5ea63e45e48daecd1117a928cff7670204a7487cb1f8b456bbeec7d941043985d3f5dc829512eab9759ad72fa25cd98f8fd79bc2695891b81841ad0b287de327;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f3e602ba8308f5f96dfa56b15aec765bc6bc918b876db22e818b7a12cc1a5ec27bd2126d64e32c75f42a3519e97c825f07e98026639ae3b12200ddf24456380e9b92bebf9c9ec95d89f59ee3557412c013e6fa0098dffdb3efe2e629d3ab8eb8bb9092bfa943c94f5ea010f0077d7d14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb491e85153ef823063b29bc813d5b5aad0b3749c59333ff50fa35f8f9cff6d2857cd65d0e310e5d3fea39d67c845d28349684fb7d5d43cd6696b2917677b661fdbfd827ae698198fe576fa0f565d33b3c6be566fd67f6be23c4e2e05d77399f89617321cfdaacd661ce0ea8fb552c087;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ae366abd0450ad6a098d6c9cd53ea97bb19836b1f157e5e046c422fbf96421d26c8598ff758b0a7f9ecb0770d750ec2eabf0455130fca07d21b7ccb05f4f7923e6377006ef13d3be46ef23f00433f1aaa01b05302ff333089a03e4d7a5508d161849eeed26df0a8e910178da3ca66d97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8879f98bc6771b1a9f9b2d720666846ea18838eb7c3843d07c01fcce92299bc630ca5b45117b218d8dda5d0c5953acf924dc02ec3583d8d893f437647e62a440573ac3514f8246d2e45e4af83abbfa64c37ef0e981af88dbd1beb52d174cf4e449289e1d1afc2a62a191f1847882d2842;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbba6420b152c3c38ed07a8026ae8c54ee296e4103894644b240b44d72c118f4e59600a9c22d0607791bb5384f32215f7da44ad0b61573a7294878478b3ec1f9fd2ab281d77dea39954ffc94f0033f19ad461ade9406296ac0d0543ad994248496c7f7554b1f3a2535f8247290e25edd1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25852a9688845c5576699f3afcf4495be19611a4ad0fb43b98cc5664a047304aa3c60d3bf7a297d05c494b50a5703db27f44f75f657bd2b0b11cfe18769a81ceaf53bc9547b38d776bebc51a735ab5f16a27858bf1079f4c2b291dc14f7d8258c7a4c6ffc6d45a3c2defa5b18cb063292;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2718815da32a38ed168ac09fa9128279c9f8a83807ebfd0b42f378ad72775f5059f61d27affe2325c9cb2d520f81138ae7a2644e6f28d23f193a0879262ef3d011a797608dea407ee8259bed0d4bf9722c03ae09cf2f7c1d3b9419f3ac9e24d3bdc622caa5ddc2e5bf9891458fe11127b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd090e1a9359a1fbc4645e93974933414b86e414f3560fb48886733c694eb8153b5a6aad128370e5e251077a5b5882b204a80916db2dcd697c05c6a1b353195d6bff04a6c7bd93139f6b7cc1d245566fae1d51a1bc3cc584dfd3b2bd351c5a104c682ae5cabd7fd046de7a60c49f43d785;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4833e81ea44069f6f26c642f83bebd10263dc104e18329d6acdfbc819cf9f606198c49ff9f5c9dd06698b5b89a88c0388fffa2235acf330d90efc54c13cb52674c858039bbe40848c5b86ab1925899e513cda3a464ec92fc35283caa2420b2fd120407e3026daf5edacc75cfd3cfc18b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57fa20c769532c10f658c697ade3392f97a3c91224d2bf3bb0b61380c695ed8bf91c0d0e3917e08e8d5e9be63f26ce0cfa49b14301ed6385f8c438bb78b68b897ef22673b4f700cc7f7c05155a58640ae6119d8003115dac902f8f82a517b7d64ab7d70a36db54c1cdf85410ec4200a40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b28ae9d16930ac6fe121611b57754066d42c28687eb41672858bd75d7bb0986fb567e35c03f49d45cd022e2b3326333902c311d5198afc0ff89fef942071733901f13ff12eed88c5773d2895104062710fd0a0efd20258534f4c42bef07c9f89e9065e576b7f8507061347de8ec1c3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h925ae46fc9954c626966851556340dc7da6504ee8619fa3d27d0d59a3ca8b675c116ffea191adf2948552836fbf463afece94fd21b6ab55a7c44d6d72c02e9bcf88ac94af9d39acd0c693cb9363593fc3e1d5075c4ae403b8bb4553a379ea12f25ce693462022563e76c2e52842c66b1a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h816e5878e4532320f1e0c69de57e93ecfe960ee70d1cdd63ebfc7ba1e65c3dcfae4057766ca914a2f340cbcbf7c9b20ae1ae9683620364aa953e50b226eced9d10961ab346bb1895b9339d683f690ac3be479abd84d23b6a8c4f678b686db54b4e5cd4404599669447ae89eecac26968a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61dc26be9e225891f28aafcf9060d97352264309f7398f3ea28f393f76235762f2802f3191d580192384ca1024f34dca8a4942e56922146413c8a099c460f3c1e6597d82511a2ae2ad5ddcdf6a24f4256d3602b227f45dfa89e7c695174af3f4ba9b833c16705c168da072b4c80d033f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f9221737d9569bc3e066e1fc974190ed78a91c8e91e16f759801c821fcb13fd04e3bd681da07c615ffec6df158f6bd01426dcfa8bd461c3dde05852319a0eee0a0e633fa1de4c16f8f3cf6ad962720f9ea869cb096b604da291ed45b6635736ba3b604b30b45fd5f358ac8aaa1c222b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h216623f0d11c338842a7c52471cc1f0d3128822919533b6b62bbc859af248c7d5b14286fb8367145080bf2dfb4b2949ab2d0686697073f4e60439cddba42208e35fee8a847652ef85a97151733cd44b3946323bcb56abeeaa13c123a5e675be7aea0d53fb94d3ac340d85a3596f47495d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4306ad8327e07cb031b9a925b821c1c406ae6a5ea7dacdf483aada23275bf2d9dd16e16a5497117ae8202903c8fa00081d8a8dd133dddaad1f9d2b1b13e6d10eb6ae62d5f846dcbc6a18ab16fb49fa9db91dd1f89a3f14219ac18c511cf8f7267827cf0b635c39dcd8165da38a5659d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4d796314861da0fb2db916f37eba5e8705a1376c7acdad30f61e83815a17f2aa87cbe9ee660736fbbaf21af5dabae4476fe27ebe65a498c2eb391d3ece13bb26abe9f30b8064601936d73d7432cd26fcadb4d08ffe4921613105bc8b8545c171667f9b6bd212d0f582f24b6a0a36e0d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3980d2d56bed60a9f9af9cc56f8ddafecc7406bcd6a22320064871cb5daa4459037402923948939fef9d6d20d9a406e5b8994395d207ef1405523636e275afe409e752caaeb69cd77aee6178f72fa419f96776c8090910b8a6db85fe6aed0ab7fc1daf945eaa6e94ddadac00a6c1381b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67e6e9f8d4d36798757f132873c848ea810768cf59178d1c3e35c069eaf3908bd1ea298744b6b758f644502b8076a3a27782070bc8eb128846a3496eeb40499d3efcff73aff537bf9c540a31936bb1aa44023dddba1fec823da759df8c75ae139ba847136e267665be5aab94014d42c22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1648d662fc7ae17f00d65956bd395b83061ad9cb15fb5219128171e51d375476a38f0314d3dac25cc7aa638313f414ef23c9c37932bf768de3d247580314452758fb079da5e2482e6a4da97e60c89e25fffdb1965e5ec7af195efdd99e4862320a00bc64becc3de461253f1659640bf6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h402f66880e315f6e7bb145ab29aeddb8893e28f4184c8a7b2b57a8ebfffd34aa9014ea343c571f4558c43ef6ccf4f7a07836749f39b529bdd04398e8e1d84838a80a6f8b811dbe5f3244e959c5ac8fd60aaccc2560db5f9edd7ac269654dc3d864fbb04c5e3a1ac6131b8bdeb5e5ee856;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd091ae92254e6ebc9c7d09a2a878a629bb9b0f6dc356c9cefd66b0af491d65780359dbc5500ee0bc04dc7e36d27e0cfbdea5a3df16c52ebed8bc4a94772a7cbc073fb65cfc9f2fae965212d8089b48faa947676326048166d3e994bbd87f2388824be2db4e0a988afda91db68902821d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9563028f915cb05a67c58f9ff48ca413b6bf8bd32a6819c1456f253324802ef215dbcdb8ffd2e05337e8c800ce28a583522dc93779dedbcc616dae24f6465cbe122ebf058e75ea3fe9bde4ad3cef3254b2242003b13cea0cb57f3758694032d03702e4b677d0fd9818ee1e04aff1a8f96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd855b4a6b9daf6eb4995067b9280ec89c24ac33e9791e8f15a6f4e86c55f3fba24ceca945c9cca034d9b5d3738e21cf657ef2326e6cc06dbc898172fee83be3336d7376a231ba245da28c3fe1772afae85f7c38961dba036eeeb06a8df68a9d4a6b899777cf2ad07277f006dad6e412b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64e9c766e3ec4b11e97b68f045ef18e089366b7e074639001f353aefdfd67679beb05df4d015ca7f77d4efcfcb31d455e70b7bfbcccec67af1d4b1d94f8999a80fa3b77302df38044d44afdc3e3013a8aa7f23c0bb09d5e9178c17f1da065a0fe9451dfb153d5cc61d83dd097405da0d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f8ef20575fb21364c97305f25af64985fa58b24fe385fd4ad3fe02dadfcc22fe9a170d546c73e977192c4cf13ec943c9d50627352c58632d2e69b8a1c903d47546a450efae98b4c81bf714418762924d9e6a27e7b9bf03d5f560abcbee7585e13fef825eda53eb133269a421630e49c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12551cf07535eaacc0b4a5a0cd5590e97c6c9da9e149f2e88be9f3826ff13afbc2acb920c013e3c84b8a0882ab4581b7cd6b99a75737fa6fd2aa19a6fe54bdcdcf67b5f5ad3b8c77da4509c4ed836a01b41fa15ea9db66d87c6323cfd7781643498d24eb241eb0bf9f47c7816e410cf46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2841f064cef637b39652d9ea7a06d18eafff3532f3b27b4c329aee3fc88abb7892d019fe31d569a9737d7de4e96c22c14c3383e2f5d27d9969b3d535a907df70d829192051e6d7f5c4ac217a17da130de40eeae8da2c3758c8dfcd94e6e5a8311edb54bd1f21b886f0020efca5383d8f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e1cf14e50b592f765f05b9c824a5a4ff68877ac4caa2ee18c9b47bce8e96fa6d51181a9bb99dfd523cd8071366f959f561216c921abe346663f38d327f994c180a3867a4499552ad878b355c24aaaf91752c70290968eed3190c6896aa8cfd88ee65f01a78bf69777e189d2070b94577;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37a55a56bf9915b42ac0295c35d9da4eb7713d2b10bdb16c2267b50e93807856142b4f494ac084b4e0b632e5789e7a4d34fcfd82503f6d06e74245c6b729464756acec26a0bccf8377e209f76a9851e9ab72b99046a47b87d488f2286800173803cdbafabbc783c77d5d4b79d202230e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf4bf92151a50189a23d68c8f4c7cc1e72e6cf83bfe7ab0f0a2322f2b9b60534d688a94c4dffd0f0d3dda4ff55c84126f86f86c34181e86dedf9ada9c6d589d3e9d7316a486a0354bae071efe27840d8a7e59883c9be40cdfb86fd7d1305dd781b98c4c13cd986284bc05ad1614b96d25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d6871d9bb2a1199f3ce1feccc480c5eb70867033a634d4cfb16d20ed431f4a19ac9e857f528b42b32ac377dc0c19dc12b1a8f801f9e0d481bb5daa4830afc9d3b200af8087123062b292df42fc448d30b681aabd8ce3433b8a13c7c70284eb8b9db8650d7360ca12640e6662c1d9d5ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71cd7bfe04cf0f38c2ba5d69c85d9242aba6e97e1cfb7e743bd25a12b1588008c392436d67c59f9b5634e674e90f4322894fd1609094685c565690af239ae64eaf4d02be883e7cc5eac466d4b5cf4a72f8d81071b62299cf453531db4a4977b14891cbf2ccdcdb34f474fd89fded3cce9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c717a1817ecdd83bb69ee68e41edd4b65451faeb63e6b463e2a91ef6cba03ee1b7dbcc000051274bc3e07718b62fb8a33f61cf75523a06dc6a1b0541fd654ba0785d8784c1653290f7a13abd7767dbff10879ee6f29d1aae85c34cdc4036fd152152107ce422a0f1fddaaf5624304b85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb345002761b018c308aaa85045f7103f2078eeb030e9e47ae01a92178cd7653993fa569e1143021904d32f8e61e2a98475a2d128c04de085ca43186de6248272e05bfc7666211a2d10e5e38146500997e29850137eeb7a7db5d038b5489b53e720166e0a8384ad03dedb91279c64617f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba7090de2fbece2a3091edf744ad69016414ecebb0c9bbae81004f7d1b7691c677502cf17e3d656cc4f1265114a1a2c8a451ef0b73e4afb101088a9dcc41e36b7124a439f2ed2771694fb9d2f66808bfcdbe6f7746cf8944c67a913783695ca336df77b66049e352fe56a2de8af235019;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cf5cac46d14378183c22caaab466fb6bcac03ccd33f7f9c44d363e2fb9546a65af3ebbf0b1608b3b4cf61723af2cc8ed2c2c6cae7b054f0900bf86a3d5fe093c12ec35f23ff0c75d4f58d71deb6e299feb7b0c3ceb50375d56347be4257306498ae2796abdbd77b8d94c7cd9fc8ef553;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe2ebd7f2fd2553c7aa4fc1c61773662146f51d492da1fe47c7a0b8e1985246c244128456d995b3d4e0a8ecbaf66147f1c2ff5dab467d03df7134a17a630cb4c72e718cb6329e08d5ad2f45a26d2e3a65bfbbf127c238828d86800d6818e649c72cfd9ec84e7a79df5e68c766d5e8a186;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72a15a905598053c93af30cc5011946f3d3f3fd91b954449e8506cd64d7fbe081b7536c1a5b00fdab0fd18d8050b17298480ceeaad674d035918c90c31fd7140c9df04c050a54b52c5de8e76bbdc9cabfe845b267cc0ed3d0df668fdba9ff8b2247dbdbdab7ecc58154c210b92a50cf14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d987f40c85a86917fb2d4d91519094cb6e52497bcda7a3d3c068f69d455705c9fe0bdda085bd696af41c0605b03e2e83ac00ae30732a7f1a18cfb8cbf52fc272b4d0847c5ba8606e16032174a4164d2404e3c2265fa086c5d1c35969507fbb342ef789dbe11efd0c2ed0eb01a6177a1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a99e637335f91e1c606c5311b5615332adf737c92965425bf3cc021cca940b114eb05fe8a23d65faba3e56122eb9fbdc1c136da68d2f8311213ef81d813cd0e9f0c8bf9e4b4ee206ff33176129623da7c625d93c10bf3d56ffa5b28f39a911f9f0b04486eeba7a38ca9db1dab8a7b56d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f09c2bb9be48f85dc7ea353b0c7e977b7b923fbca658d274432257dda499406da299646d07c4c4db10f67aa7c030d5f2f03bbb5f465d16298c61555b94ec6cf1a2bee99b8059c2499a1d1dea9cb546610e01c4abf6b2727795987528e62e6b25ae3862cbda81e7f464f46b776b1ff312;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacbb913e182924278c430c7b4d2288f7a14df7bf99df0c963599256afbdd82bfd10a85cdc967e473d96e4f603e55f46ec0878262ac7e15a445c30a748766092724c92a6fe3d3a62747503c74faeee5095ab19813862b4f814b0afbe7bca12aa4000ebee0c70a6b0142e95dfc6fb2a23ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9b190908f75c811289389d3acc964b237ce6874e7cfa7ebe4a18df032f7d9f394c3e3a7877535a2b2d1da73c3a84315222a5e84785080d04cd1fb0351db1db1cb5916df427da450c89477ac4e334835bf568db405699f2e146d4b5eb2c372f722fadae9e73bb8d51d87c724af3aef244;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha626feb7ce30a0638f10f1105ffce297922c13fd3854d30ee0ca5543e9cfbf72678e69f6baf41007a207e23bcb4e6ac41870b7db72b3d2b8549e7b522024d7b6acac5c9e0e9b630f3d50ae75aa7e8065afdbba847dca28de7dd04fbe9d5f5a70e4c43879c2f9d794d5305bf6fdd2dd067;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7626d3ab158b423ef02f8f3859450164cf8d0632a34fb14054b39f8342cb09d65eefa57befedd418d0c74bd4e021363d3e4460b906f7051f8652efa71c492bf2610f7d1a158457d30ec9c377bf8d40492c972543632962647e37631dbe75ecf3836fe59ab4828a44dd391e12ce5b76db4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h668c94657d301a3d3ff33c6a8ac745baf681e3d23afa6b37722135011b3cfb65939147d22911777f31098a9fcceca80c12213b36157ca93d03b0ea09d962c148cd262e287758a3c5813b00e7a9eda030e965a990e23d0c6e674b8d07e9b87ac744ccf7c3079dc17770ffc651d76e11894;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h763f5a9d40c0a26e16fcf29d54df164ffd33e9534f91892a275dfdc5a95b29550ae389f0a4b665b945bf874c137a421c03c8bdb254ac6e6366fdaa95aa51d32d438c1da76cc51bedaf881012a1c5658cc2ad8a347e3f91d2fcb20c892b49949f25ba6eb7510860254edddd6cef3794e4c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6638b5372bdb0aaad9114cb80510d189ba7de138322f72916f487f025757f280e92cde97a1ba06401f5bc95be6b731289ffb56dc2b7174a9f9dc33cfd5e00b8b609643049bf2faa13f41b207feed5603432c204fee3dbdef808a1b81d2d1ea4a4f0f3ecddd8acf4bc99663e2b7bfae0a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he01f5438fecb1e78040c6cb234c972d9c5b01730083e7e6371f28ec07d12b77c9c6316fda96b70d32b5016c5fd1b6cdf9c32b8b3875dcc2155a7567e74e8729c3a3d7c7732b9222e7a6bc7abc74ea5d9d57feb530a013b2f7e6d5ee131a962b884d864c97d04a44407803820d6511d0e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bba177de7ee5856565be7b296d8bd1459c75a50e9179c96dc7a7756df68e3a076ca02ff5578a22e046fe057effc11226dd5a094c63826ce450b92a335af9cc64c9e33bbba0a3a7d56dc1ff4e1ce3acbdcd4a98f5c8d7b8fb5e5debc90adcdf8c633e2f1d57b5a9bdac7c4aeef2f596e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9ccdb60621c68a9e30a8c945fbd4f4042d4fce8d610ad7514693aae412f21d24c75a0b1e393b372adb94baae4f34db5a422be397b57b17d2e2459b00d86596fc5611bf89edd96dbeac4be4a76b495172dcb437be1a9867739794ab91704def144e07b27b7a892a7293e11fe5869ce26f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d9f728cea9b451abff50e7e0b157d8c0181f9cb494701feef8939400f2faf3a14ee960bb6973702e97a1da65d367d0f5f667d60eda7604056011ec8e2de64f86e687b398288b669ca9abf5c21f0bfbf22ac1d5774317e9e1d5561c6d7c4200cf016634640d2b3f2161a4a2d3a30cdb1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb188608780cf4642f384b6ccb8dac43de49c81a3041cb81d4dc68650c0df844781d61032e7fd263244caf40b99051e357ee991cdd25e677e4f204d2bf98082d5ef86e7d728e02fd307ae66a3d085ff86f39aaeb9b379ef580d4c71fba50185895b13b7149b297db040806f0a930b56d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a6070fd07ffe35f606be3a48b1d98660275d9dad457784e6e95d39915407ecee63ac45f638853bca17c2a2503f95148476b887eb675431482c759ad4f6ec0d7483b2dc1d8ed99fb9ff886a1e75aa78d9a0f975626cda225087b079dda8f2dff90e3cb1db3474a3e7c7864832fafb08b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a48d5bc579ab2bdaf4822ce7ce087cb4619506dda4556d9e693e3349bf90f304ae9b4c9f41dee4eeb088e744554a489deedc56b4ed33be2f93dabef2327c7c7e5714c11135635258bf8d8c01443ce1308cf12971f7f2b061a208f2bb331b8a40ac1aec5952b6fe8c2582537db7195e99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a619debe1155f2ba7ad65c5d19a9fa901ea119c43007eb52a1f47f7e7d374e912b3a42a248da12ef344b64419c597054c7c02ada7cd8567839051cdacafaaa14bd021e202ff93a34c63947ac539129e6a57efa7994163bf3fb93f9c5b2d027480533bde208ce886f7ae04ea8efd9e76a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c9f20f874e20f00e5fe820079826675c68d868ad943a03f6a4ebf03898e2a926bec749c2744efd169e0467c0348b221993c9fc87cc7afbc1433a7d900ace69af3cbc4769ed7e4e05edcb718c2f2b2815b4ab59c15154ab666a191459bd180cb5ad2a7222c72957668ef8d020e8e87f34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb648ef90aa0b98382b085dfb0a1756a6c701eb20b8922b780a2a5c5eae31a2b86350a13f7ef86d61e74fa507cf62c626374e822e4025c6e4724af1b2ff7702750dc8e56d92d41a19a349e5d9c64e8575a1e58bdbce10ed98ba0e3fc9a0e0d53e31bcbaf3312f2911ce53e445d112df57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95505e31c64832001a96809cd7ad66ec22e317753a619257d72f6b42fcc90d4dc20097a33bbef971ed8193d8b2e04b9d46a6adeb9d6f6fcfaa0cbd0a6263e86cfcbd8ce70b747b2f39016c64e6aa294bc0e66e56c2455d84262983c177090d80690124ae9fdf479b56e5c387e3f7c9f94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99a141431d2c576058a4385ca270f0230339132f2d7911879689b33950fa5f4a16321e2a8eb9aa3bf30cde3be3cb89ea14dfaf7b7215a97f112351a2e18143f0b6bdf62f7acec6af8e5d196a1d8204c47be141164f3bc8219418493487ec92a9443cfb4ee855df410154a6f8c9e217f45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a2fccf4b805be3111d78a4f4664dd85eb574816f3111404d066ddaefe58bea7ea224d5ed773fd99fc42968bc09fc6e34fca864568f72b0da1b88853e2e41839b0d35891d111f5aace2ca4b5116512acd92261a7a197db730e105e836aa6a025dfc8821a451902393decda85e2c8c705a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdc9507239f9b7ca14cd5f4a575763691f3f6e3570f680b864c81c43a77b1d70a03aa7faa9e287dc754e34dcd7dada24dcd12e59a5e8652bead076a89e8a067149da43abf19b5734ef36b2a0875538dd4815248d01d80bc813c8a18ecbf7e3b2d63052cedc47b4226a9e4992767a46645;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d61b00d21ef99553107100abf0eddf3a0795622dddfe61de82998a2615c67307c6b4bb259ee76880ca5908e85220cc5eab16b9ff3b54ef363700108f7f66e5752b14560e2f294dbbefef7aa6aa47b36d602ae516dd16ee31bac2d1e810743abededc036cef2d6ff967f574d840850de3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h116b726ad7c74853b568c813b5efcad7afc67d7e4d4df895ae88fe1d6729f5f1188c7d37f08d756d3f4b179496c88703796fb4994e70112a61ac78aca914d6559d0c35817221c4aa24f598011114bd26a71b391501bbeac4eba623ab88498d6e1a5bde8828e75cf649111c2a64debbeee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb466be12c8a0b44360ccc76e9e00b49c36fb49626209217e1d14b0ab5ab7830c52f141d6fc51acb54ddbc93c715365c94c561d1c3c55eb7211fb3f705f7dade8c246828f0d5abebc0f9e2312f1c1818f60d156f68f14db8fbe26383af38799a158ccc739a5b4fef621eac9aba63f29ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14967e283fc6a90ed8fd59c150635596966d1c24dbe805c32a5ff5a5a9630f165ca9204e964afe45b33abd96c762af59060a00eb373a29430991b921d52fc0e77c86b4a36f95c7b7ed787f05d3c80a62c4b96b5ec6a2bab5da7235ee429c4935a00d5c1f7a9c787dc6d135bf8c2d62348;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c26b0fd8756f2bf7b4bf7af6d24e83df7670d4aeb3851c5118f6897bf52e4a7bc208a3aed38c7893d2cc43402a4c7007bf0aa03657c8cbe6093d40b029ff8f6d9cfff54caebf14675d626a5de9010155cef607aca340c0c0205085bc782c29b6f2e0fadb3fa44361fb29b39e068b116c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had01d607289a82ea3108c7fa89b97be3297255b399e62c322cda74ea047abcdfe01d0b0100d60e5949e216bc63eb3605ea8015ebb1a397008f1674e273bdce151f198e7234387c0c22f639d9bc30a677c9076de17f7668a0cee394427d37a69b464c05de00042d7ac5f489a9292f69220;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h927850272b34c217117ff01911cbec932fccf52ab0dbfdbe04a1a3226ed37caccdec446030c6dd8006d340e30a7691ad640995f684d369d3047cda370ac65e7848e85466760f76b6cdda5674de3cd98aa9ed70b250d340fb90322239692443a5710e21de71d077ad8d9a72bb975b0f9ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h942fc91702a7dac7ed32195ec538fb3fba7e1a37155617f99260848b97208da2c7e8e0eaf1ebe6e5ddf340e77131adc89b0f1d8c8a18a5e7abb714cfcd35e5cea602bf685bc313049028e2f487219d84fbe9a4c614863faf6f9eb44ae6cefe9997b61d233676c0782004e832294800f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1db7a033c9ac19c684d7f85b6665ba88c841785cab0443944bcf1c0aa07f9010b6a7b737eef7813021b04eeb29743c72d9ea6acb0f6051a59eaee9d459d47f3cd5fce3a2e0916cc1debb23447b5b9c16e4315c40d41af3178e15e6fad5bede650f2a096e9d140effde7cafdf6f7c7fed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6032650aebca11a336b71c7359dbbd80b97ca9048f79d044135c19ca7319ce108f4891c4c26542cb8fb782044e94a37afd0451173e9edcec899294ebe592dfe52111903976a2807def75a5e750e82acedfe850c17e1fc55506ca48dde28437727dce2b94a4d9a20053fe48adc3fa218c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he10561867a5dfe239eb0a5c793ebdec114d0d13e28053cf76a2542956e295dc5060c0b212fd14acf26eb86b2da9196e5f20cb4a20ff8cf06b73afee356c265e4dbf74bf28c857b3a2f2f9c0f3a944d7ee9ab35bd0fbe83ce9fdfd7464d8e2d46198a3fb64bfc31873adcf625810ba3cd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66f6d88d855b227c948614c4b023acf6ebf40336ad2cf93ac7817a12657100f3c849b72dd904959d6ab3e43d818a3c43c929f5691145b4263f3d7c9cc8c3faff15167fb369dfffff9a8a115fa35636dc7b3d6f14659b1dca75064bbbbd37dde12b4da9109ab11b76ee31e766956f1bd44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dc4cb3fb0c2e1e5427abf512c00c7cb9f3b7a14651279d69d883f827af2ee4f50e97c240dff807f3d42348f42333148a1d4d052179f4ab6b51cf8426d64722ed2c689b2532889278aa614de7691bcf08a6ff22b13d4f1a8a9ad3faef3bb77b322d4b5da1521d1f48ebec85a4b4288a1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13362eccaf5bb9c2c41b82ed30287943e1b246611aa0dca18c0212b70c33c1523ac480909bf59ae373c085d1136d31fd1e16832408e5e3664eb4bd80e56ccd99a9af71581eb32aad171336711da2fb95aed4efd5b8c90b76778f3cf06020a2fa12ba5d3d3f15a2891c7316ef226691c82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h826f773d6c9b62f6a783548d6a9968dedcdaae2d9a768b75d25fdd43e321bccb970d79b509ebf4458c9079686fd2bceff5cd7519be0d6014c5cd7ad88cf185a7ae0709f42f0ec70b7a60cdedbec99acf62bd42547ef4246f6ab830cba3e673cbff2dcb5fd04efa882e965224f3a53f1a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17f1d9c02062584e34d45e7081a10a0aedbc3a9dd32b924278a53942e5fc670fdf61a75b6665e6f5824dc4eac9ca9539a25e37b03cce2ec953793aca7b622bf15b13d93d7f03142f92b32e31de68cce1ad54170b11029cf411a6378fbb4f964d73d6a71a802dc161fcab9dadc00dfa0db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h543e0b42c11ee11a910965a5a789439de1fbbb990f8eed135772b34a170ba51dd09836cd161eca8a7a252c7e42109538e16df0f2729b78d08ac433496d436e13151b98fd48ef09c914650b1af437046267549909170b6b42d1869be89fbb7ad7f66df4a60bde7cbf2c473978801b0f34e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h695f54ec47b43e593b2cbc14773607ea7894c0dc0d03d7be0a810c04450d76c46d00c147b17834293e01f639d6c8eeaa1413157b1beafb0808ddd4850b7e3763236e58fa741725da599a5e4973f531540d29d6c865d4c76fa2b4d15bf52b73c1c21e178fe4bc32c616450982365faf140;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c9cf874583d1d62dece77e2281d0e007907ae1c6d85da44c112c03fcd384908f15892191a2f847d24d5fe64dbfabe567fc09deaad9e22394fd8ed6eb99dd2808f26d5de2f906686d775101848d6769a493c77b852e846cb191faf4766cba09917d3237e3d572a9f124a17982ea9c2790;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heac8e8f0f2b2242604051e903f4413005004e23a8c45e6099770f0b163d4c689fd1c6a9c120fb94007f95b3008a843c873a9763e07c9e1633959dc8940bc90f74cb5bd3714f361bc34c49359bff9e72cede82e853b4893d2d45526ca40dbd010a6f0996b986845f58f5aea4477b198c07;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc812c21c865e51c8440e9f5efda8d8e27c78516f72fdf694e294e733c35fa7eb68954dcf02d6dbd44718c72da13764a3720bea19b42ee6fee401319423f0ae7bc6d09c8df3595676195100b21115cce434284ab3a3c3c48f16e15b47e02fa8fc854b1447e3a02d55d4f17182996642f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd22cb29b0bc0cbadec34d031a0eb35a0663d0e4cdfadb88ef59666cef3399c19016e4573d0537a6e8e12f0672ab5476736250cb1fac4db79c0ec0404f14744a23b64723209d47591219ab543e90f63102f3b48bba43da382ecb9898c09731496194568c03a883faaa12b622039a50f6b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f219f0a61dddede4d8c515573d178a7a6d239eb1ee6c88ce3a5a1572b3c073f4a8d3fa9fdd9e52de978f27217a5743e169cfaaa78e3a37c4825696f2eb61b5b65663a47a6b5239007a8a01938b089816e97b6df84fcfb44967f1b086df8b9200bf8a5c595f798b54ce411e6a3a879659;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h780c91628cc7ce39bcff6b24f8113664b759fb878bcf693a9190fbeb36e1e5f786146d37eabcc664cee66d35318b894239affac28befdd68e5e4545889009dc15eebdd101762acf77390600a32de6d4837abb1d561a81e7d3a5b080aa98f0cdcb9c2d90daa3241d7eda426b6620837c93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb4c698d3f958a327af3c7872698a746e78cae92a35906e2a949d89a130eda0ffeb68e09e277be50f2449749240274b9901e68114c15c83471e8badbfaac25d9b3d0ac38df06f0dd7a5a82d109120fdf9baa27ca23651a4589c61f307522127a35c2e9253c2f7af8420335401321b53f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf3e695bc08e917518f852c2260e1fee1f0b38a119a2ae85bce22858a842a72beaae572550336dfe62bbe729c4c9791662b8019595994739542caae1175487ac2da162d48867ebeac9a62f4a631a2ba6f332c2e3d013a04cf21370b272d410988c55613cb97fea3d0d1a54b99bc5962a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7765e309879c69f2e79e264da357255a236d297fbf62fe1303fcf979bc9bad68507d46f3681904a9ee9e2e5f080425b3018da6b4090a588beba2d1653ba15c96fc5f0d209da1281118f6f4fa045f93697996df881620ffc35f252c8bf9589b9523aa5e055c31830919cf14539f7b0473;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he016ac162fa18aab2e12d07d0b3a0280f262a1f6db9b3760e273c7e1f9882ab5b377386a57d94c5d093a686a1a599d3226a370a765b03b35872cfc2b82e4c62aaa383db99249f344aa072f12d35ede862451e9628e20d5a314d0b6baed6fb786a427e8b37aff1daa9511fe901e31cdb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2176bbb883e59f7b13cb9f27e73c7a01c0a276dd35fbff169e2952024d3fef0df90af20098ea75cfab185e7ce591ecf6eda5a9663edfb762e4a55a691d8ea824214a64723f492a3d20909dfa2f2d02b1d933728985fd244c807afd0a7b9310fc337f581287e83c5c60d3d3ecfd835cd5a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff198355819e597f2c2721e38ff33d0b510892a3a9047ecf0421c09a6473defaf832f9871b7a097a1fb01c44d3cda38b8f6b0bc33976a860188da91ea87a43b03272c2c32d66aa608097afe73af26962279465f7d2245282b1d5b99ea12406ebb67c3ad2f0a3d7b3d8afe5795692fba55;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9829f22b310162d5303923992fecec1ee9e1c27e91e71982c53773d9100e11a216f25aacedc0c7cdf0e1eb11a86ddf552adfdbd57f06012a84098c9e2dcd7ddcdc35406f6c971ecde414839ceab78510ae9cef1d30ee1b1f36dfb83ba8acd335d491da2b65546312c917ae635cf12085;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7771c29e14bc8889dc506e85b3b7e91808cd7f8aa8e23b432b95ed34e3db40bd573b4e5a930b966040c7163e2410f810218d1e4b3bfc354844f702b12ace5e04c09bb9e4e923e7916bf74e65ac8942e59f70099944db473343beffc74c03845e69522cf9dfd320a5d911813f01ac2fd1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb71ad35f40431a7037e2c61f1c3bcc38cf17a6a44502bf97b28da29121601879204d5dc73c7d0ab9e255d0c4e03abc7d51e79b527de070fd6ed8d7fbcaec6f7f1c493c31ef5b72ad60c15aab479235148eb261b70392d3cb001d8f8d8ae2626cf1374ca21c2167db9ca27320797cbb1f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc051061b45dd993a970d82877042083243c7664db8362e7517abc39260c07021d7258a3a60ab7f6b2075a2fd7c5098f5ac78e3c72866f68218a8d43db707852f01b372d2b7255f640baa242e2fff65c24696f0162dc7d9b02f12e71d4a8142f5380c571d02ec0d02629b623fc36edf11b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61b609c8f7626a35d3e7b5e39e0412552e440115561eaaf52d6e07a4d156be396742150c02d4709d09adb42d0baecf2e65e1250fb15eeae93aede3d626375f03983d74acca8604bcaf144d5428af8f2236de88213f53729848e7eb9ddf527366b87ba811a9a834c484f39847dde114bed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d31edabd9a399f9430a5ef882da3190087dacb196024b182b77f62087b735bae0f5ae76062089c0ea5040d244363a41ad2d27eb5c28a6e73065aae7b04ea4ee7f09cb25a185e98f7f1d853af8520079186b553ee18821462cc4d1b17a1ca58ddffba5b713348bcc70edf8c43c8680a3f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd83f2fa5ab42ced9d7f91d4d6ba8f8b46fee0402b9009b1235750b88eb17468b34f7d5e3c42a15f7281d9f15316ee54a78e9dadfd28149345ccf8da6bd40f9f7fc5b1b56deeddb99b98d7891a07dd42af34ad23e330ee94a6854438522d123c2725dcfc5b85259c9d99631ed3a4d7bd2e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6550cb744bc41c1df35f62ac23b613b5f4af403c76625e89503ece3212727f3ebb9a447c6940c539d38034b683a5503761aa78b2e713a233ac9813bf536b49d526d3a5b06fcfb278b9e2c1072744099051b1670ca8fa6426169e923303674956b4eaae25399f6c3fbbf88fb564796ac12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8058d11e7831e0c2c058515b81eb58721ed9d8c64a98780438dcce60dbf6802ed5533cb91b83a2630e8006aac3e4a1439a2350ebb7e5bed07e2ca2d9f9e5ae1cf4eba95178b9aeb60357403e5d0353ad221f8e28cd693a45b1237fff85b3dbce2865a64b7e4720246b6553224aa17ab62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19df5c9717c0ce2c404c54036bae88d7d139c605ff35a46c247c8e7de7012582d70630eb8433de217fce9a6c445e60e9309bbeb32caa4b3d606ea771c6f6980023ab36544f588ee77a330ddf5b21dabc451eaa5836a0fafda67860ffa0f7991c681e0aef524ab63ecae7877cfe136658;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd22e46e493f9362b45092da47f01b98e410e9e9d6fcccc623db7a36810d55ef08472f961142c921ebfd626c1c65376855884b900d22cd492feb1b74481c3733f03eb90c89848a439d59a00b4963e13d81662e8080219b79c56c38aca60bdbc4f9936f8f537dbf40cce66b21f5b461cc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2548f235426b3e3b03e019f60149e6b2dc1f5adb75c965d5dd3d3d3f464e43e5d6c59e7f26233260b5d157d5ab5a44fb85d79ac79727491496fa456f6a6c857e4254c17f51d2ba800cd64c434388a83865416287199ddfad7eff9ef45519284d58bed4e3252c9253cc2a50d321dffd34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc6909c435e7fde1769c2b1a04c8ffd216870c9960072af8f13af73718b39cbb282b8b0ba0bddaa8289f92a0fd7d5b77d9a88e4b750866c07d66b8c0c5a8281ce3c316327180f8f476b427d8f94e0d9bf3e1f5c4d5d2fa96ee768be9e6823b40814596762a74ada9ddf4d62a4bb59e367;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89c2a14043d97ad51fa09128122b53ae772ffd098967a4e4a558ae4ac6f87a7892cf7342dae77a25543d1ef846acd82355df3e2696d24c4095e5b2a6ff8cad1bf404724e9fd2b71f44a155fae1f9ae05771f7ae593c642e0840228022bd4ee9217df7353a95426d653ca6a35c84f1595d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h916ada2eccf9bef6a735a5c8ef22ca24a4f10ed84a1896a40863e1c1c588eb026df4fffb5c76ae7b516adaf4cb8394a0fb1f0daa8252ec9c72b5e1ae42d955bfba603b0e788646e58aec4dadfc71874f0ff20c62e4ba0744afd70fa021edf0d3b9e4738fbc4c2a858634c9117fb78cb0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88705b6b6196e2926897ef46222fde3b287f95a98c71191afe516b961b1d3758d0a090941be9b353897a9504785a761b0cfe1fa4e9af70ec0c9e555bdfc24d83607596725d54399e820e8e162920bef2527c2797e361f11cd040986660b17574af383fc62b907a890e81948180dacbc43;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha48d3fa46a7f53b13485b9c40a2e53d5da3f4fa977b090c2360778d3d6ef63f46be147cb6b9256692284f06c91ef3531f4f81ed724aced8047516d9fa3c160fa9e5292e6e84a1013bb3b4bbea90026f1af72f7d5e96e881e1cbbe5dfe19e3cd8cb912dde57649c0ec52b94d2a10408ca1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc75dba9bb0820d7481d801a894074fc9003e61616d19afb3145147904dfb60c2ea60c9c322f3c84297e4eef0e0c925347f59c527880f44a7053f742a780df9722f81ac0e6fce32c8167304299e5337a4682ded0432dfcacbfb6fdc4c33f6b07c0b8ed33d52ef654e69afb0e906918e886;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h812c93844962f7b3d4797722b50f0c2c1249a01e926c69eb28e06955f8ab41aa576ff89f9d21cd0b56937752c36bf664804dffc3c2bacd3343d848e302f56146f8a8104f121212fc43080e6872bb325519886242a108838b688f5a89a6b0551b5f94d6557acbdd03980c22b0d26d75967;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h368439117ca0de4b085cb5ac50291551342d9c8792cf5e1b669140f29c2ba82baf8d8a0e42d943ec88c9dd362dc96953b3e0119d41a2fc445de3ec02317d525f664f62a383abd9b9a6a275dfebe38fedd81825f3f2e549ed0ccf5d24312f6edf3a19206f4f5c8b831596312991c2d46;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d905423398137b5d7a5cc789d52a683bd3bc77ea88247361c46c7d535f2cd6a85c22e46515c1c8d62771654cc3060dab8514bc7065c2f8058e8ec33c25ebf8fd98d43bf79defa6cf0b06f77982e4e1154028e5519fdedf17b8b46d4b18d3738d74a73b7ed44e60a0eb31639bc9a4c1d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1c4610b88b3a8d992ed667308ef0c7edc1a395d503f2ae8e273e04af5a723a6df4ead06f06288703cf27f97538ee0348062e7d68de4e5850d532f9073c0776de3349dd35843d46a06b0a93f97484e9c3970483f10ff3a362720bcb8fe011e410e0785e112e257245c862703b6700f6eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cb70b2bb9a8cca55823a068c525fea3b54d7ab2cbee491baa3cff9e0999a85e0833d9e778331932e9c8e84446bb2591be08d4def8a2d12bd83fdde29e9c88c0aa7d6ef73e52cc02c45a74f46b68e7675bab22203a98fa6b3047deb56db0c03c87598816cbb3de3e37f19977a395691ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h523ecc06c39a39a78b4406312ebe143618bb7ac9de18ab15d1661584c68d07e46fa947a493e6f7bd594940030042671fe6e317642cabaaeb195b0e9961d28a46110db72c26452070de8dd666b887177e00be3f94abb60321b8402693f16b3d2e800a4c8b8e3a9ae33b03ef1f4dfa076d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h704d7c0ea319b3d45ebe9b05be53936f949c97175bcab1c786502d1f896991e50f8bf91325ef71dd65928b797c6defb5902090eb3dc110ce7ca6b24d2f0116906d9f2f7d8df9917aa87058bf9b33e1e4bf568ae0dc258140e1d2a6304d4f804dec975e298fa55fd57f82457572d5c130a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h376fdd2f6dd61b022fe554b1a8178a4dd1c73f6902b583982a8b960ec3e8ace59615b373b12b72dd8abe2f932b3bf377969cec5931cfe8918a67c868c74d42d473ccf2f7a357dd61595ecaf57e58c27d7bb0ee8a2b50322af8616cb1fe9fef48f3f315e075cb50860523bb11c7d491cde;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h884d71442b1b9d3a2eaa9f264642f082528fd755af5971cbf4ae791cd98886f4c2048b29c0dab0c3115fbeb49225aed100833a900dcddf4a36197a3541a11778bcf136c0c0336c45b9cdfe25c552d881cc9d7cd96838f31c7a8db2c06fc784ece5c30ec4269ecd70a9f57c99fde6544dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77ed24d63d0c4a23b07752162a9bc428758a385e39b7824e49f4e5fb1bd4a053efd725f19ab9ffcb81be907579dc6164db221683f86dc9d585de5b6338685dcf7f12cbff5004067c95554809f29ae129641e1e41d70be831c6fb1a86c291d9d4e188adb5b7eaadbbb61a056165d6cf791;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d37d501976965414dffbf415f7a697828ea80dd8a754dfa6125c7c2d1cee1b2a7ec936a6ede328111232fa83e181710339d435ac008725d0165c4c6c9b988ecad237dfd958d3e26dfd26268cfed7740b44332c82ff5da3f86a22bdbdf441acb669f660d38a633a7af8b3c5a10c1ce960;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87b42a0755343a4659865d4f2ff6245e2d73d49d079fa70a3115e4c6efc657912142a7e3f67cd68308dad9dc439a63465ff18053b39649c9b726ff5b12bb43f60c8c545b337d06eeaed38565890f15473d52a34e6e8f637b91b0abfaa93855a75a39f5ac878930ace0ed04a2e146eff83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf93188c30ae1983dd792ffb1d30064111133ec5e9b3a41048985e02ff4d5b4aa1c32c59d6a5bf75dff28e6edbaba31acc905fb4122f8e84f55c3ca706b3bf11e6c74c0a3f68c5f56cb9d812b425e6cac8a4c22692325594d09f4006e739bb95b50adabc71ab760d8c3220c8ff62237789;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2dfa3bcf369885f7cb3b5ab96d5b94acf162b7a9a1cf7ce07ffd8389b14af3dba9832b6cc6e7ae01fce5814bc81277dfcb24825e28990cb93854594b3a69b923febf99ebdf562847be33753a1950e44aea5cf17685358c3806019baceb200024d2f492e6295850cd757588e8b5bec08ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9db7bc813f0cc2cb54525c07d653f63bdde3d02865628408ef308fa015faa1abdb4119c498e7e86e08554d791fc4df6db645d0e67a1ac46b997720dca3dce1a082355a2eeee3de48753869eca82875acb18c87673c5436ed6066763bd797d97ed40a2ea06596bcead412a50a20e290454;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38c44c72b760dd6ceeee079b5fa03af847b7f94c60457684ed7ebc15fcabfdee5edac488ea6d5ef088529fad67b8e89f67333bdb34eaf0581a6334b8ab26cebc7f6a74c5e70c5354df55fac8afb25f9e6d02bab0ffecec478fb5bb8c2b1b8b2249ba6229e0003fc9635d27ccbf5f29abb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haacb027a679b047095018119b67c9088e0b62947ee9a17f956ad08e84113fd755ed4a55e51b72a70af6902d6e583ca3863c81e2b1b002a93a3a406124b7271e3af3dec2db4f25a44da2405f0a6fdea58fa58d3d35cbcc07bc26661d34b02cdef680979d7a7b02b3e137bbb0100c3be55e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2365e93ad5d136c6f9867311c71465f0b282cea0b5b56d147dddbc7b57646406216e1ee5cd869cb7bfc75d7c56629bff405fca55decaab493f0f748605f798eaddfdc34d2de7dcae5fdc1c251e6451be5cae7d161f4ea45fd643b85300275cd077934199631e908b58332a282e3b0a37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb79894d1c69eb9369cba3ccdb823c62feec1d6ecf1062e7f0ee5da38453cb4c8772242e2e98605a2ccd8d6f92f5b2ac66a95d4b1d27344cca5900a46cb1ea907dc7ea2f9a2f0faaa8e872fcb1bf348b758e80621bc34d872cd4c19967a3b4c2fda06a9c8ec278a6ade8a27e39ae16e561;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97a1523c2f69e5ac86278d9777408f98fd01d7720fd8ae3f58e7cbd201bd8dcbc69f231430ad3b98ce6c89493b24914b770fc726869844bea543d4601e2d0af9e96c9e2870e37610c0788514476e080d1c1f16bf7537e79a81cdcd4d5180a39aee59a3bc8bfc7861dbc814540897afb45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb006be0def19b57a8dfb5fdc6d172c3df4e05f1cc687b0d81b2c97c5fbbd03d61e1303c5c07898b115cd047a5f1ca58327970810fa34a3e82ae09d18326c031b737666cc7ea173c4e1a988464d5f5036e2136c9b03dc464f5ef4a0c837cd0c8eb898722bd3c04c0fdd4813d2df14f725;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67fa34ef309a1809c018e88caf8792b3c5b24c7a3795eb7ad071d442a145b2d16a3c4bb938b75d32056363bdc96d525db01bade1b70d3e697075e8d3056db9f7278b992ad4e6a3332db77c8e93828dec2b2b8c17156b492ee84626c01884ddd4eea714cd55e73c0af39cb8eda2ab21841;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39e6d2e79eb720b309270dc323cf0523eb752be86eec5a0de3e84eaa7fdc6a1cde830f5ab9fa20fa39224ce8a2586fa717aac87dbf55bf6de14127829d82a04747b13171dc67bd8371b531c8a31a2f74b96033a08bfda7ab07ee33af2cb6fa2640e90cf2d42619342743f661322362102;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c67ca87fd6c24b1bcb14cc848a238555008c6ca35bb3bc56467084ccec2586c8e585238b2d8366cf49ee9c41383bbdf9d5c33f7e06336ea8b6d5dbad8d041099b53a016983ef50c6d718856ff93046238b6bd5319aa2091737dfe67d45aa1fcde3155ded27540acf60fb9e8897c89119;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd15ca7fe100b7219e9dba38ede4bf2e58e24f94a90d924d0cb5015b1499e1ead52507a0a33664f90283ed028d1809ffa9ff960e5fe0414644e97a83fe2ab5ca5ae3db1daa769080b0fd00814583acd49649edb908026769a7c8ae2faea87e695402a1d7044c1e976ce175bbbbd9e281c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ec55db0d383b2d774242ef51513675ebfe537e2eb52c99eb5325cf390c2f7069e5b80c1e15f8dc13cc1baa0f1152fd5750415b5e42d4b78f319afa4d581738c71323813cd84e343855ad2915eeb8b650f21eec54b8162ca4e849a79205eb8056fd8153fd920321cc18f4b73b21189208;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h832c0d7f4ae36027a87c910e5876064924fb05ff9a9f640a020153ca1747d49965ae25c9ba8640459c629fe50f903c8a6c05f879cd280e7213331047125e75e6202afb2bc85621451cb5b9e2eda313ae39e2e0a2546c0b6b4c0d3df9dd23bd478355e735e41114785ea13b5738bc040f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h447cfaa96d177094d89db982f59db01dda902fed5e4e622f42d9c8bbf87684a72e50aee79a10a415bd816c10c588fb8a0b620d650ea90dc908cedec1a296e160f28a5f2790bd339aaeb3afb4a37620ee39a4e159128fa62f22ef72f0dfb465b6a9b03e0cd650eb70bf0e1395723fb09c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42c0d383c988339b546a08fa237f22fe3f199380b73045753975e8f31ac7aa3fae544abe0b5c3a208592675d98a22695777d351b3a9dea100c3e6e3c734c86d2ec524ab7d046cae8ff042d2cd4b4ccb4656014ddac6ee6e3dc5ed322d90bee829ccfa642e9ac89b3b21116656426af9e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1090473a5e6c69b094e17bc926280899d53c35a4d7bc9babae2d27d17ee65b52f492ce42d4b73da9dd8169c87e136a3c0937f3d186b349d52e16ad1e0bc1814f96b4580ecefb5fcc2976df087892bd809624e1d97abc9ec14fb5411a0dc8e2da89930aed6b03d48aaf2ff21bafd688b0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebe9ee12d0a8db68536bd676302a5ab15ce9203df9931994ab19da1dc48f7c0d986a1534d9472ee4a0fb55dffdaeb368197acf6dfc11fd25d0d6b1b39bfeb943c586e7cde303de7e4b4d8f870ab1ac755865698414794f12fa97370760d4326c4f3b6f96578db35fac5b00bbfb4963bc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e850915e35aedb473955df51eab4f486dbd7ce5ae722d30706d844a5516a850cebbd3e0a9062dd8b3b434a04acc9a06b08e6b89dbb59315e885bf7db8677ad6e7b33ca2d4160b1e29ccbdf43e03ef62b3345d20f4355c87e81f2f24d42fb5375708b542be6c88a717a4e210e4743c524;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd115364ba1765a4065f9d4e85b98f0568e6c2c27c1faddc30f33e672dff16fb637683a170d57f15f260fc14747bf92628f7e0c2db94ced798dd3c98eebb3f69d9fcb91626fc7e7576b1fcd93d98810e769e056173b3d9bd85a592568fe2c5298f262a94ee6bdb804ae820963c70011450;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h390f32d9280cfdde20166e208959724991eb72b75caebbadbe8ce7ffd96430936e4e80619ab22b95342254b524c80857e2d9e59c5b793c3be74d2289d5591fdee222e6309b4935a4cb561ee526687028b026e05ab1f1d56c4f5c53daba0fc8966aaac32f6abed3d056623b04ca2b7ebb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb59185028be2ca08b72159eb267c48067680e5141d0d8d7f45a4b5b1e724596582ea8d7fdf26c26612f18e3fe16d2a55d8e237c2be66b675815d142e536efe34bbb3a8d682635f9cbb728349bf954d8868eb13b2d1e7d8530f779add7e9ed5b11c1eb6b8b3bb8a417e04bbf313306af24;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h516ca4c95f50103125283eb3f9209fc19b1dd0ed1a6caabeb70346f31b4c3aae9a5cb41df86ad10a3a4106eeba72bd77b29445b0d27f1eaa15b0b093449fd9741ef4feb47288afdeb8e162c6255a15ee1b949e58f33dfa700bb026a3a8611b5c05433cd84d64b98281cb3344494aca8c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc927cdf1c2c8721acf1539b12281b820d5003064c4b1b067b034aa9a95c8b01edb4475cae8e98c3bb4a9032668c609daba733f7e8d892d609cfd25329fdca5ae3add79899de55a29102bc933dc69e2837b96605b3fca77a30b4a76da20a1bbc4ffe7e3104f1f24e665a89070181810476;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6216e9daec841bac478c6cf17e67f7f0b34ec56dffe965b564ebf6236f9270c370b58bd7265779ed12c54947b6774ce7e9162f38986c9f2cc2f10c3b06fd2b65719725f720bce410b3b01593eeba28c1bba3ee64c82706fa1f923ab1d97883600872c35751ca93f8f25d56f84068ecca8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12a666ef72f303cb1f9358749a129cea899f2e5e5aad030ddcff5ad65380743b4366c04e8e75425025a71615e29946e70eca6b74a719d1bf90af27eda6f7cb7863f9a35ca9aee50f03c11defa6907bf2d2ee31aa6b9ff84d789152e823e8ea87b566d40badc06cbe1fbb073654bcc7589;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26da232b6bfad62164691b79f40127a6ef0e7e56e0aa16d4cb7e5cf1ddb1e2ffa02e0984c4c35ea856aa643aa3f255cc10704edc8d3ec3598cabdaa3b30ce83d395a446f3b482fa5b922994db62c8c87821fe90aa3a1e8191f498ca99278df41cb1a70634b57829b8b167dea3aaa34425;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h646a37ff8d29b29cdd44683151aa1b59f7196897bc7bdb5294d38bbd79f2e02a7a1234f60f4e7c753fc0cdd97211bc06847b0acbe37c5ff3f948199fde0dc5ecee45ad864f2e9f72aa7d5fe67d04145d99611e1f3deac5e858db37c9e05279eff73e6ccccc4e97a6662ae163a73b71abd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h520ed6796089425cca16e9ddb069770bc74e98b0e9b1d6f18fb1b4ddd35472478de0170f09abc970f9d60313019382585337d60da101e7bb7b8995203d215538202476db1bf467593a0d770c655d8841f24ae27f0b8c0c288a7af6c9d45d522d5a358016d507d4135820ec947ce4c5782;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b384f5aef46dc5d6d7148b30f2a08a8cd0b0a9b58d723a1ee5d30fa7ced1091037886793f5b40f7a59eb535775bae274d76262b73ff816410a25bfa246d8c31055e7ef01c37f30ab792a94ca058d2abf1b270c7f9561f2c2a15090c250318bbf526dc1a2fe68d990d8206d6d3233e05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3eef1ac014ae744ece96ce53de566e89aa47713cf6c496f7223e4f97eb4f79e24dce4977ef01a4d62f0069e2df8f7410ded91bd23ee6f341493a6347ff84ed9a2e975906542b4d13451f5a96624b14066a909fd55837a87e51a26057b4f2a5f6a61ae51ab951d765a0e690e117fc4e118;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcb53d1b63c37bc2c6cc7f338876e8df7b1719870ac1e10c649b253ec819da19f8efecda9d45042b74dd4f85b88f7ffab2b604409e24e2546294f462eec7adc6f84ecce12ac90ee518aba5d3f4e1deb0113ac5a64a5d2000308b90160e53465765f1f2cac9bd266d32dfef1d4168d13d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83aa86837739f06d1e5fbb68417c1452dea08b579c8fb4dcf44b8ad16e53f91c73601c87450a3a6f0c15440e4429895c2b7cda1387ceffcc14e6228d28628be158a58513b587e5b62e30bb23783ec8571cc0a3861153a3d1f799bdabe0e00b11bc951ef62351dc03078d48e2f0fa28486;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a368f2a75caabaa8f89f4a057340baee6f020386b4ccb67b3f858fe69a7003ecc3a6776ef7d2ea3fb9ecee684d6dae48d9da898d8fa726fe581b5986a7fa3c264f3b620c726e65cc68936fe6ce24990f4e47868d5a073255e106a8f25801e478478a40fb8598d48f947070598a5bd78a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24516e52e2f4a9aca116b410042fd6f6d7c473ff7b0dcee645bae8f3a27d0f1d2cc29ef8c5039fcde69120f8177407ad488dbabd5b0d8df5ef61cf6c2b718032314b7fce1740a154d994e508136c86b8d1ab215b5b99a2d22eb207aad2a66d0a29e048a15cc7d2400e12eedf05a7e5564;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbeca2736ef5332ba7918af4e2fa909fe16189ca03b86c6ac3415226cdab88a8ff3f3ce8b8ddcf2a18405c5c2cf0648cae0ca641b3590f7ecc5212bc3ada8dfe730baf44554d92db48605a462ac217d6f43b0e7d90d26bb706fc90557012fd207382faa2decdb9d39f3ae292298da2b93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7440cde7263307533f642d1ad9cffc6adb04323c5b8e16d27acf67fc7a89d96439d3339c6427e9fd0e42c47fc2423fe978af2819bd0c02123b46c4f5a30aec8a3bb3c6339080920678060071047aa32e7d392d20d1b70c5c915c4c1ff8f95f093d1d8c7bccb0f2744e73246f1eab1182a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43ed4bc4694b8c844cf601f1368930d5e5cd33da942eff72b7158bb66500dc87f5a7f63d8db468ccc0e92ddb6f5e64dd0c516c27431f9dcd1f0dd5f8eb9ca8f0e431b832249798731c7e3cc13b2102f260581da4a07c8b842be7e3716d863e7e9c334068f09d6db28f785f0b1ffa6f91e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6db9769240aa6c5db1c545b9094b0d0f37bcc4942f4b4f19127498e9ba40ce5df93d62f8627ed57f8cd50f9ea194023ae912cb40aaca5d594fabb355b274a6a76b4d7bc4483ce265b6d6289226a3adec4f508350dd0ba48a71b1c453ef24fb1d58d49a0d8572687d3477b2a4413099bc7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf457ebc75072cb20c5a35153bdd303dcb6908268472f964246fefe949f527e0bd8e8be032bb7d63c40c6e1a7602d1a1a4921322b7fc568c0d56805e707fad830d3f6b37f049e7f81c8cdff48d2dea0c178b24d4cfb9138533a1d4ed19cd63435d83f2f25f8e51bd060faf9d0a09043f41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22e8564f7fda6326e21509e528028b7d4ce2458688aae461b3a3fc8adc9c80a73bd67fe45185f55dfd430b6d9afb7a4b47f7af247cb238e0f38fed0a781ec1f477510facfd2bf64a48c8b89a167b7e5985859b43c08c2524c61c7b4f34283bd14b0f67feabb56264bacdf0c2e6432eca0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b7bee3f4a4723a630ba87f8b2f4cbb7d6410f68bf0dabe34789c229b81fdc0c87fa53a11de1062e8bce106f1e869b4802921b3012a53635376dfdc21e3baa18775b6a6f9cfe1958adf59240392e153ed2de91fa760eb65016109a3269661d60160a6bdd1c3a260b1c657be84db32529f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0713afbc5a6aad6926d79991f6ded9a6ce3878595aefafe2897229c6f3b7ac1ee20571a018cb5f269fc831d8c79743fe950b763ab303f16314c331bf030dbf1360877c8367b932c53befc0a24408406bbc3517e3ac08ca7ea7ffb6220140c677d0032be11a0d5c997c3332c5904c0a06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49360aca1e521992fb4cb40036b5da8aff0e18b2c256b6f11d590a7ad65a9958cd35163a415730e26b26010e33fb624b204bfc7a3f9df605537546ab60995f71c9703dac74d14e30aade22e509fff2a5ae057d320cbff0be2594f998a54cdb9b35641aa0ca3e2b44a72f10328dca461d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ae9e09087cd4e2ae0ead9845cfa88f89097b2ba3baac5f226bf4af7f571cd36351264fac2266f7ec3fb358962a5c22fad983287c503b6d66e67ccdbd733c1a2dfa3887965ced4833d179034f7e2309fae6a01b309534f64c551cdebd88a1eaa81919145f45cbf7912a9d35db2deca4c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h918843c52ed3f9889e2c4955f1638600b743ea622477d028f0a5f96824baa1aea86072f5ec43b73305f5ec5e7a77c8328c3f4a4f388020d5e170c19d8c36316bb142c76d289e593fedcd4a89e5fa984beeedbb489aaa20b1f248867d8a02929a7cd4e649c7f1cab74c145e6d7095c0639;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31a7bbfcdacff7167a7162e669a9d492b662dd55d4770987dc118e0aa82852d9c9b83105c7c3608a4612441d8d508fb39408aaa31966b4ff05030562528e0edaa7a6ad39d8de823e0379c6ef36d9383614d2999f8003081114e05c89f03a03abcca694685c19b1312e49c42dbf6eb5a32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbb17b3e611b99486324715fe152b894216c5ff3f853b41905acda67290d9a5656b085a378b3049f3bffe47c03d39743066f55bcabcc153c65f5f73122a482d1110ce911a8da66bf24e6cd9f0c0da85fff6a00c9edb94df1fa1e6ca4db189868f3ba4e0622ca117ef30338b1ea6c79e3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32ababd70f791add1369ef37a7b74bb5d3c38657d40734016c80bfa7ed0dd44946c12dadb4abfac719b50f618448be92de0c8d292b991db433db94c753902894a6ee5c8a8ba51362d0fbeadbac6b25580afcfbad9822f534293435dafdd8fcb1130a0b75dca80aef8c9e0042472a417c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf83e765be7ac7a0906923efa3099f78a68d83ca8b11fefe232142c5e9a6889421ad187c70e1d5613e8c607487df9f112e14f37178b9c9f924a45f8080bc4e962a0b990bd36310ef20c4097938aa589b19c31bf011fa29508c30ae20f3b724032e2480079f35f5243b1b8e9cb845de80f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7caca423c11584a0fe7eb8ded25c7e377ebe9f8fb6e0366068871257f3063a8802088006b6b1482bfaed18921d0f8107f63b17bce8d7a4217314925f54a90e7ebd0c3199514c514d90a7018f898ca98cf2aaf2a2e8a5110e93daf77f9e81b433da3cdc3e4bbe825ce1a805b98ad0bdd0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h164e9231c97a688ea66000e3b12be0b93a7ef9714448ba54b7114298bc22139c3f349c1265a5559fe53a06468da57e85c36a75e90b3e26b4a2c01a0cc88f0a0387d8a9dd96fbdb06eeb51236167ec4b67b39f1fbe376d74d33e139500d0dc3fdaf34fe652703b345b655fa1c485a378e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9d57517084cfe44f748c971e5fd323b9d24c0734b8bca00a50feaa97b3d3e1e2d558b9fc5727e9013a21d4e06508eb255e938e5a1b7b0149bed02f673298056de7ce93c59a2229a7d0c0253d242fb14c15832a7bba8a93e49b64ebaa1c744091a91d59daba74bdb3e0b52fc0ddb23b09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7ec3ee4e06dc19c59706f0af9dc589324afb8c69cb537c3609ef31ef6cab7cd5916ce8780c5a3f0bc44cfff662f92098a2d66dc1a290869367e80864756f61697d68d8954f52049c25db3f1c241e4f8ea1e51adbb9e57cde0b5c46091d541e20e8eb5f00f2140c8392307cae30dac345;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce09ef0312b1f5c92bd5b0db6713311ae642df61eaa8e190abf281fda6259e17fbf6806cadc62574ae7f1e8329d3195ac10e7f1463f7766283d5570741664422f6f5b0db0bac1c7244638513460f2ca9cb51b2c9c79c379c7dfc00bc6f2b2869153b620d11e29f157024aceaa8e6c7d00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33cec14b08740397af0d5377ac3184e0fa98dcb588a44d272275c97af6bfb6489b858051c2f4a73edc470f6d1d452142dabac9912f60fb38dfe1e0720f04ac0be9e4dd14b6b5240517817b237b4a39e41bd8c57fa64f79052480012e3daac05a9a7e46ce61853becbccfdf109275326c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc621ee984de242b44eb4f545a79137c0e2d3d714cafef346f27306dfe41ba58237a591d83fdf83b1f779580d5f5d122cbdf7db384af8de0affc6c3fe44b2a400aba7f587bfad524126b27afc6dbee1efe66f56946e10e750d9b4a4fe7e7b03bcb038945b6ebc56893ad131822b849382b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h231f91461944de6fcba7acd00b99b82fd625d7d22a17d6225061a647770bee41005580f161e07fe3bebcfdeffed0793decdf5f61462c2659dad1cd008f5927ca0f5b964bddccdff3529bc6a75118a1b14349ff79f434210ee203644078aa0447e0538086807517e142ee699c8ac872db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43a78acc1964bf980aefc779cb5044905e3c3a168e77af71827b8534bd0e87e0323b1a9934127c183309ff6c4a7e14523122af03d523dbdcfada806f4810cad8f42d5e81ba9695ff6a757178a79698951274e4efb5f0fe389105a32bc3a98fc86365716b4862c7e873c99bd5613010ad2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h580e34fea0b5fad7abdc325bb57f908082e5828549b9a419b97315c042e90584ea8ab83b1b0c7176e319d021e004fb618859b8519ecaf1c314875adbc355b7806470f5c51e79d02ffe5c3232543c2ecf4f0bc063ee7231ad6efd1e0c5d76a1860d37a035c3998bc9f07e63f62a697887c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94c3ddaef25b04654712159d204d1647204fa2cd49b6f7fc044697e2757417ce2472cbeedba12d90e34a7cc43cfa1e2fba16557e00337558689d982c140e1e43642c759ffdd71b74f2a3406b6329df169f62af961f1ed09ceb7d02f6313e396fb57385d47334a8cc4fb5044eae2860073;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h519d95c2a0be82719763dd4b935f82f396167e950d1dbf53d9291f9df660ccbdca40b6e7365dd2d85ebf39edd46a6f10cff0b55fc71d1a6a70ca99f2bf93faa5653bc83f0e79a9d6ee7b591be7678ff1799b4a55ef4e87a537ffd5e158d3e5c03e8251af17d0692a4f792b55d8f856951;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15a3d50c66c3d9f473ec0e9bda1462ccda9a35e593b06d823392c3f1c19eb32678f645f2c23d5c86c16cd8c3a6f5688dfcf74403671199bb8bca6acbbaeb0658d577c3227883f7fc855564264a79196b0aeebf7e29345c0776a57cb8d01ed6eac2b136c2f6ff7c5b2bf10efb7facc8f66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fc84813b889633849a63571f060d1b8ca1ced67def8a260aea46f25cab5eb24aa53a2cd285b92dbb2f2f55d3751f444758da913a7e6402d0be976a6b4174971b9975726d4f8a940597ad06b5ea0f88a14bbfbc259e2e7ba21bd571bb3cfc4b47f0d7ae0dbcbebf1fa07ec11a255da376;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89823a92d1ebe858382793bb6c23d6d7ecfdae8147328e15633a1d7911712b3401eed26275fa37aa7fd433f5ef1731e6e60dd9e467970cac7603e62f072f0b7b877cf5205679b5bdac8b05facb5386639a10247f92ce9b8d0a09a8dd8672f34193a11748c0440fae4b5edb5e07f24bc72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7c0be6e59d8adfd1b086372fe7023530b146ef738150f3e1ac78d8221c91de38657adeb3726a74f293efc09af436603890e888c219ff6cf65c126099165699ec1aec4a123e0de71b090b7be598c118cc39a6ed26ce4ee2b30fb48385a23797ffde6e8d0792643955ecb6610a82c3b9ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h790f20e8ac1ce6ee7fa67080db040cd916866493191972a4ba1cc4cb173e4452c1121a94746744f818a244d2f56a8d925afd81dd7f378daa40cfc5bcbd844a761a80b60d607ed7345c79371cf9b6054713a5f30d1d608dcf1ef8e9b8704bc3795cbe321879652239c4f8b03c2c6556e94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea5484962a9cf1b9dcd3d23f1adc8a7a598905528f1cf6ed1942a63644bf1e357a4df16127232aebe507ef733e4e271cb02f91c9ad523a46578a0acb5fea44929543950879658ea7e3f47e63a0ce519876238a83ab4d8d768e8c7f5386640893f58ed0ae7c437e1f8910e6960b3cb2843;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13dcd53a999db1f1443601cc05adfe0ab01fb35018311ddec8c3713b694955854931382827db18b3d486b8ef46e0c9ce38918c22aa16f61d2a4ae9287c26d3bd2de7b11980073e5a5fcebfa62e7141cb44ead0171467baa1193008a6b0da13b75efa4046c5a5d1829938e6f3dae4efc6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8894530e58f3e93a748a3f6d87bca35c2466e73800f8dd2fcce1518ab29d29c7ae9945bb24bbdc86fb2deae452e222e1754bc5946b6836f0e7007bb7917492bbac56c023a756932b0887eb7cc6046e58a6bdcf1f0b519a10ad79d29d417675d1a3aa880d4f0e840a0b961f4bf637a7474;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h796a677a35b5b0a76a503b53cc0140d90eee631654059a95608453eb5faa2e1f7256e0215f075aa9ff79c59d3f8eb84613d55bf46a2a921dd26e810b1913977944542591aa95b8bd9689b64848373e3bc6062c72ec84aa79321de48a48a4c418c21512b21f6b7f7730067e2bdcdce4164;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf415dce4f6fa05e97496ada5957316899d969a4a6ee4ab459abbf5a8841ee188164df6e3860f4f61b37464b1e6b707db51dc7baed91b9ac0dbb9022f6e01e4c6c087009961fb053b659b75b455b818003e1948c9e47e5d1ccbae5a245fd5bedb196d9280a3af3c2866ffc5082aad4c19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e94a37f9fb292ecd95d223d4f3737eab01c46b472038858e2e2bc942f37b1778ef9d5ce8975d07eaf939900cdcf6f983368ecafc2c916e2a4f7587d6e70b42fee4887bd7c65c4b837c49eccd3fc844e0b23f684c880a6e38404e8d27234b0f7e6b89beb53d142eaea7a1d3f19f422f71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8cc2c3a67b8aef628ff436115b34e47553207085baa1e047f885748a5f226c56a12f99df7d0aa23f8888dcd31cb3a975729b133c2f1549c5b971a39b5c3edde93315fe88ce63461f11162ac3c050e92746aa59bea6bcf01946dc1f330fd088989861221fb195a79dd6a0e8f98a8c9d08;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6228fb7ae6f3bf5bc324b8de2bc61ddc82be8469df98841d17171d6debc261d38d8e6dd203fca4c1046c95a9f3aaf5603cfe9a2b696f3c5c53816da60143c3a7ee97698a92946613b78ecb8c8dc057a9bd28df71b1a4b1fa485a117174208157693278c3788c255b345926475a755635b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e74a29c5b67bab7e071abc225d79430e119a5077b8adbf0ee528ea2e2be868e58ba73e4a74b0f175ec87c6924b2063ceab9c66206bb73e9781899004f781499afb6a1cdd557870596dae950fe65eee914bc2acd6ad520938ef2272b29a68a6cbb18fa627bdd046cbd868d9308f277386;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9db28a8ef6a3fee7f0679b1cf9750d13e796dc839793da222e929091a3cdef911211c8eba7a91b4d3e897375b5272515a115c18d503fd40aba126215d27d0966b88ed9efe8c61c4339481d67c4137931d786f9b147c7926d5ba4a2fdb14ea794fe039315e9156a2907519dd0c69688771;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5e6fb742bd8659ba694eaf94e84e0b275d6014780494830287e446ca699e1774e2cd232daa003b06f569efcce69bfd5ee06d168da4a356a0ef3e8cc41516671a7d5cf9d352e9eb5edf1df6d42209290f69ee77d464f5d321ebb271a598e766eee4364c87c758bc37083d2ad8a814c162;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf5be41388c1208b1a84c943aee0d2fc4fee794f90cf873d509bc6db5ac1e9cb0bb00d46f7803975f49ebf5a0b39666064f09aa46268b160b8f7d8e8d9ff9c9e0b080ab15d74896e18561352c065b61714f081a16de3c76a0fe1e678580dfed1ac2169bb14e3b0c3575ee32ddf14a1717;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd84b8880d9637f4a5703bd20481d299d2df0ffe254fbfb62552770ba0679783469f4d81bc41aa8f43696a56b1f75a8f5175b6d3f20efcc2e93af674a5af41dedb43f186f1b06ee7ec3e0ef851cb00ebdfd0b6f1032524e27b1a607865c4822a2ff7ea05f28465207fa5836a1fb353580;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd889f3e0c398def9b62d237a89bf343de24ce72c7df6d33866d37de22f5300c7ea7ca6022f02835067dcc4065c41821a6f0a13c3f1d42899c4b5816e7affcb99d627c63b74a37db1d486562f738e771db45b0c7b9872f055ecd246fdba0aa6fcc4bfae7cddc7d671d68081522321722;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d9c2c9dabdb4d9e60c5d4ad5dbe5f7353bf5d9b467280d9174edeee53f8ead738be326fc2de4400c4158a7df6516b0b45f7e02628db9ff03f3e276b3b11408be06fa376137e5170ce54ff7c4a77dc5ec72de0f883e63d14689d7df31f9fd9904fa5d5606d8b48c386c651e76b994d3e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93e33b5854b1704ea67fb463d3a8c12753132810967bd4c7318e25580482fc62d146bb78e8e2e8a262287a70b8f143b6d764770747e26fb1316f6982d5da4bea630c43a584350820097ffa6ad27c8dcbb78ffd6e1168a86bab991a44df6712ee657e0c9414e6908a6df1fe97e272392ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16e4e531f7f427a59c1a51e2bd8b5a47c582191705fde75c90a6a04274557dafad9d5b8a7166315e559d07e12ead140fd54181ccf7af85bac7d1052ab89e07662ebbca53799abf931ba22e8334fbdbead82d74a534295c2e3fc4e4af044b021801d4128d374a22a9898ac76381b26680;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e65ab669a99400268f54c067c9fed70b2aa45b290717884e08fda8d5d45b3932cf3f96f768203eb3de9b9b52882f825ea3d3704b2627a39619fbae35dcf1f897f76fda92f611c09944a2c6ac94ed186e1c8fec6690278b981fdfb1648c9b110363d80925edd99de85b98d165bbf2fe06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7cbaecd59fe60d97ed9512e141acbd578ba999d6b4059755a406c6ab9ac7bdeaab35906b8a7efccb69fb6d8eaa7b98657348b2f7bba3c391a5d221a25f0ba9a70b785569f9ed06936587414177645760e008c249fd299b8ca6838e385b3c83288385b0810d9b06d1a2ad524963102101d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75c69d8a99f1820bc7f4d129955972d59554f6973aedc50f27a2f574941e5f67d2a4db0e35a7fe0bcdb7504d9448fc3ae1cf9393350d767e1f0ffd9b4e041563ce89fbe6e9a378330cd39b0c79d2cfff03fc2be712cb1e2d875198a6e63ed26483bcf41d0981d7f5a7b9f100cfe648a03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe17de83fc1453072f8fcc97fbb07ad7842e78a2cfaad21698bf66e3623ada370085bda47548a493ded06dc093639f0fab01373abce580fd5e352f7e70eceb7ca6a3b76413b1301ce919d14ebca8abb220477589e743ccc645147dd2efb28a89928e1e1256ae489573dc744d7fc586555;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fd7e2ce4df3595dcc2c82c7c586e77b02f8bfcae433c102a5e1c2939331b061d4fb182f53c7304aa10e8b8909564a819f4a01352d618682f2e6ffc8b7feb9ec51b8a5dc793cd5bbe3c18ce78b92d5d01dd098c723fc2d80beea0d27a6b049e9d7893611dbe8da3b6cbe6e46b3ef55bc4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e6c440a7921f6798a9e5b4193bf9102960448a9736b640454e5a51e8dea6b9f27475496986cf35f688efe856b51faccfc7507aca08adaf5f34ac2d91226601c8cca5d293af1acbb88f2b1e1ae5163f48df3d1518737a6f9e93504a4506db42e20a19a1546a95ff11e79520ea52517908;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0e9f4e43ce986467b066ea3891bc073fdd457359e6e5baf1e0d3af383c998b78cb8118e2a1c2c1227762b547690876b480e87e9442f88b7be3e668ab0e9aedc4fd8ebf771f72fbef49098504bb05bf75cf1e28039d33036b8ac90e79f4f20230ebabed7fa87dc268d4cfb26aeee6a5b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd048603acbd98ed2000508902869bd7334e6af1859f807d927b49a501c80fc7998030814ed7573f2dcf66b2156edb7bffd1012ed67acc5025e5180b8c7048e609a42d68be5d2b46672c3b84cd7fb298528b34076577bca4c78e2e26b067af003efa5cdce8251b6b131afb06ca2defdf8e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe9af673ba0b67bb0b175a146a7f1bc6ddf631e60782ab8679f65960af18af91e553598086b8777675e86aefeb8e4338fb96b87af2a5bfdd87e50855bfed71ce0df1a42ffe3bfad7a431825e048a80b2199e1e383495292046305adc0a0e7c70ab85d504cb670d84c9f22464332a7d264;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65994ccf5b306a87838e45d08cb45838eecf50ed1058377e61bad21ab548c84e5d9a1871daac6174a97aed80bee3701b996c5509dc2b57a19fa417c9b110e83009096afd421aff58b274b31540277d553a3b56b97528a4f7a74466d775ae891ce83d1e3b4615c89afc40bc3a3bfadf073;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb660ff12a8b7722be689bc2d83b1a3fea72edd62745b4a1651bf47089a87e50c8f4eedd7a7ae6d979b03c794f3e06b6a6817a80ec72c4a1209effcbc2d2f0a250dcbbefb4c0d742a77147e671ccf874d67f463777bddb517c839cff45d9bb0f7816f6ddd304a4ed458e0b15532987f82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c8878e3afb181fcb7d11f9d5eb95033dd57154e2dc8d15a245ed06f7bef4b3b1ed1a2ce45dee191bd27950f6f7f12a6e86eda55ae805490eaf83da793502685e90ba42d25c22e8a78c3c61fe802a8eb17810f2cc8a07b71859397ed133ddcb9dcc0aa7bf5cfebfd4b9c42d3056e78a5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd04edc8180b55a73a1bc94c0636cecdc4150261fbb3e31baeae7c6f41cdfb0a28e5e0ca243cce5a72a43b52f411d07f6b73f742c7b76a5d89c6257bf59684be523a4b4b3a6fef1c340719b5a3e9f5953ef89e95701b9e7feea285f69ee508281dd6ceac90f3e6f22b8889ab294d38b7ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h324df769a05f1879dd58ae35633e615e63cde5c701d418af2b859cc6d859b20df8e77ca56d0a68286e6bff98fdcc9935537b8ee71b21a67fe69a5986f5abff816074e7114a16fc157b218ff579604ef2ce8a48b8554555e7c8f1749ff2aacbe9a33295ae2928d799a85c7347c11080401;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec2e846e949a4b2072ae0d8aef06fbd215445c1e03cf99176bec700ee7f4930cfdfd128fcbf985813d2270c7bc3faf32103b27eeefb344e9c6ad8f7a38cf6ab50819e024e9b52e526c378ecd68710f1102474956d6a65ce8c56ee28bb4556af4b6ca5e2ef6f6a5f510e8d0a7d1585c880;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57432eefd66cd0f4e3da42b05277109a02528f6ec4337779363498d1d51d618001e1d0701debe509f37e140e0a2bea226c035b95c9c28d743e6d8c9d1a6035e01f98f69e35995774ff6f49ff300827ac8d31d5dacfccb34367c5952e1d189abb8ee7aa6014eefd88e306bb2f8cf59b222;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had0dac7d43be66d7476c7d0681b42b9db5e3ac3abf6020776440498909d4646b53ede40e530e18b6e3408c8dca4e1741b3191d2181454aedcfad132bcf62bd1198decbe75dab889b3161c85a3512688685f8e4e61d9ae1eaa8500b95f929067c0f68e236b59c1c43956c1c8119d387ed8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf19183acfeadd86abaa57eae6fc89c21f8366dd0d7d3f9d143d8bb4368d6b3785c369cb85e8efcd3faba3d7b2894af1db85e1e9f1b7ec00fa0024a1300e9d051fc400f905c816bfdeea206b9e0326843d442d045a62d6e76b527a072965f012b9227e3fe78ce3be008f3545d4f2094ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43c13ce2e84b92f427cc14f8cb34d65b4ff08dade671205913a336e32192da6b5a75a49a805f49020c612ca634e34f88bafb130a170d8030832f7f036895b3d8497bdfa28682bb2c5dbc838223980fb2b2f7aa18a3e19208ef6460332e40daa1a651bf3c25dd2f75723b6487f639fa143;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52c48b5f399d2f55fe4323c19b1e6a68ee495b831830b868d2ddc38b490f1b56c12532cd27f04716229d2358f7e831e0005713f5fc0e878ca80f8d4e74947cc16c0b587320c367309095ea880ba0612cbb73c48280fcb9c88a6c913f4d62fbb9b9be65e47c2d5a121ae8dfaced5127cca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bf9eae2178e1333f5df28779164a129db95367bc80a928cde7f0809c53cff1427825a56156c7e6f4387425bc9fdee31b78b15a2a2be8280fe5cb50328e4027d16c668c15ddda889d3ce14cc2a8aaa622d3e216f50ee4f1b1ad4d330a92e0db14fb2bcc217137d2fcaa752774fc52fa1a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc22c58ebe768cc8a1e39b83e8f29b2beb86bea599f702c2905f9253b4ce5137dd7a0ef3eb19ef9655b274c0c2d141efd50e6133418887e915771ac9908f26aabfc4a5dd1c839911b051baf5c137791f4c7cc65621f80059ea307a3ebdf935d09f97909c72487a28f08a0c34daf21e159;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc686c19f8ca2a6289eba693c2e37146ee59bf478148805c9fb29191e15628164f5f9e7a4bf600aca19ec74e4c756cffec91a27b9ce5dc9c32ccb33f7046fc42dd681908fb1e5e5720014a01913252d4f3821414f82727d45806f1f19b3bc30208c7b0064258f13f954476522162830b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h997ae63203c4906315b2feee6d500420121886a128589d28c6451147869b7d6ac9467f0c9da1dd74963abe115ba52115435f94c8abc373a7e039c43af34d9cef7c6e396bdde5f5659a05594f4724fd4a6be7875175590e51c8c8099517944db7876353ba7a2b116d4050abc652bd0cf57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d2c18480b082fab309a1055d13ca31db938b1119d0b9adc8bd5461110f25a0e2e741ecfd47e5e9cd97505bc7ffbede9b0ad92d4fbf5318fdf6d67ebb74dbee1eae1a2956fdd412d7ba6073c8673a52c6d6b18ce3195a228dc1db4fae864d28887b4e65fef2303c03a9d3e89317f4aeb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc73734dbcd47a478c9e90d27324412ef8d149bfb34a2dc1791b435a2e18e8f6e2fe3f6581a9e61f5d5fc9d9e3db1e9f5fc97d4a72feb348429a7935daf8a57b54a031953d1b7854bce8ddcd1dd12a97a346b93abae22a047305a35b1f9276e349b9fdac5e12a0881db0163e7950e009b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h745cf9af52df7ff03d0754ad5a0b8c2140bbeb8fd75dc1c24ff48cab3003f1a9b065d4d95de3ca8694a7eaeae97ed57253cbe1529a22b90de345b2fe3b828ffcce7afcb0adc050d780b27a0baaedbb9d21fb8e51099df231b3fa1b8f9dfd1676a36cb461a443e234677dee9d802d4d618;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5f57b7fbeeed2203729fae87ecb3c44155f0491eeaa7acc7c78ff8a29e50b86fecc04d1c92c2911cf67d0210dce9c98a0b1020685c0a8493027cc116915de910f93376f8012411eeb52bc8631ae0aa95e301a55b37520f7d61a75cbdf8d2dd5ff44ee1d381c9487f1062c3b5d8285b4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99c10acc176c6be53364ca91c77da58e1f4a509fed6cab79473d4c4f615686e45f45e564a3b24a700067c5a50473f5d4fea155c991b0dc3b6938ae1a4f906c6cfe18fa26cb104df19f1f3c303c4b7e47e9827c533287078d8e75511e953e4db31aecda0e477a685465c35f46d70e0813e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52efe88ed6ba08345a9a4537c461d16e04322723a05bba2f507138a748ad484c5503daa38d81e7ca813c4c07f720c3371eb173a55464bd5ec92efe6b2cf5793c20b43c64e70470418dd8d890d3a70444a164652f81a0b53602982554631e962755b378c67384b0c4b5c6561c8c00b337c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5afc51753ee3edbb1eb1157a305e65ac690a61290478e6d7d3c06de78f482c4ab6caf845f9211ae211ad8d4621e48dab607dc31ac2ef0c42346e9b40c7dca4ad94f460245ec0949929f55df8b684aca3c7f5a6dadaf85dc045b3cac4b6b1809a25a736777537f335380fbddded756e4b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he30f748272faf921519a3a3a66cf9a1209be77cbb9200feba4b55c5d606703c0cc58d388c63b1d8d749ac171631b545730d2665c4e0b7705f603dafd45b2611cc21ff4d46481ba50ecedccea97901fbda7d57791940e803736ef85a372e8e39023a7c6c50b193e67f164490c2e0c539d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1b3cf60250e12ddbc16eaf721f56e87aae3376dcb50ca063a90a61b86bac979a3c5525a18888594f1b5ece4f81487df66f6e34cbc274894c10a923a2da28812fd4e9799aaccdc464714f8895328226a1cd66a0c973bb38ae0078024417f506fd3053cad573f7a1d0f2cb347c13ff94ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51ced6c925f028c4def50d69ccb18ed813d2e6c0198f9ebaa8c1c22acd51fbce9881d73ba84d38a7a3675d2f52a7e583ea0222e29147a6b6b78ab6e40b4fa60dfc2514a97dd157b38cb1990e80e2664946bb72ce416806e6c0ce8b2c389e938b6aa76c7a96b3c1352c73fb71b0d5ed6ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h774771588725ace27daf618c9d6262d7504922b8824d43bb5ee7178d0413ae501ce15dbb36a347678d082381a7a36314df5e49a6a0c5f5a3bb1a0a042489355fda32c268940764aba749bbd62dbcfe3a219f986979163026b231bbf84af62d00928490d6ec83e4f2e628467deb8f9ed4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56704a9966056cbe7f6556664e412af17478444f5a0dad61954320367cb988ad5946bfd5974f45876c27cb391d80afe2c21104675450db1e8b05e1f02b0633435c380e813199f70f0373ce81f49d60043ef5d2f618d3cb6960212be243c9f26e1a294e64578484e552af5bd952ea688c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11a898fab1df410398ff1229d09820bb48e2e3c6eb5b3362c4a9edd9c187c122808cf6dfc2e912ecd8fdb561345e9f5a0ed6e663ceb04beb6eaa61d6b22fb9f21f2bce7af094fbcc727ca4ab1c05de1f8c74c0a909d2425c772e2f196832f6477e5f3ba868d7159b7e68f38f8fae074c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32cb90b69415ce450196d7e0beb61694c4f1cecb0cbef8aa33f71700a6d28e6da7efa19e708751db5486fa104c6087349b19df4d24a430b0935af6107d87ec06f8cb4447b0e60c5a72878428074403ffeced8cde1b7590f33c58c8635ebf135af0b052622d1307dae484fd3f867939588;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a78c4260ae7ec72e0cdd2c2c08ef6fd3febb74a5212b5234d003d889319c4b27c332632c4efdc721cf5590aa8d5bda1d4db7d73976a203732c80b949f923f41e6ec5e65ebd5250d87798a52782d6495ba1ab966f0c52fb2c9ab6749a89bfb7f948389b3ffebcd47555ae0e191ce72197;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf04dae491296eb6721e2b01ae36bdf8ce563724d71c4845f226e2fa126bc92ddc76d1752a8eda24274496b23edef8eaa7e32c82790f9fbecdbc6ae8e2221d72d815c3309d9e237be1f9a595b85eaa1fcef6414c87be88dd934e7245edd75250af6c7c97a0d5ad51932f472824b4d4f42f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbef3d75075a11e7eb819702aaa87780650310bb9b2ff5bbf4f565153f93ea5bcca812b9e6d0cfffc5a0a96bbf6590c916934677364ee23adaae7fc4ae9b6533cf414109cd554540c0e84cd5027161c40da36a4f01ce1cd50a5d85c0d085d682c5cc74c10e8ad874f8a4c74bacebebb15;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h101cbafce69a9e322546f55709479549276baf7af3e9b6846f7de3c8f08ee19cb7228842e95582831a14c6b202f08b75d5841b0e0717d27d12e8d2900b27af083da69ee40ebf449b6a28899c4c0197126be57d85b47f2e62e64f403700b435a93818f058c7b20599e7ebaa6dc75de73b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bf781681ea76f255b448807ea884cf79c3dca2ef3faac6659ed47c1cc00cd6b8f1d426914d68720cbeeea4cd05141efb3d8ff7054b6b9faf77148fefb326043330e394bf2299573e46f5960d869ce137fafadee89c466c62d64f036c3ddcb9a1df7ffa219ad4083c0462dda150cd49ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60f8db822e348e72e163e8a46cbd14579f41cec1dbdea15fe5452e990e5fb3f37279768a7f1408924ecf7ae726cb0403f5e0afcedf32abf48dbe140682737c0bd9bb14600542b03d380bc7445534334a341828b61740e68e38c3463199d2f999423c885d94b82fa11043b782359cd3dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38e60387c01a06050bba091c59ae02ce5d3d5df66e527da1fce1b639d36bf8160b0035c50bd67ba399b8ccdd91a0690b0e063d1f3a95eb09f4ad4ba79b8520714029e7b713f6ef78c6e238a16d3044521a1b7351dc6994933df60e114d1b4c70ed8fca9555debdd80855299ab83dfa65a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h486698b0488104c48fb6cba1178a5c2a24607d7fb7f70b83735d68d98256b5c5d9388b3f3fcb93cc3d835764050ed06215cc04fd4597438f77c15c9933168b012ea4d3c9366541abab1d78cf6d26373b74278127cdd69c502d034aa3853c5b1c11446d090eb53404c6fc764a7acd71236;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94ee3310a865a28df27a9a7f6e03b1b59af6e76835e5a5b0daed55c1ab3923021b09886a45fcc84957327356a9050411c66ddbd8373a98dba7bf64eed0c35381e405e3e07054509638715d5a886903a80cbd4dc53a5a3bb62c79079b97afaee030af0fd864e71f4113d3033f1fbf67752;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a8c497ab9bbeacfdfee90080cf71f19db139397c44da9908730d380ba1210580db1d7fc26ebebe2aafa8acdb4da7565a0d79b06e42f0127529ec2a273701e477329532f48be6f4e790240680412d60806399cf34defe44855853f2882b917480b0e459d5bd7c50347bdd7f210c42e10c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha874bd366d069d0607059a4e4661c8fd12fd7ca0d1406fa1e4d8909e22256b28b85e12287af887415503888450da13cc6bb60ad32d87327df3c88a2544394f33d7432a9e17a9306c52a06725ca7e8f54062f72e3aa5fb37e2f6bdd5643438c83169822362188bbcdd5ec445528d730d25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c26cdcb482ae69a6611307919e492aa21e55b7da355ae7bfdd91a5b4aa8e0f0c13fbe06f75ef0d554b2df0338cf057e67caafc2a96b1ec1b100fc8484be5d49367599714c96ac36f02329c7028e7ba6dd79d61c30c22d27f127d26a38bc72dde11e6a69107a13cb015207598e913e5f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbd1be5166f033c06e484076d88cc29e7bc324c3b295675e299e813222ca64ece9388ae3cdf395e1b858f948996c15348f1534aceb9a41e4efe728fcdae05ff751f49eb237d44be7e787244a23df51a94a02758bfa76872a0d143be255daf58b0da2af0b54908bf142b122b91af9f6f4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ba4467f8d84b6c2d99f38585d785a6f00dac0a8ab9cf836e06f9b680b66613fd796f25e0a0904670303dcfa2aaa9a80bca03e889d6e69fbbe312869877518fa57b98e41841b54640aa5bc4d7ca405b0373795c8e31580e12f61841825381638f20ba44c0ca6e957631bc567d2ce1b3c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc4477c6b059992408a9072e5c9a38f988204a2f7e436db8634b11c04796e569f1274afe6770c5a8ad1d3e2f29ed3f9a66bb08ee26bf3a4f5609d60866b1f7281a47249ba5fdbfb5ca3f7705d62d89be841584e75bb404deb98ac4980eca47811e71a23a1177d2baf88cb1177ff60f480;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1e79a664ac15a87fdb83435bd17be1ffc68399d4ba75dc1af93194cc50c1c2669034ee624d0131cdf36a7f0821b5fb021d12b7dcb557cfe8a715e1055f6a9591423cf0959053ece1ae7340438aaa379c28562b1981142121f13d5f828e305703e33ff8cf2ac1e9d8280f8ed8880db9c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c1ff1735d213f369528503f18cf28d1970b1d97ae82272dcb996457b566021e104752057b8f87ec3a619f7725d31a3e8529a4e0a65a13d75f0ae776bee9444c59d85e9d8f4db7bec19831e2ba633edb436df9e5041ee3ae915a30b568c2378c18fe36b6c262ac0518817b0ebbe0da7a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3e1d23fcfe4258d088bc12927d263fe57c65b272cc9c155f2bea7a06b6040a31b46c4271f004c79fb27e39bf0e01dd55bdb2e0e805d5ccece700bfe0afd1b0ac2f77282211376934eb1798bffc34c69281685b7e725ae2a1a94503051037db6e41fe25d9611286aa37fb69828fcaca6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d6094c575169b36c9c864166e2066aa1ee4e6a81cb7a36e0cd02043a068788f9fb8166ac40b2f02ee256977add4d64612ec04505b7b1ef75ea189203ea0a32b151e9c32f903755d057f314f90253ca6915d6f30c0acdc91c81b94b2a3f6c20a493e5f46a59c96f9cfcc7c386c397b0c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6786d9dcdaa0980615e9236e2397ca088a929029cf01d9e7be728f948c26aed58c42cbb28acdeceec14958818d6d71aa692c9591dd41a57f919e0034896701c1e2975408f2c824c33c0635f71984d98ab5f95363c75530adfbb792490fc7aa27c2a069a5dce2f973956c06d9b5cab3850;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5273549e1de8b3a58dcf2dc5d002f11970e9deeddf3eb9a8e37f1959ea61461179d26b6ec93979de2c4e383e2331cc22f4b421d479f032ca6347589343774c226a5aa59e25f8fe94cc585586c8588e95d34fd4bc0dd890c2a60b85e9475e2cfc7a7b162c20a11c8caf2543b37875cf38b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24e118e8341507637a18c038f248fc6229ae930b1071151f3d26900c1be0ab522cbaaf7cb35c291ecdb37d9a3fb3c0ec2ea61db8706fcd6fec2985c5f1d78bd5bc945258a32dafae33c800a88b1f6f0059643fbc9e894742497067e5b01fe844fa766a29dca4486679c67340aae219cef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40c58556ee80273869f4661ca2cd1026fae56aafe6668f6fcb0b6b3bcf69aa63cc64abbf3f23dcb6f32370cfeb150dd5551799c9265d96949d944e89bd4b7b63ff412e85bfb01f11d9775932f85fa534bad699a3ef63b4e75955de37ae6c30ca32b294b2c8fffd874e23b6699fde062de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b513a71c8c900099f30aaaa45526a775f07f031e5dc21883a04a606c02af55b8226519b7a22539ce040d2598477590df04e650b6f4b061dcd7c39b03cd2bc21be9f0c0cc6ff526b040ae6ee981a55e6048df26f92b8cf95b93645cd1c00bf5aeae75845c94f74eb03f71748d87d111a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cc3c14492889c25faaeec721438ffbe82c3be817faa1f82a3b2210e8ad6881f9be36635d6c9b048373cac5947c9088f723dde7d38fe40860422847f5b77e30332a71af5d06b07e7979d958b06cd87fb6e0f225a36396f04fe587aa633d9a659ff07ebeaf6b39c7ed47e1327ed8ea1ba0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a723632f6f8457632bc0ccd77f32a4a84652c110bd631f7d95bc49f4a4c0073a5cafecfc2c83f1646f55a256c8d875ab1603b1d28d18725e58ced588bd4fb9e8caf3cb7ec49ce5dfc9cd9cb6e83637369d209aa8e4c5d25ce62dbc17d4162ce735bcf1b3fa7d0f5cc1c58c4541fdc908;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5580d0181083d8666c05c254b2508a34944991aa4d0f6a6f46c51ae462b0fbadf2d0a73a3215a31118de7923a0fab3d5b74b1fc1a02f86077ad6718d5a89b3635a7e1ab502b19cda744776638890f39d166d7aced5287668a388e8e4a19cf6a2bd71cc7f53ae064de435fff4c2cf7110a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce3e585d80da8462fed163cac0d1289a8a9bfaf04b88f72425c21a3f3156873eb7b347b90dca74cbefb4f5a17cfd98c958af650ff5a24e204d13c8efe9180a3094eaf31d40648c1494ceff34595cdb88d34b0b186140312f31d8fbdac2007825c7edc81e905982d6191633f23ebe8308a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b0a1b9aebfb2a5825b593c4cec569f89789e42c67846ce755fe4c26434a4c7e575dc13b2c12fab3809daeca3bf652209c2debe5410717e36c8bc2e824f26e602c1f43398eb420187f621b10fa035515a91d624e6fd80230e4f4e2c2d17eb62fc493da617981f50261204d7c8952ea7e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9fddc3263f31fded72b07e8bbac4d41abaf3d9b5d2e633b83f72d8ce2cd4653a0ca580c25c6725684c22fbeefa8c41a57e0e84809125074ef44afc9096def8d37cf97aef720fc7c8347faefd0264fa866e3517db31fba9b5c5cfcbcb12de0ac1c2a14e997d741a3c43365bcce1c26f5d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4516f68b94cfb055251c3a2b728cee11d5bf1eb27e67fe84b8a313db06fdfe984ec80cc430048abb3a335aab974efdadb8ff26f46ac5c5b9cdca571221c5d897122533f7fd89d72b66a0daa6ce414ecca2961f4356da0e4a6b75cba0bbbca3f0514e0637e5cffb4285b0cca18283674c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e52c45dcc8ae2b318314021b295b3e8fc59ee680558aca1a64ce96329adb673b0edfd9573a4552be9c90d8661b3208d209dc5b4f5c14924642589a4acd64a800a97bb242110692424e20278137550815dd2b34b50a31e17c5ef401426332c89483aa68ec5eb0b485f840d3678a9dce19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5dce5d6365be2819b412cf1f26e393b5b3d1d1a66ec8426bfb03ee3abdceb9a2be041ecc8d26dd6cfca11d74a3b61d77b1c4ded3906391b28c531910ddf1b21c609614ea33166f3dad835b68b2aa565171a05005cbbe8c1052ee85a61481c38a549f689d8bc0912751a0cf55647ab698;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d2d6cf2b9f3e285497b780b4c127e347e7a19060de5c92213d00299960aca5f42f614c612deb1ae85c5a962234b7ea92078efc55118a64b7c3c49d68f9d46a8b18ea699261f552bac47382c0ede7b18152e64fa4cdc9a6ac83059cf16741d4ba886beee27ec8c82d4f34fa20e38f5b21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4f5e3c5e86cafe9ba647be784f3c036c9884474bd842ad24d04eb5fa0ec01a154ee50df2a860b9428f86d7a75e7588f608ddb51a8d385867bd2be23755421494531f0235c186a7758135490f1d5ed24983c7928da3b660b973deb8c2c353ddb27ffe367b11bc6211e7ce3f7ff1e48510;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb491a63c1979f8c517de347d164eebc986f6e7bd1f5bca4cac5afe657a746088abde640debccdc8be8f2e7a8a6e8e74172e6d562298219be0eff3e423e7537042a09083eed507c2c010149d15d0c30423c1274bb91a3020e810cb87f40dba47ee3240bad171cc5e8c84fad65387d8f51e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcd7ab191e6d8236a27f9d8a77bb2ff001f3544bef6693331f5be2a50275c2c49033e7d5b685a56a0fa92f57ec6b1d956653cb58b4729bc1015c2a1d107af91845837f291a12bffcaf928f96fa63b5b54caf4f345a772ff7ae2fd7c86b04721df52a7961d43f3e51d0086c5ce19856f1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf59fbb170721f3613cc895d7b3e7ec6f7c62637ff57fd5bd5c477e69a4fed5d807b04fc179503847f7a66e035c444e7b5fee3aaf452f5394830f5d1e838da832905563f3e50318a58b0861e4b9077b5dc72a3c95a5ef6b59f7b81184882618f09d243f06c915f134440ae42db4cb3177e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3281af889c0bc475dab5fa07dcece9b5358d9b18d8aed9ef81347b2d8d5e6333cfa82ab26c1c4cc6193eafc303259b15427627899a65f33af983955c8a4895d98090eefb82f449347d4e653ee6f6f95e0609c7560429ea3dc53713644a45f2293bd9340441eb645511342de8163a5f01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31f266660ee7a86049b2cc8ea81b0e2aeed5b6cabcd0ac268519d4403211638e80ef1932bfa07f9e44e1133f9c7fe0bdf3c27d991929d46b5230426edba2938b94f9fc9cfc1b2808c1b9958eb94f0d03487050e36c555f966881d9c5e0135c136b9d7add2299fd1abd53e65db2fe68fe3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ef5bac54aa2630a40e6648ec0d41ad583a6d719da1564b920309e27b07ea0586f5cd11d1498a8e1d4e1fe77a875170b9eccfea2b47fad95d9c442c10e196654195eb16501d01084abc1fc6f115c9f024a4543bbaba6abcefd903dac1cff8beb01417193c1f45eaac367d7eb39ad6193d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4230098182e380ada9108ddd0a1c77e9383f2fe53cd2fd50485919fbe11304c258b290d597cc7d9a652aff2cba364ac66bc2486d9856d45567faa6b6708a57e5552f53b3f60a0da72e58c86aa4402ac3a9ab6c5bc9e50dc5b8a7eec42b9bbf7302f18c0766aadbacdd0a4f700ca02395a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc584456bccc30eaa25fb33caa6c5cbea1e4cadc8e545cf1ee24d2653d131c02a7de21cf8a4481a23d5260409cb8210ef46fac1a41e9cc5edfe6a4618c9d7bd28cf400fac7818006435fd7cfea00f441dd1bc31af264eca6c77e01150ed28802fe7dd2d5843fff6666839eb01024d8f014;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f633d521c4a06f222470ad422cd3ec99287e2a09f9ae500e4787eab50495ad8286b95ff05d953659b14fac552d6f9ac506508342e4539253bcb33371cd31ae790606518ef6c8f34a4aef4338f2458e783a1f15e8f802c6d6382e720e858e81ae684ca69018a550b9b4fffd25c3b5caad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf54925f910d08308c38236b5877ac846b9b8bb1adc03c76d0f56e353a01087d59081dd2aef504167af79b850c7ead613e3374ece5a93602cb91f577000e62efd96804352ce8e51646632c3102abce1236cedda76825838cc31f12b7d208293edee39e62d35465d787bdfbc9a46075826f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h836afa28658b3892bac01e66c19ced5b853164de21c2d4026bf6ae269deb4835c50c60b600e5056575b1b33920a2f3e2f266f2741f1bbba02c0bc5d0bd6bf2bd9f1d9e88cbbee0e104626d67feb6ada2d6799422056ac5199e22d44b994d632c35c6e6233668c7b64439beb2f02484312;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd38c4b25391e1586af5797f868798a33279d7ed6c2f9f1bf184236068305d51e855cc687c21a32c2300889e1ee7b43a5ce2cafff8d1fe229de3985a12bf2034b925279a86da4ce7ea3eb112b5f610a9e1a932fcde04dc36355e1e156c0424f3e7de95d14bb061a3f91dd13cf85085c699;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46e2f45b231e95a97a0147a0e15b789f08d1ee6c3db481d1811ebcd37b1a0395c66d3e351092ae5b2ca81613935306cedd95de2d8fe4dd0116cb36858ca0cc8e0d9d5593ce1faa52dbae438fc89acc4ac143efe492a0e69cc87685509c540a5465e80cc83a66842e351d202e06a98fd9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2980a46ffaeaa166d739032ea2504f9893674ec7056d2238712c0548fd5ce7d874c94282b9d5c0358db986a97d4a884c1fb7f162c518b456b2d5977b9441bc232fd25bf6e62440976ea206e78821906c15f8ae06bc79ed2365f2d9b188f079c9e3802ac36d02346a8a8df3463ad6886e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83596bf214fcefbeb263d8a6ea89ef7132b148c4be9e1eb87173f0012d63c2b2495cb492bc7e8c787f49886743b98ef8d08e3ac6d5698f82322f076aa1965b7a5d967bcc67317c89ecc9723031ab75ab4af8facd4bef78550ea97159c43c37452abe1b2d4f7ceb6174ba1071e046690ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e04f7ff8d88ccd662eabebfad4146011943c419a5025cc46cee667ef0adbe1adacd172f661e91960d5a21a18d37723595f93e710afcdbe5c891196ea0bab0ef41279fa6cb8ed02c5138dff5a217a7d72f32fac2324cd145fe0667fe4f3a32a6e370edb81ba19afc933a5ea82b548197;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0198b1b48dfa2122da379c3a4ca768c364df6268d7a9fd5a57c72df12240a7aac1eb2fdc2954a69ecf34d47c9cad7314b9cd39553586444946576b06cdefee9df826258d0852e8e7e8d4a80488fd6bd7f687a2413ed819f78df5bd09c8eb7374f658aad72e04f4ce0129784fde27440f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61e3251eb8ea61e93567b2a4e44d8d1c278d990fbe0a1ed67346747c02d81b276c64ac110ca817ca015b8e01feb70a9d81504946f0c88b6fee81e78b8fa190c67fb555a5e1b3fccab798bdeedf947f69119a82ad588852634e4d4cb30ae9d0720bb4719f41eb72eb2eb29732b369a0d6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28dc3ab6217a3d812ab931d39172fabd8dca6bcda85f268d27f9fdd5b9810782a853758da2e7b586444e16ab12a5182535696ad9f07487746cf64b3d0fc82c59c0e213783be9fe361f34e40a07d910a87c0e5ddf44f4b9776f368bdfd38891e27de85e2a4a8d13a42016ef9c2af6c7fe0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8cb0be52cfb7366019f021a97061637705af0070e35800db7481ae66de66ee200a775692dc3dd8cc4b2aa8c87089bc9149c40f3e358a027d45d394a3820b08037c82c95ffca60d4765790af5e3ceb379e846f8b1ba69540cbf0627882e5c127d36f4806a968b2922e85e63d52b797cea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c70ff9e96f2de98fe34c4016a001c591316d9b0a8bf7fd9f70beae90ca03410eb8372b8841ea8cc179637fc8c1bd785c78788dde9dd6d7404dd73a9b6ce4ab3bb97e1caec86d2a91aa97441392a11e528489e0883d92bcfe7b50a96969c847de20c7d10b0a66f1dd11218a79407c38a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h274e60d3756d07b2bff1ee59bbe55f8ebdf3e623ec86d0a2e925f68eb41abee47c4b52b34970cb0ac650e1ffffe52abb81232629f8839d8e330d0cc581bc9ba95e2705f544a4303115cf0b55a3100cb62f8f7c2e1af24364387946a133b3bf25efe8e4ef4e7e65ce674670fe697cdf3fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h956d5b2a9020ba2c542bb4cf56a0e2c1928d2b97a6e83ebd4dea29f620afbce6b86fcd3c130c56f7beb19fce5b0c0d1bda390d7694624931ab88c2db2d41773bc44dfde9b872e549a4bc6ddb79a7bfb9df190946a7edb7133055c314b21be7541ab3bddea1606ec43d34fc1f12795a702;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fce8dc8be4c16f8a3a5d40295b8c35fbbd3ddcd5abaf77f6d1f52681de415202f148a20e320156b54a97ec0010773daceac6a25ae6a6400caec111b9b0e2b1ab43b7c6e89ec43cc4e45833a1c0325137c61ef852ab834404f1eb5df86d29450667b098a6b518353b6ae08faa2b73307e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b809e592015a30d1a9dd1844e715fc73eb219078867dafd5834deb90feba894904cdfd5d7770c239a8e913a302deac4baedaa9c251f704d971ddcb90600131b2efe403c6d26e3eeb83b92608329392c459d6c601ca44d7ce0a86c8f71e6b3e093478719a273414076fa9754c1601851e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h404443b5557d41a0cd549f1dc414f56a76ba091a869f6848a694842dcdeba0667d1ab55f51354687670414c4e4f883df7894a9f7b47ba38dbd8a3dfdd5bcba0a4f359bdf1eb17dda1b3d9d85cab523bdf6bfd332739ad028e412c08a5738cb12cff3c9aea97074da877a55b6fc3d2430a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9324fc946cdcf23f437d5c190a53d344bc09952fbb3d10d6db1d499eba0dc9d72dda4f611665198adf3c5efc0f986c753c2a89bec9c147ae387432865c09ecb0add664f97250077c9ca5cc6d74727bd4c7de9fbb2056841a3fad1a81df1f7b94225f7c158893ac9ab907827e00abacbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca5152ca3adba8892317606c022494d7984782ea7579f4feea6a50b68c0983a05dcbc2808499a142ea138cfcff7beb689867e647c3858499e5e46c0e3cb29237e280c02b883c8fd143d601154ef4054f011b84df7212feb7edb77c238c9a362821b05ca2bc7b0ffdfaa4ba496dfe40b34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc857aba1741962a7662ced879146b5671d2fa904a37899402f6bb0edd30d9585103dfd8286693962353f75c39d90671602026607b83c52c78117ada3d3db688d0e6f2d2562f03626a2c91c760719ffe3ea67f99556c000b53afae0ce34e69ef49465306358f8a5a7e2d7134b4eb9b5881;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h100e5483b2c439d6af98e5567d196d17d1a78112e3dd4fc397fbfe8c0679d3b6461f691d62a1a6ae3cd289571c223189e304caab1dc934d7e0aa1779a0f4a1ef26dd753c8a503419884df6a1181fb69219d3bda506a6a77cc2ad50ed2f8ebc6d544c6f87b8346ed59c1d0a21825330af9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83466060ef00e5ae49a91be3f9e89606e28214a4cf75d6339e7861ad355a0a9f700758db1d1e3999f78b3f6b7896404f9f850536fa3a22c350acae43ad1d210a6549d145c0595f1f2cfcb670b45c89e13ce9abeaecae69be5aa480238c0097c4842c07e064990239468365738d8ec4306;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcba3950c038d40df4401faad66f1e8660a631941d423e22c15146deb9625b256a82a490cc02f24337a494f921e9cc2cd7a69a561b0b6b48e1f5bc7f2a2eea05cafdcc06844f75205afcd6e37043d376f95228c2ca52be8226b01d043bb54bb2b7e20c1a65345ff5aab58eaabb1383169;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84d9df961d1f1c64aa3a0921c4677b7cafd49e6b621513a6da39650d4c27b5ca6259e60c1854800e47a1fe21193bbbe0b86a5cdd0bce1a56dd7333403259dc6bd6ba34ac32e482df5e7c81d4a03555bf18d8e28b6f3e513177b4befdc167bdb7bc95cce69ed70099e84523cd50fd61981;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h539eef8f645869fe29f161547cc48f413941267e42858a8f71afc556e5b70613492b68200245fbe739bcb45feea1226805bca0241052db3109f62c48fef30fdeabca52d83e743d036a26d13f61000fd584b081fe435a9abea74a03744a556380e3165f493ad454246cd2ab61284dc9469;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb78478773ddb0972f88e900303fa3bd52a15ab2f4cf72e07b5bdc49e9517dad2909d5194cfd360927344e5c2a7b7d564facb78c878bfb16650339ce708aab0f3c2fa3782927862c5358d5ba5f44be3c3f4a60c63651cd290b0e8a9cd77abad7d1d2d6cc82304b6f00b762be7a4ff915e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce9a8b39f68c1d64a8f2621cbcbb3d2312ac4d7c45677e07471cad4d7e059b81abdde3a43635bc8dfa49711058a629b96ca0cbeb40b3c57a98caa6816b62684b7346d5999ec9522186aa73f40331eb3da800553a0c66d57da4773bfcd03389994689abbbc4dbb5c5e1350db0d1bf5246d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27684c9f31436060d8d3f5f4796da112a0504fc79695e95069b3196bd5a3232675fdfff93635bccfe0ada9f6f3886036f98f4aeb5ff3e4a41473886edb77c89b83201c98d2c94d4fcb52f8906b767b3a952b745793106398e293f24f37f4f5ce90c378ccc46e6222cb3b40b5e0300461c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71bf25b92fc2a45f6fb21d60b4e2a4400ae00710769311e27cf744ee13a47a3efed8323cb49106436e78a52aea905ea019fca0dc5e99e16a57cc55a97db9675a15d0def9a0a1770f2aefeb2d4a57454178f3e6973bc4786c6a1094b69cb4cbe1a13e9a512fd61f5b5bd3471a83411cea3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h955a0674a3ed6955a8742df86696e760453883414db9568ee02ff45a0128093f5ba704b3be81bb0146ecee06ad6348b3ffd2c059c34f618410498845fc4715e7fbe6244ca5f13bb9eb1f0b599c5f79d0469895d02dc9864bddde4943bc4dfc6fc808462e74eae3a8ead01f77cb257195;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h773336514f6c148b5d0e8ba979727e379400d28ec3f058212663cbbb39bcc47da01885b4c046239da95eef4b73b7415f5e70f3cb0dfeaee547068c528a407f98c6277985aa1abf4b8aec9afa1a7420d9652f00972957b41ecbab8a460b09ff0618f03cf978fca107867f1e1247d294cab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed8b8dd163d312159acc8d507c569168d69bb59f346193c58d9d38cb537bf391c17b5f29a0a6a886ab5cea533f24f5fc3ec5b2ac0b808b758ba9a2320afa3be6cfd43c4f203f214cad4968502e30fb77b53874c6cda0b17bc03a7e562216a0dd8c7c615401c0fb306147695cb8497b7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f1165135daf1f77bc6e3ec8ec545fcd7d578dc90cdd7c38ba00da84fd84179c82c0826b9dd37e5b816433a57e63c58528a06c697cc8c9936d07a1e8a0cca710ab7a3dae72683af47f6bd85b9efb84bd5e55318242e0aefd561e452fad5330179a19de64dc8063bb9ce66c2d59eb997a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37fbb5caf9d5c70dc5b5beeae9aae62da22d60d4ec2136eb8712b93d32e46c5282bda1252d1d33e476e14fbf3131889de57d5ecabd45435538339c89f03e48e2a598d5e7be18345e4d267f14ec1f19be796728af8ba17ab0be872bdae5388cc92d63969d6d66d0b75c36029c405c1063c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b6ff6500fd7f108101f9726cb15bfbc860f04f5d2b0e879b9a8f2b95703ed1a7593e4eaa4f3ee9363c3083cd5e1a1ec6354e7bc925f129a9f5a14feca7d0fdcdfb0b86b07ddedc7b0c3e314c5a4599e786f1bcc0acd9fb8d83565ad3161ee74d008020401322fb1dfdd8962b764af4ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h200e6e975b3c404880ebbf0785c43dc6b08c41d9f7d2793ae90d94e9bd6a472fe9c3f5d8433be7285598f58aefd41c35e1dd1bb4d0da1763886bfc283552c5e96be30e0d85fc8afc2c01f4533ae30d36509ac92ea2399790dd63e1c7faabfe6867ed754f8c7cdfe081ee8e74e4f5c8ad3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24ba79a7d7d6a1751142e9da6ace9d5478047d17ac775cfc442b8267c49085e53b9ddda3d87bf007f261600c46c5a996aa4ad6953b369d1bac928658eded170da1ad9670a66ee0f6e31de0948456bbbb1a9a03b75be4d33ab5f295c12b055e2090cfc273855ac5881085506500ccf1197;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h356dda7dd0eb1f8da388fe95da5d0dabfbc2120c92bcc4bf286ca3336fba00da1b32767951039b2453df06b53d1538d7a94e6011d7d10cb20fc38c300b9c9999cf5f2d93802fc57d972df3458eaac3255f3a571b401884a2c372662b3ef6198b99e626bc02e67af612c2b2e4f5d8b84eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fa5883b36ea27c19bd9940f9fb13fa0c19d63b28c6a88de2d3d0210b2cfe617aafcf41b13e6766902614c4028f54a9591989334af2a6461c4ab55792bde176e4897cdcda547c9185ecf22ff8174b7f6f60382a459fdf6c99955e57443303fa916bde28445e2a523aa79b8258183b8122;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c1a48d3c4d02b7484c56a56e4e9764445d89326a33ea977d831607b8eb9303d17e73725c831c4ff2eb00f571aec6af44148897932904918309fcfab10974426fa204db7c77156ade83b5e516b47b9929c2ec937f967df0ff644cce501dcba7e26a485da0e6a7e58c170bc87e202719d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2afc1ca5250aa20d625aacf0edafcae3e285bc836cd0675d7f4ef71a342da0bb6eef98a53bfa9f5dadb0e45591c89b0a6e3d133f376f467951748e19688ffc88caa2a6131982029047c5dbf2a887e3056ca228731cea0ec1dce2f7de51108f16d112456e6c086031a28943b6cba93788b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8b59a8075e6658d39f9bd5ea4bb32ede4dd438ee6c8418a7c78309eae7d429ff5d6be188155259fefdb5b03348f489428769dcf7f440a3fc0cd9703743d326a62ba1508cb2ee751bf9270030803a0f64bb88dc64525e69da82bd845fb76c2c2d92aaae7225600e611b6bf469a1702c8d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf770a7ae9f23d09ac156ecc0d7b34d5f9ebc14dc0332a479762dd811a66d7a4f0a0185403a7dd50eb59e5ac1d9e7bf8c066047fbcc892a1e48808b0b2fdef0c1bff6847c5de7c4d7166530f139d7d04995473d438a87c4a3572a1ac6f9b5eee53419e852201c3918fed40fb6679a0f7f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a2c1c0210c4f8059d57449711411529ef42dd5c27e0f7cdcb1577d5e662604572b795c79cf2b3d908fc0803d93c09a50a8fa2e726cba67c9cfab55df7f81cc126592a482e0de78f5cd57ac53e051557e0aa8f2f7b26c4308efba12c14611a8637c61802abedf6b9038ff2e524fc65449;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17ce563e623f9caee6d054a85c8eb3000bd785548d1829b478b67c607dd3217666462e3b5406b2bc7ad0ac5ff693f4564ab3680bc22a298872c096eb30ffd727cae1dd7658d7da7ad51b2cf7dbc3c661f79e05e2ebfcfb5ab854d4cfdf309f4ebcb0aa64fc53649979b5e5288b4e2f29f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fe78124d3cf53b25f7f81a2bcf628a5ae2d2c8a4a6cc121f4fb814a4692f0872121a504c8921c78744fb1317df3bb4f9faa563d90eeef8ebd604dc31313d2a8e2d2ba713375698385b20066b94a905db0165f1eefabe7a99ef736ca8659cc76558a48d36860d506ce846c6b5c2f68b80;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35e5d5fac7877a50bde389c210ce09079fec7e48d0223f7b183711bf8b773b7550f0c6d449b7b6fe5563601595d97489bf1130f7825d5b5e385957635dde7358e544a8d738aff7ad8c1e023f46fc9968281b108023afe2576ad9f61299a3e7bad8512a519f399d4822543b39704f9f21e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98a210b877aa7640aae26cc3e05c0301ff037bee2ebfff63ee82204b48f398e3d49880d91ceca538557167a32f849415d3020947d8dde534cb43ba2a8ea93c0e5e38712b80584052fbd85432275ac7a33bd131e0769c1ced0e92a02154d21edbe8bcf554f2c595097ab8d25acea28997f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9778e1e52397486629f59ffcc3fa7bed0b0a8c3821a04368937cb6c754306907b98ffcc4014d3a3844888d09da0355893eaf9d6ee2a7fd9ae16399c94d508f30e24e5e8697c82843c30798b8520a9338b75934edee983eea0fd7d6ed49684e3584414c6970a175284b155913bd18abcc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef66ac17536452ee8658e6cc076efe99acd75b5fe60962bcad51cdfa8c3dad15121fb69fe06903c37f61e0cf135bb333b14f52f86caf1b7486947f74d401e39c4f012ed378e7a1913c8152ae513c83fc6cd031982b6aa3a44e9085e756b2419c36f2061e3af6424bf5ecfd9f6f53b2f22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f2180eb06d300ab1a8372c9ed2755472359cf13a5740b16a8b6b7f623fc361db048d9e77db5688ce75b58e0258d34769dd5cedb8acca480ca2b7e35ca1183e93c582d3056f82eb96cd9e51ee57fa6ce7a88d94402ca9abc328164c8ad46e5c5cf11152545d7788c4b409855314d22b3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99f023925e335934dbea2ea44c1eaf0b193b95f913bbdd1bcf5df223f23eadde3899ccb91aa15e72c7c2c9b497fae3beab05a5e014344cc9947d7e7ba922da85530774dd1c2d99f54d9b67445eb165a5a37c373148f08beef267d8bea0ab395e36ff8e6bffb4ee916aeb800143b855282;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95ac6bc48317fb13da0dd842f82f47c32755b49355469a66991bdd34658156b1de91d301984f4dea9fe3482204f86428120c785122d83d7f20e9520baf31dc21323cc79059bc95463220fe4b63abc97e8847bd16549f4ad9911793f472ce08e48e8fa62bf89f98c9a56513fd4c21cd54c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a78c6e5a3c548237e778bb6dda59b32bf1295db4268f8e54610ae95de87ee5a017276f38dc320705274ce66f2c165e5030a16decef27828e624fdcf5fbc35d971a831391fef5d244b9315776252cf3d7904523e23fe925da65669240b4cc386042362f7034fb66b296c427415d7597bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcab41e2ed453eb2d8f00ccebdcb6dff27601eda834e76d2160c944d09caf2778abfc592cc3105f03c3955e7e1d3923a51a067b395de23bceb912e035fe4cb84fa2770e40e9f32deb44aeae56d391c19d7cacadfd09966843da2e6710e20bbc02ed0d98e4a4935706865929a7cf3d4f50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b02023c90d062ba8038e92b01abf667ccdbfde8c833aeb53b21d1032279d6f0200ae81903e92e02f20763d76bfeed7bab0bfbd4899cdf91e33a6cd350c7bb3c741731fa75ac07d0353bad5a3cb4745319ededd3c2058f77572f7d14c2662d3c63c38d456425e2c8d7ff0e895648cbd47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f7eff285ec46e4bfe4db371eafeb676b6c1b7e5747fc96ae04f2a81890963f30027203d4ee733e098647a7e9f80fe1055e2d76eaa72dcbecaae86f032b40e084f5ccc38218fac8a28f20818f3305e81e692c736e0a5b2f8becc8936c5ab4012341ca79ef08730d71b93cdd65b4f73710;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4305c61d1d8d42f32091126b3ace7380d246626da81500c0a1170c5622892650e561d3c4cccb6a8317749145ca4e77e285f74e7f99fc7335dfde1e210381e9dd01f897b11da78d03d59d95db2473cbbf7d22b04bface22ef8466941970e559fbbe1d914c112dc675392d9e1dd7870e89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h506cb0c46867892dcf00c955e81b64f558fb556e12d462b443e92bfae07984105ec13975690f687385fc546d8421c0c1856eb3c62543e73449c942e6121f81d6a4b5376de09508f8aafb1bb852fc06bb9e85dbd0e61f4d957d682337115042445b56dce52ef42bd132171d54eb16b4fb9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h186f89dbc6577eea8a1dfa4ab60327a0167499ebc201148a7076fdc7fb566d7cc66432a9ffad8f61f8d05ac3ccca985224df1079805f9693ec1effddc099050b850d00189ad80c8166d12167968c3c5340cd1f3da1031b2097d6b98b3bde73ef44bfeea5f401cafb7fd126a4d71eb4816;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf946f0cf57f036aec01eb0c8e0fc21a2be6f702abb87bcd4ded502dffc1260dd072cd9dfa0671384e0054f1795fbedc178bab7545e0e944577b52d6371b9cf77385b6ac7bd605bfdc6b69aaf4fa0db4e51ea61d52c3e33ba691c197261f7706ff0a6e614a7a47ce2275f0fa27528e613d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'headb1e2c872c6db7fcbed0688604e50b3278042e773e62c6e01a977d54e7a4978098b41dfdb768820cc813f3585eaaa4bb9b2ebafeb4db4a40e177d0eb778bf8ccf949abad8acd14c518cd7c4a107e17a06408fed0c36b8a3ff09bcd009389b5ca34f33475d2bc2f22b2c2ce8806a3a00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b139516d133089a4863e67f3361c34bf893c4968517636fab7ebbdb40cb26b79b497bcb087504a1d28db2a7bbd138b4e4330c0fcb443e14004b518130348a9632ab2433e63c954dcf8429406fcb3dc55b0961280da6634374b4b7eb4ed0d33641b2adf8f6da7a84a56827193bfb01c13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46af2a4b51a9b1fcbd3c0ed254fa1c36be1d0a9ae260cb512d94600b69f6dd8b19c31300d796d013f6f65c83b9f4ef21dab4391c83dbdca65ac0f7770fb9fada96c4498c71694a242de56b4f8e86e57e1ec03d7fa762842de02e22e89c42e8dd926b98d0818a750e65b789a55ca32d90c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2a9f55019c347d65a8b79825e9ac131ac752748f4ad2ffd0a0e6ee82744ccdd2a1b0c01a36c80d3e87dd79b39ec6dd8aeeab71fda5c5c4ce141b803e0fe5f66c915adcd5d81705e9bc7f9e9ca0e5d6dfd7c215b03a3142f283ce2b6f86ebb357996833cd29f7721b23a4f0b0b07aba4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83ba3cc2c615d5298fd12068a411f30173370ac341d2114676818c0a8391540ec523708fa70d703a9a028fd06e03b01de61d1e3101abb90c832587973ba4ebdc263e71dc5c95093714815817da9b29d713a4a07f92010679867812145de699ed64a49b6dfbd5fe0cf3ece35222866cdbe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84f492b7bad74cd00dcf983023c0d61df7ad9421e5e0235ceb16ec58cf0d4431d2608bbe0c404aedf4cb1908ebdb3f359c46aa5ccaf715b72c4799a6fc360ecfc97a5f8ecf0449555c198a1a0829b7643aab07f92c5c50727426921e98402aa77e6594fc8402856f7708b29bf3a3b7b3d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36f705fdd2381474a532f437d1a2c94123f8904a42132b69f4585e18ccbe7a6bdb7f9ae7e52fa0736cbcbfcb009028883526a7f3bc3f8ea5915b30421db72256297659a3366f4868a01df22feae0373e6b3bb867f9a9018e7bdb937080b724a747651817809133c7faf55f2bdf5b04e4b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4510775cab22b4c877b21010e374632a99ef5ceb6b52574efd60e713c54edea69e9aaab46c4641fcd3a5ec38899733b04fd8bf11d6d4e7d4dafc3836930c05d3bb4f8218d5bef0543711e7de45495322ee4025f8953fad17b846b2ccf6ccd9443e562b6ee88e0acb793eae287cfd379ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1290d8fc331c89746d1fa45fb686aadc45a07bb2644a3e2e0d72db0ccd67248aebd1cb7b28417dcc0a430c3c322cec34d1fbad93cc7a26e5bdda38b4f8dc23af71f8efb41e3609d8ecbfad88399e3172ca9f638398338387fd6f85e53df6bfb4286b52ad86cfbb89f7766f35946d6c233;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8be87d914d84eea2d66654bc8ae5bb80321be1206ed4bf9f2e547d452550fd1d1f4f20a4490fbd5546dbf998429ee563d8cd3c79400ed20345bc100edb738f3e5b5460700fbca7971518d051505de62ec80f8e204c6275735cb6238041e3d91f03a61591d35ec6a5ceebb0aca09a8cdce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h738aa6fe2ace2baa03e4bd5e9e9ef67a9ac75320dacd0297efc5ec9fd8666ca6d7bbe98c9e783988eee50c50bedede8371760d73d30ac3679e5b20e95dafc9baef0703c415d53a26c6ca3c5537db24f9b8e5ecaf9c304b5413ff89e0b4ee0959eb3594af1255a9cbc8d33cbdcf735391b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haea81693b37e22992dc7a8d1099fa211873714f87b913f2494936592796e50c050d8d095928ec5a19acf4e20766da02b8ef6f01d79ef275fbe7d5566bfdf6413bf97320e689da6c227b76d1c6ecb9a0a32f7b8d5a97cdbfa366610aa2942b8e1a34a0cdc54c2372dfc082519f07a8f8cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89cd169fc7e9a3686308fa00f13351dad2857a2f1552563af553e7e27da8fd0352ddcd40bb8e83ea5eff159f433aaade23365e8200b44e62cfcc61793940fea36a026ef252139675102e4fc27af87f87733c6418156b2939710d87b6887666008462f1d9e88a25d7a6e90fc3fba3d67b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd71463cf4bb9a694e66384d2429666c698f6ab769b8a2c4abb4a8a377eb914259f386e085b94439d8a0d817fc9995e5503c7104d5fa02db7fb6473082dc3af8a782e1750b6ca48abd4f08589d1f642a28c14a9cd2d8bdcddc63c056dff43165dc2edd534bc29713f743930fe61db8a215;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fbee5671487ed6f9b8cf407efb4f162bbc86d116306392576a61cfb768474a67205ed5556803fcacc371bb2b3da852cd08960da408cdb0af379a089460488b8ce2c2561b9a64cec1be418c81db99d10162b0e1367b5340fc5dcb7cc0fdeea69fbdeb6465cfb7ef9afc8621a0eaaa840d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c13f3ca41a151b8fc986fb9e509dcfcbcbdd473f5be26810fdc64c7859ad706d35b31bf0fcdbf81fa4c4d61254c9aba4f75e17dd6209267765b45adefce485ec6bf6b52dbd06a5d26be262da947deb090fe158bab819d28b5c60df5ed2db9524590f48f89a7c105ac2764fdded4ed398;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h508e69cd55d8cf016f3e7ef09063e4280c235bdbf53c7d85e4125fedea2ee3d56fb82d79743b8295c8089c2b5cb9cc32af91b517f411e0fbddfcf58650b221da3bbfffe0cf2e5388bd665e20b5f00240d603bab92c1f8222a9c0c683d54b057bd1f2bf9e36c873cc384a469fc91cd5351;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5419511ea9dafaaa6ac3e5e5cbb6c36ba399badd8baf1012fe763645b36caceb2ff62392e47e935f7fbba30a71ea2905a7a9bae8605ba37ed96044647faadf6ae907470e3279ad4b5eec437cde57a2d9127984992f3f32c2a0dfdcb551473c70ba93a2f6afd3ce34e25dc942b79dff8a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15a0c032777389b5997a5b856f69f98d8b9f28eb9574c3f5c60dd3ef21dc02e81a49d6b1a52e303e14a0bd691b0972d48e41584e0d62cb3f7ca796ca073735b570fa0197fde0d9b9fccb4ddfd26c1b2752616cfdeed992513363a8089848f9ba797283be8d5618ae6a0f4fdc5ac11e2cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc6fceb39e2c37b0d14db3fdfea57baa5f564202c1b6fb29a18457b1fb82f201cd91f200ff604ef9804641a5bd8cad72c6b195cdef1974b1ed0490299804f9f3afa0b845fa7ad7649c8c399106d67343966d7114d9105ae5872da353ad62aa5ed79e2712f5003002d460f61c531522f44;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf455e83d8214b4c1bcceb8f6309c0f29bab7b568706ba4fa2635ddfc121421beedacabce4e7d05157a362d300516a955e4be72bc223eb174d6badfa3f731dd1bfc3e01970bfe7ed4da04647711d76a89b4e2acb31d24368c762817d32f897db013c55ef8ce2c77b6a624bb358883108e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ed5aac60c8426f7e519dcc3cfc6ad88a0164466652cd68b8b67b5e9e1bc9bf8035367107baa8ba443e0b33f55535bce6b1c51320f017708179bfa48f31e50b31094b2926c5bead75a6e6a5d8f1bc513e8bf301352811f0d1ad2a574fdef2fbbcd096a30c4cbc17628d095da834671a64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10545144c0ee4cbd0fdfa23b3624f493115858f56a2bd09390827f4b0c4a7c10c4909a5a4316b38a7a98b96a4a0a11fa1533ce9fe0eec65cacb2697016144548fa5de907ec1b28b64e23adcb2e9ed3855876f5509e6858fe66ba9517cdac266c1112c8500ce09c123b768b0fe2147461c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd6556c0b3abe569047d1f16243839afd8a55485905e784536d748a85aa688ce5dd6a05bee2f73efb3fec81f129ed2495a432fcce533acf449dd421784df777212b4b053bac9ddf127c5926d7801b43ed1d4b437ec101aeb65b34f0bebcc8882537b797b744274a9d0a0c6fe6b482232a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he46a774a03e3cb16f6bbfbb03b153e6793ddc791aad60bb66776bfd6ee24c760aa76b7274865aa48bafb1db9a5ac2ae97c0bb24718a20cff4855490836cb94241749a75e1446a5d5dae905d26786610a9552bfdd9db9934c67db0434cf712a45a0ce1f49e66a0751da378b243c1e32281;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8ae19f6d32beb6926857effa23d37a0df182a87939c871691b028ac945f521ac1f0008de54446e6fb4c680d71f090048c46ace6839a51d1623fd0a94b7a3d20e43ec26766a5d8698858672cbeb5c430adc2d7714ea5576638e9e3bdb45ebe1f755cae543be6b143d1e546fc3443acef3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a8aeeb0c10efa8e4e1d76f7e4f302408cdd51580bd711b0c24705c21a937048e226e1cda4282fb6c9d58354d97e2330fefa735c83021c6d8e7f47a48142e2780425c65fe86467cbde7842f8d42093c8f9e176954e20e2ad3554c93a9bbc69814d6dbbbbd6cd8c9147992a45d19f81331;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a571b48ca9be8b143f0ef40c7debdd41bd289d02c43668873d6b640557d6cb8b5c79528bd7820a575484892fb370c45f5d953c9bde87a1af51b323e0f80efbf5bd3a1aec17b93c5ad4777a618812eeed0e33b5edbf2079e59f1a61704daa51acdbd6deca19dc80435aa5a7dd3f59fc20;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6266b0aee2cbd0373db238d3165d7448612fe906220a1eb401adf7f0fad22730347d90dd83a614a0bc179c4521bd97bec4e5e7b7520254d04616395103f1a3eb75509ef8a1bff8980b31b208358d3cef41ea78dcfb4d9abf0c7208946ddd47f0c84839cd6e264e76e948bc5324a5d9ea7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8d87b60da79b96823736b8a2358d32ef861eec775db6cecd3cb0c90ebcf98e34531ad6d5a5055bcf7a5fcabbd8c2d3649c937b41a11553fe6161a0f72a44607117bf58e241d923c60d35f8ea2db4898cd06b0e8494da8b7f2aea88af803c9b1d25e21e541fcad0948663298869760b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha171270096cccd2af2c21f707d24bd2ad89d324607042774a04458f1a574009d851778b4ec29dc9fe4b87a246e9d012681b33480d462523f5f4a1042c987b78cfcbb594bff28004095c118bbab3266ae52996690f94922de0660d15244fb209b42b4f6b2915b25313afcbd20de69abb61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ccc65217300d37db5613197452976bd8dc3fbfc9dccd7ab6239f269c9e04c2f033d61c72d709ef750f30e544de0805a9034138ef5c6497bcd6d23be9d3a62fb3dee2b3b130f4d7675fd954a4cfc80cc07a0aa22526e5a314bc33452c5d8b159ac3057f9578e2884a0e076f23aa9a6db2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aa8ab879d4946642f0730de02abe602aedff12a9e5486b3229f4c63374ba07ad54a2779ce2532e66e197f6cd6e6c06dbe5084e9f40cbd566465121cca9f47e843ee18ba79751d169d79e9c7898c77eadce83c5a2286157ed8e32773dce7ed1f53cc308093e377e770e259b917c124761;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6975c36aedf448bf0d5da4418be6d4b76568056e64be1492343779742ffc57579f73fdeb7baaa2b05a00389354df5f142897bbfb9ba1d4caaff2d8f8c3e510d21e77b5ae4bc500ad40b4d88f1b3bfdb8dac47f455664fe81d1e48c985fa1da0dcfad24c247f7da7f7584f625556830ee2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3e70c59a79b32fbdecc26f9e45b85ff6bdbaaf67743b0b2e13b8fe321f6acf48c9dd1d5af7c172ab5cd257e332eaad879d31b9ca99d072dd3af97485c7c4d54165e83798d49d26f19c66c768c65170c6411ad57076261bd619ef37026c6dbb7df42893876e86ba01332e3f4cea9859aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c13ef061f99bc7d7b4cf6e85d31c99540db1b05eab37b30f67b212ff4abbbb0eac97803f83dccd292cd3146cc0fac946dccc4cde777d30d24a4306c3e2db09c5428b3ff4df2e2cd89a9dd3c4058e3198126448e31c5ff6a54124afa63f7bb135c08195f14ca49e91c1d5dec3292f4ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h144db876184e8b1e3fe012ff2d6767f976cfbba32b2f020340a2203972ddf578b77eb06499f8ce344e9aaaedc7ad7d7c70758a454668ee6adb10f0758cb7a20ce3176793f7e69e2b15ca85359a2e105ede8172b279c49fa0bdc972c27970599979a41e00093d404a7e20acb3ae4c593b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haddfe5a6d6213fc91b3089fd45f6e52dc0c349c80f2e7a0411d67b09a57fe1b0b50226887abc21aafdce8508402f9467fa64d7a69b16b6185010dbb683d3850279f1786e4ad6d7abc00e2f2157e1cce584ecf6d608532700273ed2049f05bd792d4a12173ac88a7ab3feadcba33bd1290;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43d8e181b549432f6606ee4d3f05265962d720385d1cd4ea49f80cb4782001f5cce3a9314d37b5bd7a9a025ebf3a96f66b2b0478fc7223547169c00b7c14796e940f99571b6aaccf25e886c90a7ca9bc3451b83250243bef09c4021dc54848e1d852ff1e7ede2018728425b040b57a664;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23994e171ebf8641770dcebc8f05844cf67140266caa9b2f1e9aacc8322da5ccd38890eebd5c8d5745f49971144cf8d5057d3d53b9eeca34674a5c3a0f8adf556e60ae8e1a75cc12f651a3d9af913ff7a8ff9494ae8db72900dd449c2cb3e45f80f2422a443352fc1b4451d421a2c14cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3301a5b515bcb27e2170d73c8089656f79378d1dd6dfadd115b2dc4e7830644c8ac99b5b3de976d82e87c2a71fc33139c1d818c2e3bc3f604435294f0e21f0111ba210c16c1b28a3de686dcd2842446586b688eb186231f442a2060ae77eb08deadda2d5fe2216833ea9f8b80bc7ac867;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfe48baf33b0c35184a7cae24295cb94a65f057711fad7c4dc4971f627c44d2e2b022c2937fefa0babbb1d74bcf19dc5ad504cfd4c163804500d5bfb9ba8728d1966f327057382a188f37d57bebf1b58ba62f26878aa7a2737af9e303eb27c66c1211c575d20988ae21f94c13551aca32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h289d4c698c1db1128793539cf2a39089701018e161d2ee1e56710cb87b04aac278b67e1b3ea7ab3bca339ed26e2e3c1a1d54cbebe60c167875626c3537117110b9f57f9a5d28d763e0afefea67d2577132ed6a49b6176b97d91ca910469258626f8137bbe4b5eddab5e88c18265e7d22c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59a4ea7d6bec5120cccab188147226e4576e0705993492f82a672e30d7c0a9ab3cd3341860e284a75020729329845e509bfad56a78f13a8236a6ab4fbaca483de4837f2d22e60bb3ff87100d4e8f4b75cbb3023b62eef57d0a84ce17e6d0b1c40c1b00a81e77ec8100062bffae0255846;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49a07fb7d074f07f3db8bb7ba0685e0635705f609eddd455ab147d42645344949f96736d810ec229d6e9e781149e48722b4f8b72b3491ed18a57034ff3264c84b052236ed4fbf1c5d8a94ee6e4efd535086df4213ed92a5aff66f2401a0bae010157d0b0719527fcb99495e204b49e337;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he295dd977af7260348423bdc6b4fdc1be2504571251aad763bfbd4aa904d09e7edbf6304cffe89f2450206bd6e2ab438ba2828bdaa5390a5ba68bc7e36fa1df82838c2ae155a5f4cc5d9c269dcf68548da1e3938c16e91cecafdd7ba113b2455ab7828722f3efd161ee028cdba011e8ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e258948523680ebd1de00d2f77e0235d033cf21e40714e53a90e82ae32420dad032699317491629d364a692e9ede71bf70b80a9dcd0d2e80105bc442c3459be38e50aba068c65502ea196a0eaba2aefa9f5421f98676c2d5490b9e372d4ff70c6b1fca0e2f252e3d560ae701cd947907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf38ed829580fd22eb426b0e67e480d3e86fc5426ba2b09b6eeecfc07958e9f5041b42ad85148255cf4481adcee4aec68cde5a3af030c5c2a3bb4635291b4807f4840c82dbd95b4157997ab8262df188e0d6e4234e6cfc8ecc86262cdb96f8ab5951fa7727fcfb32c1e0f0e7a4c7cf1b58;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2b8436593cfb49ccd96651ca720d09659fd6ed085c32aaa1d325a7c11f263e54de85294cb3514d53fff44e8260584b435a46f78264e4fbbbbfc76f9ff0272ea72d825669fbcf493a906da0f60b2bd0d2cdf90cfd96e2073e9178e36ca5d124b3d27cfc31004cffdd20b90b9c442ac0d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55190bb467a8625ad353d2965e506fd6a3d98211254545c2292f3fcd9484278220d76edc5d0bbeaa16f8c55de044ae79f9d243a322faf6abef29e737b870dcb18dbbb7c1642eccb0d58733c763401ce0f26c69a411db8900b54a03b95a94a49fe1af57d99ab0f6cd3f5a1006477986cc7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79ed7193d6d4742a42a140667fbeab505325bae64444634a7b6249317d9d63b5c2d17655b466aed571fbbde20adf997462d4709cde14a780c175f61673c0393448d03f94b0aba980248dbc00b91dfa0cf33989151b5b82a9ee2e864b812b1f71a1f0dfea5f1db8bb66f32eadfba535f73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d9c0da3a9bd83430b50f297fcef0d7da4f86556a955e8df351ad36f34f0055a8059cd2c360ff2e20175c6fe58551d99ccb1fd200cbdf31275e8c7d1a57e1503a8e0d20febfdedeb4327d2d1e4ba6aeafa646eba6c16ce02434ffe7fbe76999b6ce8df7402d03a43dab925528a6da982a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6cc8f1b6ec54861fa5781ee5f3abebbd6d6d7d36202176370d3e05b45f32d3986660dd82c7c9ecb38eb65c1b8bbb4c670ba6314a1fe018692861eb27226320fa3b8d32eb79a0263fd0658e047e9ce1cad538598fbd808fb8e092b36fd9c2a60eb2c84968bac6070db48329f909cf0f74;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h824398488038b5e67370c866d1c2e74139c08881e4f23ae258c3d826b310a81900cf331c03bcb777c98095faf547b46ef81ccc7e3de1374c287f77b6ae28a8f5b1184d7ac614d440e3170d2a69244a45d1f2beeaf915d545b46f74d5ed7dfbf3f1a01cb0842722cd0474c1ed45a4b9f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b7d1e4c099f48c3394d256a79ccad027bc7eab9a94f906b5905c26898a641f7e006c1e1aa7afd1a3bec0ad79dbd0d0142c906ab242deb93935e1999d8f97cd412f6ec8dc3851a4842f11caae6f037636493b85a52589b4475169c8ec781e087ef0371af06dca4b287cbf0d40835a528;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaab3c65ee59b5ee9d18b41032ca209ae95b546b46f3ca68304f588ccfa691f12a6d758bdf3cb8487d32b3fa531c906feee268c5465571035d0658bb855c51714658e4f2fec7f618ad9e807c5b41d7c2294eaf3a784724ee930fb6d22d8c8d3612d2ce5900f909060c9173db84e48fb26;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed2f64ca25f2ab6e58b1ebbbf45b4e5e6181be5cf2376e168a529746fd114fb5a350a20075914501baef545f0ee6ccfc3dade567452b69f9c4d9aa56367ec71a40b2c1d391d759ce7f7ded2b81ceb951e57013e35c90909deff9e9ee0c83247824defe5228c49661b86a4ec7308018a2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61dbfe4c6b77322dcc5145630fcd0a489183ef746145eb9e986bb83b82704d5b8d4f5cd9cd258884ab381c389c8f26cf097322f002141eb22d017593e4481bb8b5bf896f2efbe50f74ac120116a4fe694ebb41c418758b08ababbdbff90996e32dfb95c846ee92fc59ec8024083a5a9e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h183c40080d856a6d4fe8efd10b8bdd3e7f0d5023992c38e2b348978548e66e24c866ec19715341a5d22a1ce3c8541fb662af6f1a0219ec20a1e58b604a6879a3dc5f02b483dc537cd9aea04ff28a08e4f373a0f56f79f49777aebc19be56d2e74f0e63f7ba125ed3c1ee194d3178279dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5d820d89f17f0435c6ceb208d45aff8d88bfe4482f674def9fe4bcfbcc23ff329c860161d0951388b9e6e0bd605c8d9de08cffc49041da27ff1c28c4bda8d8b3f14b66c9d677233cae02de5de4086d9bd43d8c6127f6a33c5e481ffab1fafa82e7b53a6a71cd07b5fb064770a93a7713;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d9ec5e7ae77c76bd12c704ae9fc7cb8c08ac14a1e4c83b9cf38f8d3ecbf4ed2d5c843b264c3731c6a856e723588834330b8bea6ab190691628b72410ee16fab25d9e94247cf83276ffa3a91477317d1e2137963a5fc341870188636e7a4aa928e204526a742bc1c9e751f16e913f372e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf20322dbe05acdcd216cab91f95b54993b026839b5da88a9e042c4797257cac56063b6c091a555d67c56e58688f02cbd62e952ef985eecbc4235a1091f1b8e0a896744764f38961c3adf533f732c5275f82a3cbad18dd46a932674e51591e25e80ed62f32a4c15a6696d922a1ced13c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4df6bc20c27d325b7bd78c1abd1996bf9bc9ae866ce7979cb7cb90f5354e4be92821d964635b1e1b973b212ecd3543b8b7f9281e7d2b72a353326f38518be33be3b55549d00d330a47f7e38a315e6a3136471fc763eb695a2c0709b43e6cf6d3196f5fdacc7e1a79475f4650c6c9dd0f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4cbcf74289d99cb50799c6390953877fbebe2fdbab7f5a1c71ccbf101e6ebb7a747cc82b35f89cb5bd39e3f7c433fc8bad0f802e9cc92ca79389876396842675092fd9d47f86cf2061cf55d1e9b2ccd349452d532a3fd884b4cd9e380dda1baf871ea250dd2149ae20fc475daf49119;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h326d8e56079e5fb36f690f0aa0b3061446f443b168905a90293885628ac33883a406bb72b40a939b6dbe8e04706292a27839f6a3cd52388948f5c28f0235ac02f9d7606d76d3a0c40a4d589284b484b4709444368541293efc31896910c215c35499b0ff98f19fb3104ee6091792be569;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d59114a1d8b89e0e43996078e8293d4396ad20152674eee43077ad61479d193253d25b4e1dac84116333ce6e84ee02840f67dc2813a1ddb27877bbcdc3e3c3b3c5ebd187f39a0fc43458be4818d7819b44a90c429c522495ce684cce18571ce88156f6471697f7ac5d373333a55890cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h379e4fe435cbb251cf7086d930a4d36bd3d0079fee35bde0b4fea3b51a3f7ca3a5fe22b6d73ebc69497e04810085a05ab6255fcac21fb613e4f47dd323843f13d8e51f56890955d83eb4d1a5de696ed83e2ee358d3147b310cdcf1371c8f639b32f2e6fba199eb934c83c584b7b4ea8b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8e30bee9e5896e6f5195cf652698bae22abb550a5adc07e2bca8cd99e5f5e1929d85deb6f62d413a89cfe7b8fe14a80af44bcbb3e92c943b4d2165eaf15b4886ea30bd9e18bc1a1fbff451ed1c3040002ceb0b3ffead24e88e9c0f5300ae8fd8798afc96e183f9d4f91d2d61876a4af;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbf55a96e4ae94545ac9330be9ed6e7aede485061391189f5091909a4714fa1f5d3df324ffe2aaa2e1d2647e65063d3f24ee45648c069e618d1199b942bcf1c2c2f93aceeb4532ab1e95a82811f5eadbd2f12835d387be3e23fea030c3f9bbf980abc5f973a4690d248243bcdd77770ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3f0a399afd70b9cb5472a2c9d31f6b9edb7a7d87b81ccba1f58dde221249dda69bf183b2db157c15e2925fd3f94d02ed7d2ac84888857778ffc0eacc8901fa47c14ba71e9a7976948f62fc82635afdb4b7347da188dbd0ff31a162fb597625e8b0fc6d15c0bc771845d408e93c4cff92;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h696ce888b171be49f1a95489f9a8ce34a8360e8e33a8fbf39c2d7f07cd62cf321b59869ceadf96a9dabb434cc86b222effa8ec1f0427208b04a729b4369aad1913a8e57e788f0584c076cca818fa90d6c096234dd6088de0694a219ca3e44600ac7d9ae25f194ae915f3f6df23bb96745;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b2bb79aad9cb0099bf4a17a7b2c06980253fa09ed98b07cc6b0114891bf916d18e383abaef623ee29bae9546d140b27c45999862fb6c0bcc470d651bb5e4764eb74d3703e2efc5ebcabecb0e94272dc33fb9d5802775799ba4b3cdfaebf98a3f36930bb7400a724b290fb5d830da8138;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1043e659a6a66ce366cc98a5c902dc55e5a915d0a8887cd5b3b9893d68508c236c4cbe97114b2f32cf40fbba11fef01d0297fdf7a755bf32100fc6e6b5cd853895a42f28e578d0041f82336cf8e4d94007b7a6e545fb7122aac4c39118557a62702366ff3d93413c71ce9b2955f6d23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f62a04e1e7a3de3c50cb6a6c3afce0306de9a97bc62353d9c9ce4a12d79173f95822c822d5aff10fd993e28002975e6787bc41fb109ec58dc33a3357d92d4b0e40a3b27d46787858bafab75c1398b1be3fb860feeef539657bfcc8745d1d29f9c0cbd89f4e314fb081ee69ebb0cf661e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h358a2a48526503cbb17be65ce93e4f71d1664fceb599f9e96c5a23ee701de2badad85a1d2ce6c7a7fce3795ced90829efaa8f9317d1d8ba83a2baba89ada47674c8580e1cd99ead24db4c08ec503a54b6b5f2ffacae6d9f12b05542c2136bcca21acb64f2b4d7fa494f06847dc0e57e1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbec1d4e44f2444bf398e786796c8464b1542d4084e1025789a1bf43baae70a1af94b378aaeb88fd70bdd186370cdbf91e573291f18d03229b00eb9b56191aaeaf289f4635663ce4d241da3f8a2b11b25fca1d4b800f5c5b79161404b8832ea4b117668a4bf749bedf4aaa27321ac55c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34232d2f8f8aaedb6b3f8ed743a8a14490994e88b6295961f73bc27a8c5d7ee04f2ef8082baa6290e4472d26b31c1211c57301939f72be4e0963cba90547735e4ea11cdd91afe5e99aff350504b94fe0c2f26477654c5b742791b0d7ad2e4cfeb49538d23477c1ebf578c44e5d96400b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2270274884bd6a6f8f9ef873c220ed7da493ece569178a893c551b798493e5e1ac2dcf1f89f7b3566f19f69783e8cf883fd8665b3b6db30cfd046610d3959f1a9755a6f050f441a03c0cb86b5558522aacf60109c7694beb11a38d555bd533e6c29da0edab6d2b90aa31b05f00434a362;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2b605a18d8612ec1a8a91bce459c388844bafa1de11d999830a3dcc039befb930b45bb5e1ff02d549f14cd5b84928b5854fa3bd814115371037ed41ca80d7b71b3681a2cea342d66b055a7d8febaa4f618b615595ca16bbd0fa8b412989bf2a5a749acca04d7feb4208628249ccec947;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1144ee27ac9a7d40b06dbc201cbb000bf51a7be4c3415d478bfd0530d0ae520022fb6bec46bbcf7f926a507a54b041bac6c99deb6e8b54fedc8f4d49fd62c3c1a68ed0390e94b9c3b933fce2c579e3ce3815845136c6ebbe46558d53799b4d033928801c4334d66c2ccce8700a677550;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b6e77230f4f03c90c8147312d3f53c3a68f04911283c9726bcf50415d984b4e320273e6a1913977b3f529e88891a4e0d788dfed510d0e5399d315a98ce80ca2fd26e61197b3af7cf1ecd4324156a09cc0266d4a48f74dece3d3f441111566cfa71e08e365840708414ae475e3a03131b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce2082eb7399363755625783f973f4effbe55440b540a6ab18a7d37aacc717a19cca33ef1aa8d0e9940851fb2f596269b3697108a82ec58ce7d00bb9fdc5b898baf1e8a1bcd239da93538abe68cc023cdd4f2eedd48c8d70551e1ac7d584f34476967b6c678362ddff38a00a965409a40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca393d53dd60d873deec6d3c06d8099883fc5b7b407a7b9db0db722bcb617f2fc88b8d457e4531fc54f8f03bbb61325bafc1b73dc6a39713c80d29fefaec943e2295b39f3070ccab695075a1bf44e1c331f51cd18cf3bac6b4129f610eaa9a1d891e78cf40bc557ca486f4f6c780f7490;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12e3f9b10344d363ef1464978943e76c0ebf3c924e427a08d4f0c88c8bb25e63869e0543140b00d3366f1bdf37a9c8610778a4021ac19eea269214dda295fa795b5741a581bad4d3430a23c250e676cb6ce346d4f8d78efc7219e82e210816ba31dc28fc3f314c769b8fe43daa78fbf71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f3a92fd12894f6fa4131e4011d3aa78af8353261f235f50acbf07ef6c02dea1afa945598beb914482570fce3c424de20efee0025ec9c48620d11329860f73ff21485321b0e9cdd90185b9c4c27e478c8df6a502ce899653ef8e8c009b7bbb91ccfe54f5ab8d8c351dfafb0ced43b3868;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29f8896d953a1d4773a5811d015edcd20ef93b1ccd2e76e39d5e38afb30239c2a24c94a4c9b52773a4c315f82b921e8ac23a9588ef609929750dd212c9d8a3168191a151f1412c71b82a7d6c2858d6987d14c310e600eb2727a4697f7e21c0e04d589c7d6ae7efb5f7c37ca917cc25719;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56e6567dd5632fea3200dca299cc9e851ef7587204feb58239a83ba683e914be93f71213e24de4228e97df7dc91f8f95546eff78aea4a655b8eb0e784ca80d4f95618d5b0b0955912f0fcf360b4b4c80530e4287b5e55ca4d17286eeea94d29dc355d94587c45ea978121f1360100c4c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd25c1bed498d706f67845d888712d8e67227cf66e7e16cbca192aea58b2ebdbd1e5c26144113721cae267f4b8e70bbcb5bc7466041d7a57609e6ce4aaada49bf14e5341bc5a4e24a62f684d6b927164180373c25bd041c47f77a6004caea647a715ce15e3104707b8731ce108e26c762;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc03077e3dfd06b893717714de46516515e39bd8774d6a12b9a856ec7cb02b5d136f12842b518393e591dd742b54f2addc18617162222ef5a719d5239b4df73e19ef0bddaa2ba074af9a547e445a41e696ce30673a3f6ba76627c75ffc09118aa7f5a211da69f0c8d3b138efb450fc454;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf49dcecaa1a1f15fc022e3cca6efde8bd72f1320f3d27ae3ca5909a44874b789c58da8482222588f65d05cbd8ef771fceb7d155f63caff6b89c74783adbcef473dcb0609e03939246a4970322e09788e29ff79a414e8112c8149098ff1433fe9d7ad4909553da1fcc625310a2cc4558f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43be7443cb816fac460e8ba7cb2a7e90d3c9d36114a2ac57f51c3370c068c143ef13f2313ae009df85f2e932c5d5758def544af2489aafcc6918c4c79319d3ee6d5c149565a0db15367d26142d56d73e90e5c467e210904e6f9991fa5cd752bae2d316d1834a9bd42cf90732930f59280;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91610da200c2494d66925055a2a4ab5d9aedba20da7fc5ceba8253f2b328e3b5e14086edbff00ece7f05088ece262f383c678775da93a39bb7d7ee5ea28752c1b83c4a34bb76dedec7d1635c7968aee59ea82b1cce3c6e83afb87bbd06343fe1e8b0414128355357d0a602c8c5cbdf978;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd19a2974bcfcde2e0a6da8f724c75953fe9a235ec7930fdd36e5b2d20fe7c15b50f4508467eba26c03bf6087cdd6b0e1b6c636065d28c7f1ab81a890a0d6dc50a1c56a4010fdc618c5fea008cfa2a3b2ff7d611da5e92d941a92ec55be8cb146e5980269681bfc015072d7c573a4dfff1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d022ca8f8cfc00faea9697ae557815b1b40ea7937fe2e9c8db1a6da14f5515c671efb5ee2f3d35b2158fe74ff47a1d41ece9895f86425e8c85ddde39d285edc49551baf6d97425914b106d68ec2e6c0c741cc6fef1bea334a47fd44c9344c05b3af1e9a16826578d1f8f081f736d8a01;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6e330d24168ecfc7f7196546cd433c170ed4824c21857615792318f5ed13cd0c327c94b389c81cb63d57b18bfd11969d31e4aa37fb63962c7f0070379bf9ca01ab5e8e9b114daa3b8b1b11e141d43d93ee369838ee2b4e3d318d8b4f6103cda343e52620f4d4d9b9eaa5d57fce198168;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h783d454117609ab1db7c5b9e46a71a310449796144a3aaec9bf80bc7ff5a3502e6b78fa1c6bcd1e5213245ed223c63dc7e9c1e6dea647298983a44ed8d7fbd9a2d5cb484ab90658e99df1c64b5176a2dfaf4aea588cc14878d0055d4da8e462efc739591dd5c972ebf1abea4c74540bf3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h433e3260e0d559007268e0efda07bfc1a2285e4e2a20cf92abe9286876ce8f03a6dceb7dbcf9c80dda1050d7f8def27b3b984aa291cf6de697393690d6f7ac43f72e26d89eb1a835377d830b4acf63a1624cbb83fb72f1e38fa9352514fb2b9dede4e98d8eb00dc2ae725e7ffd89c33ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b93381853747c3caab203c0cd15b8de362239d75acf75469847723a5c2fd378d6b82872d860a70963b4efce91ad276c2f5c574333937c6c1a0976f47390cedc5ff8894721cfa43924d1c2034853a7257153b57bf4f3841beb44e0554f5d34a584099276a76e1074288e8aac8ee063cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48729c402a23a44fb63a2839127f435bf689dc3ee9afcb810778e6c9996a912e8cbd1fea56374d7286262ce37df6bbf0c72b090cb32a07a1e68eaef628c7632e16cebaeb4319a43bde2fada728fb58f2480b23d7f788544096d9bf3216d4e52cccceb8bda2cd20e80fa2a98219d567f21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h548c9ff951f8c0ff136b6c8fc7a5425d8dcfd750994c94a14b32c4492f34034675c99a476701698906f79c35e975b40a54f5d0df05f3ef3f942a3c3fcecd414355c6e2ed7bccb1dde82d9e1f75c0f6bdca05e28cd6c79a896e27f527c75a57114b95fb1f7757223973fed0d0c01aafd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22ecbf6426fb89566fbaff6cc6e006b607ac9dab61469e64fd3a6c12ceac6e55ba8ea315a7f959f67c944ace8e1b9d850c806509a83119454db7507f8ee6c64929297e65a29a51065dbc6280196b5a50088f6a653db6c2f1092b86fba89dde04a7f7618ca01fbe5f80b71d3688512f683;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5e9a9a5796f420a386344287210479582214353d237983da9455800a4117b37ebce8b4c724db5a755cab87cd043d5699576097e5387656322ad3e709714123707687d119cf0848135295790062e489d07f9dac5af8213746d736e143989a71e25b9714b35cee43ed76c52529f07dcf94;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc82334db6d1c0b3254bb12456d0913d2c1878c4158251fb58347855bb20e1a16451c569448f50913ce12a282161c96294c9e366fb1e822c0b3d826dcb3454b4f30a3f64a7b09363e057707e15c2fdeaa60adaa27f34e873f5b231a43ecc7315aea7408c00318ac12e175fa3e8b651f18;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e71571dc78e786af58261f088da387682dca1f267ab69fc962733eeab51223d3be847f1e2e5918f9cb6dfa584ed263f24e974edbe834347f48eeb3970e8033a38e25cf64f185e6e5319fd4a699e7ef21b5b7c00a720be7231a6518b904ed9d1bd7697c321b91e5da9bd9f284724cfd77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55523df181a2d6b45dc71f022c63d0d0c299d242533b1e999857878ef50bb28d9bd0143a73009e0f4ae3cfb4af7b2c835412174e5f4ea4473f77e16fa067cb25dac581672cc704a09e820c6e0ad7a55007b410a1e73bfb0d0ea645eaeab0db2d7fd1754676d7ef216abb010940c4702e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4b18b99ad3bee061882ca2a146d13c93897626334898125bee293713cb9d3eaa9f8efb15536d6cfab0b688de01790ee1f3ca16fa9cc00c5a250803b77d847e6587c1481407a1196795f69b3f5451f9c1eba5758e84100edf13396a13201bf3b03df06b79a14e1054ce084c753e27ac78;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h459659131307415799b7659e571f871bdebfbdf5f06761e75e857227fa309eb74daaf0081252e3dffde28e497c4c4299ba091d84b394927332076c54aae7d206aebf8c1a1ecc6843e87b814308b868c73b4b46e9946e293e9b906d43d381a3ee380aa15289f2893ed3e75d83075ba1891;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35d65832271976e4cb7af1b61d1967fa046a2e0a571f4779cb38cf8894274c2ce0a33aa6596da4327a104661081e6ca9e5ce9661fae0855004978e21870379b65b120d2eb1e4652c0b55a5abe14b547e58849d747e74b608be76c8bef3879f5d760d75cd1e1369b5d2b4a824f58470dd5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bce409a9a6668bf505d188998e1a532ca20e1bc30d9dc815474e4e5c2a92e61e6cf67b2037bfba54380cdef109a76f625be0fcd504d78de554795af84b1bf365e307ca066bf7185760f93a51d21c3c00004f973161bf47990af7991ad3f6c9704933a4f6cb6ceed270b187c7c465d646;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h260977629c8ccc32ab6a21fa351b7f4656ddee1b22f65d97a4b4ea852f8827eb55410db48f6abecda5b888ba7d5bbff86771eb13415fc9446ebb86baef2fe1ecb831c5caf3edcef8ec1ba99b161f4eac48152e4b44b8508e80d227f881e2507a1b538f2d4fac828e3d8834aa8eb803fa2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h246ee3c2c65d3b181ffda8a8ca7c13cbb7fe35c43564377dab3bb769e48f0ceb3c00da8e74fb5dbdd44f6770b50158bdff820b79f33deea22d94f76fb2601c06552c34be26545a212f6ac9ad5671c2613ca255fdad18d447a9770af173d24cdf21a62aecf26a3496a5b7f537f7dd40b4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4861fda8b9a7e9b7ce8bfc3dcd0e26857c2926356ef674917c63f4cb6706413e7f689c570b8ac9be75c23a7308895ac4b7c80d09a2f0cf22abd2f861b47c31f3836caa375fdb969ceb589a320e42bc1b88eaad4d9fa76bf99a2ef19075cb3812312b7bb98420b30f990ebf10838bb6c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50c704e6771cec8c8625fb0c0286a7d56b24e9987e31cd7bfaddfc3e5b90a1db7b07c96e8baedb2f5e3b5ab518de2849a3e8c3fe38a8538a4583ddae3cfcb2c6a347e150780e3ce622a5b406b23c6a43acece25524f4c841a93f2bdd2fe3c44f12e0b13e41c3fe9e9c96dffdde3156841;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ad79622f42f965e15876ae7873fcae4544a9e4f22453e00abd8f6bd214b775adc10fc4181c31379e3131f5f8edf8a348f1146f8ef02a88068fa3592e30828bcde94b8779febc04bc2602c88a30714086d9230d44b838f793f422c96b5da26fe2c901eedf44075c14074d99a777aaf492;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbdd6c939cd4fc88aa61d6f705141dd5014e392f71fa991d60a562f8aa9d1c3409322d372365af8c62094caea73f3ff6cd59dfa2d64d170dbfa1a99da768175465b20d4ac21a8dbfddd3abed59c145b92668713e4d8f37973c1d548b2a04d471b61f1e44bf912547968f9c8ab7eb8379f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc66dbb6636ef97b0500a517e91e1d97a8d884cb4b86151d64da2161989aaf799768e380d16f45961e0731662f527eb99ac4262fddcf1c2710354615f89729db646ec1a15073a878e27b2447cc25c23af31e702c6af62fdc0ef849f0ec3b7d4225ebdfdd698cfbb8ddfb6ad116774190e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecccf99fbd58c40f7af0bd46eb88030e3b59140e188ab78f153ba7978e14a3b05560d58b8b8199ed89f28dea9cd7e60ce05026ea0b8a051b8103de1fbec058cdc639f78628b5669c34b6e4316302e920fd8a1730347fc697f87ce995b8d37134a7c8d781394c94af195099c27f8531c2c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha75ee3c7e9d7031e52233aeb5bfb984b0edfe94b239bcaac5846dd749a140feb088935da6fef0649d6633859b8571dc3688ccbea57e6d9a6ac081a27cdfa820c2e07245023f447d0746755268daff5f1d27478900c285a580cf75572cde3aedee853f1cc16b105e389e28e25ae2ba556d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb655deee14ab16ac84998ceb3eeca2360ce73387eceb260f3487681af85580d165f2771d1b3bb650d9dda2c856ef154451e1ee8f86aa840203280dd946b3433d3f24fc424220b65ca409262d202b477dd833f7cdcc7281f9ffef602a7dcb3fdbc147fd48fbcd6dd446fa80bf3c7f7ebbd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8daf7a1049c94c79fa8a0fd321ae6b4b7db8e479e18fc028586f69ccb00fe45a2297817dacd731aa11ec145a5d62006812c8c95d7d5980c8067250c351f02a1ad6cfb6a4342b7573f940788e552f0d4673e3c16b873219d8f221921b3c61d55d73052014fd9c4f7f0965c2f533785f8f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d38aa94ad9c07601e9f395e1cf512d601542c5793747f736d9dc2b16af09997526631c38c2a1dc30a81af28ab336b7fe58e40498e3d25763dd12f87fec17ad666745d7c2e3f3c920b6c7be41a44c1bcabff944479db086b003529e47e4c7073c38322ad04c497aa2f0c4b0ca4da5156;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66b9c7234574c059dd9928f422b6d9de799e93a4b027f3e26b0f7805675b458c64122ac7b225c35bc6a4974d527585c24355b19e8d082d0e3732e4497cc1ab9e48e337acd1c6212255ab5edaf7aa26265400306389fe98819a5931d6b0a47f0f44cbd42565ec7482dab385ed88ceee983;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f3baed1ff28c47da4dfa2ad0571fa1e893cf7719b17c9d4c18e9b827b8a93c1217d818337aa5a03deceb289f82a27de92d3a750497131fd7e592bc53ba736bfe22780441a313b0fd0b49f672a4c3095b33d45b7d7fa0467620e88184a6b88e97055993c1850e0e110c0fb8a5d8e1d2d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h565091673a1185ac0c1374f996c8e0b8a85fff58317eb4744620047868dc70f2c9fed13a29c0e2b7d0f1ea085218c60d3a97ad20460f100959836be57ce217293fa4b625ad0e7dbec76215dcfd4741bafffb49dd4e589996a81c78393aae22973fc77075b41ae381e01f9b0eb2ec7fa90;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb4038f6739441da7e485c831ef574c2afb4e4ef0496e00875b14f869f10d6d448753d920542da40cb1d68f0a316c7ad4b8484e60e7776d88c710e452f4e46ee55670b342ef96fe9078d4485e0964b0c33414f7944b2dc53633c7356411efd66067c957d4aeeb6d956c57871c2a54de25;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h488542c6b3a9913e5b3c08ba9871a4ab63463c103fae3679794c8f66ce11bcff80013a5dbd1b4cf0de56fa74c02a7ced9f517750e3676216797d51ec7cd7976fc973c693410288752699ba44fc22c4bbe3ab6237361cf886ea514e891e173647e49acdf26e306c16cdb5592f752501d1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3426bd6be02fd838d5e62c08c344263b73fa789d977dffbd5fcea95067f70028fb84c3851ebc0d2fba0ef8b4dc23dacda9c17cc8ee3502a781f43c5689c13fa1167bd361f6dbe0d2c96adf4e898d600a805b2bbe4405ba47a37ec6bd09a6dc9c8b59472a0ee538bbea2ffee52a597687;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36df3798907a1a733bf872e76c9bba34436ecd4af91916ede930340a548b9e289e5f52c4f24123664342e4380e5ff60435516a28f08ea57aa3a4000e4d23a2295914c0e584ab024fc2c2efedb15237291b900392430d6c7fffbc62ce8597997f94ccdfce627dd20c5021bd9a71a8abc90;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d0281bba4dd68022032c930b4d7aac491baa07069e980d733730ef9eebbe8346fe7486da784ca15d43117cd1c131650b9cd7221b68bf0883dc6ecc24507c8770daf8d48dd0745a911944d4101552bfc5ba1d0378ba79211d9897bd9b6a619082e1ba2e7a474ab79aca1d2a4ea0e4c42b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bb4c1111a32cc66b1ca1d1fb93c5e4e518ea18bb80a7134a6707e54b8429ee0d0de80751273d5d25c0485c7a5b4505175495ff7d4d15fb235c21b8b44ccd734823d1f3799777089741c59746b25c444def1efa9db71b08a41e0943d206165debb220a14b24490ae46c8e0d23293fd953;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37b379256a7bbc96485f724c1c17b07acf104cc970a25969dc96068cb4709484ab224d1b72051ba2919815f8e6739530874df76507deaeb806673790be5cbd555a93c7af4b8b8a7d3b74c71b6f6cda7af0f380b1cf38eb89f461b31a25b68f28539b080c4a9ef39c8f466be3d71526335;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb858739d48a6c2e2812450eeeeec32f669cb85fb07acb29ed60f02f21f9b702721ec4df0b8e99c62f821d95dda08bfc6fc446476fa948cd2f48793bc90f3e66b9515f0d5cd49644540e8947b6dd418843813b6462ac8d629987ef6f2caa8e5e689dc74b9bde81ff86b0151f2922945197;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6d49b0d6478bb58620b3abcfc0853ed5beb1e4a884f96930d2ed1d364d574715fd1b89cc72e946bad4b104be3097619d118629c5386cafbabc9f247a9df424358fb38af08f88951a340df92e8b6989dfe192fa297ffccc2533520cecb2e768e483eb98f1211fcd1ba45d097302ed72f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c97744d7c9c08e44f98782f26be1eacd87f977e6b1d5330d2b1b09061ed1c1c5fd03ef69a7653fe4a7ab93a897b0a357aa2d587303edb16fadaf47d74857823fbd5d79b65ca88d5ffb748e47cf82ab56b966c90396062f0abc203edc30d1468e71d57312f3c3acc699c93fbadfc1c9e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb523bc0bd0fe72e75be13d6fdaa2ad21112fcf40ee7282fca9122588a34d8ac7e8c80a620393648b1d8eb62018156019bff117d6eb2b1bde2e5926e29eb3de90aa3d78369483e12bf436dd301fe1e7d336fdf5de23df91d803a0f695376fb03923ea94e7f2c89f95151c6f51b85443a06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd408b8e4dd11a50326ce51635ec0ace5b00fdc08793741b521766ab9bfa2d9d2f7373f369f408ac49841524df8a655e1b5fce5ed2cdfee3cd63074d23f31fab8b07d025f130e3b0151198eb7cc0c9890fca8bc3c7bf584d30557f114064ad0d781a74b42a964c520d827ee9e42d83ee6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80abfe02c9d08a670c2d9625301255cfac467bc92719259704afa1ecf195f75b067bebe6a78bf5147ac01eeadb4a52dde7d39434d87d007ae36b464d9c5f03456f8d71271e31fb57de785bedecf90e9ccfa3e018e676f9fc0d2d00750d2ca9f3d2e245ac64bd9c5608127ad738b82d834;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha70447cf6362b053faba57f546cae28a68619cf8f81912b23214b18273004062c9aad0f144dea88af036ab1317da7967e85dfdc0bbb25b8b825e4d45076314c16f1c277412e11b396e30a894233d5b737904f38e68591cccf3743e182e69e2751f0d56a75dd01d13bc8ee20e86a6363e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b23bdc0137c748b21e7c6145688e25f98257c746025e66295857468630ddfc0fbcf9c0ca8d9584f2daad4230f22210c0c8e2a078b7e35fec44caba4792ecb00a870873ef3a7e090cb663d5bdf8866479435dbb0722ade35e18cf55af02e65ffd266002d181767ea59a338bd964af236;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h669df634200dc52d2f3237f90c695da04b1537252701c5707b5e939df07082ba0e7552c040d3e46f0cc3ba3a390eb4d486af5091464907ef450917b8abd9aca557c389fe3e15efbb8232c4024d71f404e21104e072c4ff9f8d0f5aaf9f93bd4e2625414b45affa1927eccbd4be359540;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0d9a90304b4ec4df2ff644f7a1ed920d0309970cc99889edc9fead3bfc87aac57eb1e340673955c883ca6bec00689a065fec2d71bdb2fa60a7336a6570d2a0eaa439ee549517bc4d00e5a6760bfd4201cd56bfa25d40652f4d126f6dd8a4a246068449705944db9c70077b847414d0cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h188579cce0ef61b00ddbc06f6696ae4ac684d392ae1373dce0c74ca79d4f4c0d498844ad5acd366879241201d4539a19c21aea72b69c188f27753ab1c9440ef2362b9add2c3ce21269cf85e4d2b177b5392cda04a3c2e2193dedb4e7910dc4d9d7a90ab416ec0940f21dfebf6317efe53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h211fdbc53cdc25cef740d9beb56721d644c2037a03126df009662c1b0dfd46f0e39716839f81372fa194605cb3519a9ee2a5ec20cb2ba34417c525d47aabee36d453939e6491258a4aada85b5e44af949239e52e169cbb3d40b43c2449da77b9d41cf207cb5544c7dfd3830be25fcfdd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9666f47ef2e2fced186660df6b4284e686c14e213a22304e73316a427581ad2e3107752a057b2e7c94efe2f71c896945e290b61c53b7500980b4ca8422814832a73c1d084e1c7f051679ea0ad6676203d7ca2a2b87ce8937eacddd9b2199133c11e00e040a05e85f49642253fcb0a0d79;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a182f65850282afc0b9dce30defb1d31d50aa6418a6245507c9481d24a3d97e96f5ef78005b3a4439656d5bcb0cbf5e6a478218bdce6f6ef3b7c9ed5e53fb0364b768d316226a5087245e8106cfec71448107185d402495306f92a231f7122cdf7748ca1e6627ff35924427e022cdcfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ac454769a8be92934c279868da3bc5739f7c0c8010806bc7bc5f6c4ceb1dc2051f289add3571ddcd19fb1e1720ddee51d16dd4b27ecb488238d7004fe5c3c6e0c34392835761f558d627c17aaf469725d431a891a42a59424b2ae8b27d08a6c9fb80380f53270395a04a5b794a07c213;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88be28cf6eb0091238263d41a5ba8c1ce6b929ff9aa842b11941d3a34028b08c51dfac4330d8c95b45aa16b58a85b2cfb3fbcb177f2b09ce133dee8be5f32d7f8febbc5869ee4aba0758b4ba1126a794fc5874c2d3ff176f23adeeac1ef388ed26b043bcba44841fe64c4343e4f8542da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6379580d507d752dcb2543e04cca6adc689ea68b39d1cc0cd617634d448220a3d4568ee06ae4f6f01e3d510204f6f174bbfa317106d48c5d52827a54c26f513600f7218a81b723c752bff3c7e8693a6e444f5f9f8d23a129da5fdd1e33f0e18b7d9e4630626f64febdbda617d2a297ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25fa0c6c4e0481b45dfdc2bd04829194f5370d9dbfde44307f43dbff60e9ee3df258b2cd81ff2ee82c840d4fdf51630e2913d34ea4afecdb4cbc53de8bc7c5136ff37a3f5cd63e0eb520e152794f214ffb34519190106b437989d653db918075bcec341a928ba0bb618fdfbb574a1134d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91b173afe40a3c32ae4dd3c6897716676ead3248a6cd4cfb8c31af3d1a1b5f1f607e343c4c0d5000b284033e259efdf62159e0da8c4dc7e35e82263211f44b18c28870dd22b4ee8c7ad5d1ca879e407ec5a4114a516b2c236fa19456239ee53c231f59bb1f71916c5f5ae7dc5b6341b12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36408ca2eb18d89ec6e6120a1e21f0d83cf0f7c47a61d597293e4a8597cb47cec44700bd116a21ea5a32641aaf8b0cf1c18fd743f41434f6873d6214003e06250ff3e0872d2eff39dbf6a48454bb24b364e841a12c5c50d2e13cfb06529180fa4ec76f5d6aff195e769f686566b9172f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb3b637386ad5f72d11ee5d2a9d5075f450546c23191dbdc4a8f9ae61142dfd2316db9ad0860fec94f12f4bfec68b5345fbd1ec57d330add3a750020ee8ac2d02d0b435d6a9ef664f81234aa852af5e475c3a1ce77160e042e76b25b4156839a5f25711456dae09653146852c51ebdbd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1001929f0bfa732a99310bf1ae71fbc16baf9fbf0feb64f18a787307efe8374a53dc1297e639106712873a0cb84d0adfc78c122964277b37394447562c257475d514428e4590ab4b5b7d2c117bc39d0b9e7044585181b551bb9d397fb73cfc21ba2bcad9fcc8d58e78de9e889746e200d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd46b41bad2a3099734719b2d7833add98412d63df1c3f5efd5da19294cf72938410030d5611a97006a6b6c50581b1840b73536134d3d24cd94e0c677ed400873bf5d609ea9b0368b551bc55535ebb7527b534dd06e3c62c6bd04ea7d6fa2f421c09b8c4c3a50b5b79d8b8f8db5d89c2f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd60432efa74c9350540f21c094dae7aa1726700355e103dfd6ed73c5a7ebaa80f3f0b0bc0369332a8cd537d259960a2c4abac70405a2a100a1b03e590f6086db680dc211d2b61d42492c7a481a0aeecc7b88141a8643d34ba014154aaee0dd1be976c866757d2339cd4984e127f3ab409;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eddb6e005a09e6181ea37e6adc218f5b44ab1a325056a892f3b567eadad436eafc6853617c7d4aebe7e3afe6758116b72dfebc5ad2f814f06dbaebe1afb092e815aa54f0876d64368512f0c0a4ec8fd916d1a93b8b1b7b3eb8e61cbe3f637be968ba76e9449295353835584253aaafac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he72f78a9cff9ab2ae3dff4c0cffb4328af181da951f0a979973f44e200a7a31857b9603f420ee2e0f41e5741cfd686fa4f386d75994195f2b2b86a74ca58e780a69f464cf15b4e9ef895dd5b91a4a023aaffa04afa04e94076bcd0f150ef30890cb85699abe1ba7552ed0af16579d439e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h317b47eb5e2e4324194fa4beff6420a52788d19e07e9b5dfad06813b5e2bb5e7747122ee76648d3526774396d9b17e7650f25eac212d033ae97e780ef37450868d7cf7a885e64bde942561686103a0ebdedd2bcc4943e2db531bf292d44dae2602d7901fac113145026aee080abe7a53a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd13e252e64ddfb9e46ce70fc9fb0cc7782e5f803fffd5f7eb6193021ad9cd080ae03b6550f43047da7ab33f67e8cbd0b091776f0ec92be0431c515d1326cdc809f543cb9dfdde3a6d30c88ef357a914aecf45a2744592ad141d9f3a2e13fff11606bf8b382a006ad07378d4950add2174;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h898c19714334a5643f3acc19186599f9252db26c3ef42c0f77f295461bf2e16a04c2f44c9b8c0c2ba09fa104e9d160e5372ab3535ffdeb8113308d5fe8e0a09cb72be6e23daacfc556e2c2c02cad317105eb6266e46cf12495fd18fa1c2bc379aaac0aafc31fd91a6588230c1f76dfd67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81c0b97baee43bf6c7bbc8f7b14392d8e9662d867cf6901089fd98154c2f08c69ac65d82951cc712c0c70fba600bed2c16612a3c3846500b5de28132d8f0a2a8ca4e60fa7f5e6d82329edf0c4ee63a395b84900449ea286d31a1cf287175fb96a8db52fd9a287b230df08abb87c554a8f;
        #1
        $finish();
    end
endmodule
