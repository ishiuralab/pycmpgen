module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [23:0] src25;
    reg [22:0] src26;
    reg [21:0] src27;
    reg [20:0] src28;
    reg [19:0] src29;
    reg [18:0] src30;
    reg [17:0] src31;
    reg [16:0] src32;
    reg [15:0] src33;
    reg [14:0] src34;
    reg [13:0] src35;
    reg [12:0] src36;
    reg [11:0] src37;
    reg [10:0] src38;
    reg [9:0] src39;
    reg [8:0] src40;
    reg [7:0] src41;
    reg [6:0] src42;
    reg [5:0] src43;
    reg [4:0] src44;
    reg [3:0] src45;
    reg [2:0] src46;
    reg [1:0] src47;
    reg [0:0] src48;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [49:0] srcsum;
    wire [49:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3])<<45) + ((src46[0] + src46[1] + src46[2])<<46) + ((src47[0] + src47[1])<<47) + ((src48[0])<<48);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb29cb2bec023d5a17a19c6d4e684c628e67d03f3437ac6af2bfb0d09af7f098278d5c8bd6f8b1775debe09932aad7779b3687fa5f751bfeb287d416533ef7c2ca9ca98b83f529a30a2958de1f623;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e22d2fe29909b0a7487da1a70cef4fc4007c30c6808a65657d5d1d2d4881e90dc4ec2cc69f5f2bbd2fd7fafe9f72f8192173835f5c5e626e6cd1c35f18ec429d799943695081e6b0fcf5ebfe39a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce322cdb782dc145421db72e40bcc72e264c291cf2091f11eb199f68e1db25038861e7a506d59e2c95b27a0a9d2eb69e40bcf7afcb0d1d6a77020d2028da74d0119727d50390dd39561d268d63b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48f5e1c5ce7d3a606655a599d54c1da6d2fbec7f8da9b62556a693bd23e1f275d9ac802e2124063930271922d063e7c7613ec5c682e3fe3482aad2468271a614a4113f68a64c2a9eadbeff9b3208;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h365559a350a60439432223a8f0078cf824643edfcfe98b79773efc35e7e0c8db31c4a309e19d42a94be60924a5923a0dc3efee0d3fce78ec91e9d32eef83d0b0ce21534bb8f133685fd6174ff5a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1fa3392426859eb6f118056cce120e70dbec2db5190da6831b7abefced7f0bc3e90609987e43c846cb5a218f4e7f91602ebc6a745e7b36a32418f3fd6fc8f6c07a083bc7e19ac74c1c28764a883;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb39a4ed6b84cbcb4310ead3d6ca15de2158ec2cda954d10420b09ed979348df77b52a2dfe93112eb1d5f64d92fa9e40b72eb3fc547b2f6e73389c2d1f85306455a2267271656e4a9b2cdcaf83105;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12559eb99a26a7be39308c63e98cf2e2df440cd35ebd06fed2c4c7012ec04af18aea4e77a8b5366c95080dd1ff74512f0d0cffc93d6795860b07e83db3f3dcf11ef826ddf2022020a9d76d8703a17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1159c104df079fd906bdfd259950d9e3842f457ca5b1e29b2058a61338f4d926aca3c7ccd302f4d77289985060efdba793cd9ad4c3911919e725ac07a92e9565e83a9379135efbb9df8e00d25daf0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff3fa4568fdd83d8b42e649946a3c53c7116ebe84233bcf988905d95fcf517f346625930de3a7d7c0fd10f89a6fe57f8acd88da6fa1b2c6516effe59c13a68972ec8c787b49b40640b3e520b4855;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d4e7e197773e25ca449de4663f0586f73b84fc454bc63193c53f89665a60738968cf88ddfad4ac72469466b88c5aca4cd7538842c979839d3bd8b4f1dab2cb41443fe4736b3a4f5dd9ac2be9161;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eed0ca892804f21657584dbfcc980d6a95a6cc2482f3b9f1e687eb49979f18647e9be3762b5fd09d706b82aa7b34617103fa6f53fac83c7d6e52288192a4d7c408a9aea9c4b6c12770d7deb24aea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189a379589898fa0ac8931c565cc2c6233c61462f7857345c87485b67fa80bced817f4fc8d18a5755dfbb83e77f0ea488bca541ceee25278ba0015d70fe85b6fe02965aff7e0d2eccef1142dcac76;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd716838fa531d4798f160c8227cfb167d1220a2a480d7168d6b21dfee9a17a442ff04ade2cd6c6ea22da7c43b795290579fbba1a7dca5cfdac8d6cc024b98c1b77b587fba270aaa5e19659b60c92;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1478dda16a4e85d47f8b0348a1845b75f878d96bc17c14fd90b400c7c9e6fe153fdddf9189c39a9e993320a1cac7282436e60b91b459ac12cf4b58a69da67562b43f8f01528179e15df7d3c793cba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e77963303c48305811d69e3a72b2daa71f8df5b6e56e94734b2d05953e25e0bc5248624c479442e8acf5514133588e13ae7b173dc568e3b1e5f66ba6a39e229869e768c88eb718570d6a1d59de1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5da2226acf050f2f6d61b5b63f6fb9f14ea7704bba1cb4fedbf41f88ed96fabf693b8d5eb9710391508dc21020c8e8c902054a14edfb08be03cc1680ec01ce02c7fc099b783ba614d5c9d0ce9198;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36a72465b91971a39e54364c7bc02c81bb9c0e17be3ec39acfbaa9517326fbf5de6e27675cd0b5e6e188915eda3e83cc49d0901b8ea03390a1b27c3854d0125d9b385498d5f67442bcd94c8dd065;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47033e3bc0555db68c93f5a5c2b00507c7258aecb2aa55ec157cc984816c64361df68e9986d0d7dd216e601edb47a61233c1a735639cb45744565c1b7d85b219e4845f67f793091ef639c4bd550d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154aad23326337929f60aac16d8c19a31ba563d2ac292df3c66544413f27412eca42727e532b1144e35638ed7d0ea64630a8f49b34eddc68a6ba9cb274b3b48455557e452c8e8b0144773960518e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdeed6d09d7e9f3efe78242a919cf3ad429bf7053f2fb5d050315e01c2489bc5b5e7e535d1a03a6a1a3cf143cf1d4cd27985c47dfdc3b0f5231fa486b1b7e568b8fddf52584d7fa367d4cf15a04f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38c0766c4fc6f34bfcb8aa0832fdcb49ce24afff2080ef534d148f9af9a2a82c4bfb15410fe4139d5780bef35503534e35f51bc91813470a40b62401bd4e134a0b136e83ea1d0764a68c4ea282de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c53ff82e4882a9598782cb5614959a4ac77fd8b29adf63318cc957b6c496d9f9e642c29a0c16222028f290bb5f1735c59406c4334b10371631f9a779999f2fdb2679cd1b470834f738a01d3765;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89ca8f653deba6687b4b3ab99685075e3e63108acc8517da36af6f443d9907e29cbaea1556e36defdcddc093d9e4376f08e5a950eb484b603545e76c573a63164306ab41f8e68ff47886eafea21a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d212ddc4e193893ce83350e8dcf7b7dfac078cacf9341ff0320cb0ddc51a68952b9863196e9ac6d1a08f4c23b9985156c477feac58bd70ff9a8bd6a4e40f995b089350753f13eef8d5fadc33bb3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c13fab9aa6930967e3035e9e04ef2b0b9b5a9b1de313ddda132713dc2e3e94256bf0072ca75ee6a84b70d15191e7d65c53946652ca7cf97e5d2cc2dd02c0e73df9365d65e17dace46c142708030;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c96326984316806f4134dfc75ef057ce07d98cbff07b6a1ee2a8a54c462b13b14c8df781b39626c5424cea1509bc73dd8b9615301e71ea0c7ead1f60131e96bae86c88755819035abe7d2634e4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1523667b94eef594d1fac31fb27944fabd07dae024bb18dbccb351da19124f81d04a8e5205278461166ea2ab384b232ff90cde5e915a7cd2ebc3b4c9bb2f0aed118a1cedd9bf9589d2d1d6d984193;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0a7553f9974de3fa990515c58b7a2d41a1f3a1c0d73f25dfe877c6642ac18b18022f3a69c5eae27b541c2048251f4978134552ac2dd0239ecfa69374fd979729788b113f5cbf3a90630e8fff6f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14536b76545327455aa563357d5b7b56b2fa92e1fe601992c980294b8a21d9ba84ecc58c51dd2357da175304a9e82d7285e82f4ded3ca17d14eda6ffe852e8f54849bbc2b5dcc96cf0ce0bd96e746;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1853e0da35f87a7024511f5eb8e4e7a8be5da88c150c3a83e52a52bb6a1d48afad32c410605b3936b36021fb0d621fbd5476e7b50cbd9c6e19179ed4de645393d88bef48fb96fb174547758240579;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac358693704d9a2ed0cdbba4dc9d237391115e99661b4bf73aa284970242fca42820f0e4d16bde43ac7f053977a462bf80d87028974b8aaaeeec071ea569291f7d4068ae6540d701f6df6e4af79d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175eaa0a3e2a72f247e12df5ea9eb67b3a9771898c8cf64a26be0c00b624bc4036219d69241f28defb985fca7cdf2c7bdccd9ebd14756a3de0b3f0e470753fd76e571d3ede71f8df31fec5184935;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b57fde887b5a42289db7438f502936ebe7d82554f2f5f756ca2fcdfa9f713dbf7e75194053473408b6b39efe81af9003e4c34a44563e3ce29ae0a9fb016a30931889c683f8d3b6500f04b86b30d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17eb5cee6a1726ed602bafc9fff00a6ff169796433b965426365036ed97e48c7031a2671fa7cb61d31de3a1400cc6bae326e2cbcdc8ee109b8de388f5015084cb7e2b821dbd3960e242fcbec8b07b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f15a2f25f65cc5208ce4397e9a4cc00577fd4e88dfed677485cffe6329af581ce5c89acd25a35f9002ec9440d125829e037504fd68a7fc190edd5d18a68268cc27933af1ab72d4eb5c2308158d25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h554eb23c230ccfde1d848ddf59b87f23dd8ee5de7715afbd6526a62dd68d7162e08b152ee8b31ff849f063c76282d07987ca370ca49a52f576b7d0d1b32961fac0cdfc4c16282ae8ae31fe7bb9a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109d0b0852c547ac9cc28e5610fd7d082cb7f9997b141e984081d79632513a20bdf3479987977a70d80da1a022c169d9f303724621a7b0bc5c756243bd7e01794cdf68f114ab840ba9cae7c8829f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa5807bd395497a6a665edc8b0bbfbd18b789461c07e5350cdd0a0fbb0dce11ea9192876351a2d52f649e582f754a290198281a5350933f0050ef240a77fd9cb7068c1d6d6b2cd899c14c6660dd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf48c76f96d7ccc0200c6cdb5e14c7b185f6eb4ecf821ac0077e27e115ca894d3e3c77899f53438143f568a29bab967ada0fc941fa32e4367ce8d1712e298076d0329a9026c40b5ca75bd82829f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5306eff8b9daea8f733aea272c2f93742e50e715631b0a2bc7b0d6a27c40e7dfbfa695a04e5e068848f92fd50732fe5bec26909c47dc088f5f08156f69be00debff2ddbce8d40e94b8b39ee9ac7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1430e33e8e576d3ce3bcc412730058fb7236278c8f8669862e6fca40a1110d0fd6450d2be1056afe73b192cbec1980e2014adb904f50cf75bd64bc64e868aead6e4c4597d75e35ca15efbde0a45e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd54b584d4052614b0303ecde442d207aec281362778e6bb036b4a9f10ae233fd93a47a03a3596a68a3f459cab6f91e6e36a539d38543572e1b95ef5e9b761add33681a679dc9c4e58e704e197a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f84fc3944ea1c10c49707e15fe8d6024aec1645640918014cdc61f0ea8d6bc01ed74d439479877e06281079a2e4d5eafd7d4fd1d896069852fc9b0de25b1f11421f533596a2d2c89a60f3b1e550;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd153858af223c745dccbad56d60ca2c83d257f9028cd43856818f391fa8e74ccd3ef7b424700312afd6fdda104bd40739330212cd5fa295128025bca217e9fe0e250c716c58ea1c628b7f729d9be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1847784040032e63041f85e362bd11aac686cbe5a6c2e5bcdcc89f103303a7b8ab8933d2017bb9d5ae0c00ddaa6ff0b8308b61153f0dbda99475fc3b15800511e1387a10fa10aaf049cbfdb7637c0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e4c6730dd6ee70a9f9935c2ccb8f14a5cf07797e8a84ee6e3cedf055a7658917ae18a0b87840a5816323d25304424a3fac2af0d67e2dfffa573345709ba4c2b186d21c6c89839d286e382e1d78a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149d55964f5e1b88d566072a74bc8c9d3591f476690f4bfc4dc501038b46d6a8201d6c96a410700b6da92000b060a50f0f91f05eed81f2f884793c8bc70c3760b83dba6c93f45ea3d1a8f42b8b657;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbb188a8d6ae737ea44725054cdb0583ccd0fc859d8f26c0c82e8f3f561212b794859138cd7fed8599e2cd7df941a8ec55495bfcb9d9dd7f68b35eb280746648fc4c89da960270f22f04693f90a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e09e2500d65535be420b72218daac71057152c9b13e073647bc2eabd510f36670e27037a3c90f664512fe641d6b5f0286971d64568f035314a5f6fdfbe24150ea1726df067f4c3aec33b57a7a185;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f558b2459ca46f611cc94cb0d263702b4b4f739356e0e4d9fdd04a9e8e8de9fff8158e4e557aa343777d0fb74b348863e6589fc5750aa64b0b35cf9d8071baa29bad106fdbb9b4a7828ff2150e17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ec11601efd3a645aa459981e5eb898ff0e17a747b157447bda27dbefb3a1657a5bd78e0d9246f57ab0afc3384f5c6e2a28b02d3388511dcd3d0c9b3b123dc4a90906e437eabdf27679bc70a8019;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc9d7225aec15c00bcee2a416f537993a3f0c5c9a02646c5908834a58626f0c6389fbc881fcd0a143edde478ca3bcbd9a0f7e7933ee8a1056ba9802e60d318512f009ffd722fe9d051b9983b3567;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16755348193815d98748f1414ec858694c33e22e6d5ca3bcbb52a743ae55e6a64e9c61089a0ada30585cd801f4d411d7be34b277437e1567f1b4b931b1ccd3ead07faf3e30418a0696fcd770dc166;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99a47db62d5e65db06b6ac04c030a41533d8d354e8dfbda7d64eaecb5505b1ae047f62a184adf41afe2b93901a41bdd353d40a02e8162cfdb3ba4222d75e1add44cccfca7e0a1ff5274e5512d687;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18159aa28edcf4040fdd7cd00e59ef32a7dba052ed786fc880033973e9a67dfb0c46f5cdc9f90e772b5cea9d148e00c05be6eef2dda221900a6988300d7b1832b56355adddc49219dadab792424b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b31f849ed0dcaf8a279f40bde28828ffcbe6153d30ad547c7888db4e0dcdc80fb2b5e91fca9a34c5d7db366fbf0e029d2b11ebbe1b8b6a699c824f4a7c1ee4bcdee8d16f355215ef12f8976bc07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1486fc6afda220711c3ed3eb5334192c9ee480414abc27ff42f99fdf709aa7ab358035d27624fc471a40038005be9543fe6ef6f438d08bb0cfd97e8bf7fa44c6716b8a68a619ec68f84f13c8258;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ac55b565be88f33471428d263dafb78cada1b2dc87530a895c8161cd89219a1b57f7926531d61f3b71a42a9b3fb62c6be809cbecfb505c8a31af1f9c99884566157b82a2065421e66193e77884c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19748f18996f7222c1e2d004c5166cca001e3d796c3e45a95f965a2b0be261fe74331ba1e355d670ab000da0a7e8954b6731d97f6c940105f5e63c636696a784bb960039335671fc7d2f7f997118e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda85c2bea138e354fb8ef4826aa4415b65ae3b50dcfc8fc6d3ff3e32db9f15de0f42abf3af0e02257b6d8fc705d919c3eb661267aed7de4fe8bd2b97136104a2989f2822edb695ac725133dd74ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d46fc388d588ee61921ec718d44f528f85a6025e38eb49a4a11b456510b98d72d49f7da225281d59a5c278778b0514ead56252d71357f7d1ed2448a4328bdb529d7e27200a5bc61f1953f634cf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9fb06e4f8e260982da715c18f2eaf24a0a7de48e391e367b4b1118bf0bea642d6b70faae1813465fa18d171883affd12052da89a2dd06bfa9b810ef503c6fbf2652c7a813d97411e77db7b2c3f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153a33d4c7c73affa30b9958c534ae152f8eec88d1daff2b1d8e70a00c2883fa397aa2735ad72ea51eb2e1f5f8b15fd0fbe77f12c7db151e1af71d54b3f61a35815ae976032976d12cc68a0c77790;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127f89fc84dde6bd4709cab5cb93fcee07c19ecba84ac500ea9a5b2db242e00125d4c90d52fd29541afd656b65924d2c707d07a7040a34a7a3d625713def91314fb882181ac498b211bfe1acc08fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4a4ebfc026856c33f2b58a8b49f550aef186733498c66665eb2d67c4dfa86f760a26d4b85fa22e1cbb78e97d19bc6074a9f457795896fbafbaed01d1154bd4124ee493b8cae0fbec1f45c3972e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13294bd75ca4bc11f17dc9fbb39b8a8459ca3c0ae8371b0c746b92ca01392480a2a0d77b28d5c48b9c9b6fc848cc47bfcc3c59069e325d01fdd609832a0aa321412cc86e94f5bb926f30b4b1d827f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha221548c72da60bf942c8991fdce0cbf63678b511f21b302876cf79fa8d0675318b54c3e33a85946bca3d6ab6a366bc65bace2b55ad8f24682d6837adf42e92df50a8f98343e5162c78cf7350d88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb075f1cf3b1a4f3657af3cc74a24ded2fd06ae63cbe2d0015c686e4d998ed0fd9629756c6c5ee7c7a5aac83392fd41d78914f15d8261ea1e91567f67d0d3974816af4ae1002ffbbe1b57c4e1d01e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1513902ffa7b14cb59260d8e7ca21db0bd3c9d2ec2a1bf91d0de9c569b71d49667588a7574b49bf1086e43125c1de7b20820200e26d820b5dc24c3bb4e743216013b818a0b2d332919f359606e02a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126ed43a1ea3d0f15d58eb5b742be35b65b147c9d4feecc5ab675d1210b6d48002781489df0d91b735aba8f8bed442a1dae4f19a49f82cb49701b6208ee718f85f9b577685016ff6d98e26fe191a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a8085146cc732b85b2e8d5d846aafb8256a6ea3cafdc3642461d6219e20947191d0b00ce5000e547f6a2439b36f4e423fed7bfc56ffd09c2add842960553a4f86f9141e6311469fd670717126d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b7e4e0a3d25f16b5cff40c78ffe33ea7e14dae124d1e67e70e16b97556a638a0916a006ecbbbf5d275c623d1fb47fb343cafe6f0ed99ae6b5ae4d648efa736480200549919494627739c1a1a6db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fc858dcdb537f3be8e0e5e011840fbde52e6d2fc4547e4cc1633381bc918ba7482222486ba515601dbb7c8370fb3eefeb796f4d7ca6e75d78c255540df80c867425789f5022b3afea09126a8650;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7a816feabec798991fb1574575e9327e44a07a670a2a5419cb58ef18c070df12c55bc19872bff8984de5c9a747e8a1e8fa3c23280640c7f26c209fc226fff789abfa28fc4692050bc6de20eb52e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175d0067cc8056d86b322dc1eaa568c04e55c2512fc8c3871c545c8477cb9044b981d8dbf47d79f31c3fadbca391ed8b370f45971b194250130deda43b97476ef1a4fcd18bdd7057893f1115f6557;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fbafff7192cb76faf5cf19c4488d8a9d3829b55c03d72910ef871cc1f6c42e50ae06bd6bd89dd5b50a888900b0a50d0dc442afc4acde79998ce04431161c876ace52bb78f3c205f8820c3bf5064;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c191f85cfd424817a3619ee72c02c4793f65c16c5fa1b222a3bc20f3acc10cc797ed8a8a9142d55a359fa65c0cfe8b75b1f3142c15adfdc06272a9d7155459e8124b797fbbd2317c81a3e60b431;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd09a8147583f886836ce27cc2b5dd9377d24632f64b9116006860bec1f826939e0da5bd65770145f58a89a62dcbf66337d9765062f5e83d8d0cfc03eab88131ef20efa0774a31a40e52f628b9fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc51e59bb56d7b796ba892d5d8738bbd638a84a1a144f603374d7791b0a11598ac53fa3836c71a36f13879d452c9f7d201a3b407a130764f861f9908b126bfcb2063d09457584311d1672ddaebff5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1243e6c33b53b08a073d149f921f7807bbf2efc78bbf6d9ebfcd38992f4dca314d685870551679cb1d1906bf1cec87658f02c7b9848ee3820aaa461cd82c9c7c1c6a967efb6e8733c65e43f522b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ec0e69d33f3066b2187d25cf8cb163d1191bf3be5cbf56c4fae200465a3851adeee6f3883529a0c9de1ac9354dc4b9a8092013c86392d5c1bde0489c6c56a2f96a4e4acf7efac5e29d7bacdf93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1368182e3e90f0a0b8c9dfabd4152028f3758bffae9a1ffd38cb688a92dc3b61718ba2796739186479567e1067ee818254c542dd2c239986ed6a17e7bb1cdc9075c85de3821c0c3339045e5e279fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44e8273d2f149a432d0a9c4c6fd944b907eb6a5213bf45a02bb17911971d862cd79f2ab24b660bc499a0ff6e482ea0f978b439635feeb3e5e333e38fb1a60965d1d3dfa0dc8fd3455c4debc65012;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2130634805ed46f0ca6532460e27f91fd0e7e5f63a4a1db0898a50f28a183c6f44f3f666743ac49b1741d0748a4fd2be85fe79cd4aa9190a9cc91d6f58fc9c323e4089641d8a6b3e2a9303297c09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38463e135c9b116302774d4e0d6971b8a5a60fbb6191ada86fccdbe690ecca00c1124f988a48e4614a099569b60fc9caeb379fb84f5ad8791bc653ce9b9b56035083234444aba1f7b288ba33875c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h688f5010327bbd116de62b547bac47caaf6be13e968bc388a6ee8399a896e7b39900be1ba3e1f8ba4bcd716e041c4993ed01aa41e40e8a5f88cbb7a4d9c5648387851e2315678dee6fe9b1960f51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e577db513c59072083c93a139a79e7106cd16d521560e8c3fc25ccd5825ae42a2e87fdebaed99ba535d88cbe9a8bf2e0f795d1d073856f2c7a6ccbff2cc03793b8fc104d82a94ba12ca99f11dccc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee68d6699e544f8251a6c635b12843dac549f59aaae60d74750e91097d6c86d7acbf4067bd7987daa009956bb82f56b384c8d83e5d86504f2d06be25cadb149e28431f8a2ba429a114f6ed473c68;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101b721938504163cc1132a817b52f2f937ed30dac0b167121882e24e3e31aff13307c74d7daedf0d98d43efba05e62a948747fc53fa9e8e9c0f1f814f6c82f521c78a40eb463de4c4eb34d6078df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2b8a77a36154beb186af6355b3051eef35605eb2ac9d32a71097bd62643fcaafcdbb32e6c590967253ce0a4f3a0a4b83f19f2d0ed948b4cc3aee0bb208e5fd25e81549738f1b932ba729d3a81c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71f3f9e4fb6e0cc240b96ca1479fc2e5f5680d9cbf7768f84a5ef8a379fcce6c23dc47e143087a915bf58324e899530c8ab4faa50087e0990367af97032c59ba5dfe10478f08db84b4cf08e178f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ce4f0e623b00af1f682b9d306230c50210efdc8ef93e2d1a900360b08fefaef5eabd0fdec9485d7c12a967c6a44dc8f74b322321f1387971e58144fb847a0ce0636115c1515e20edb8edb9440d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad14526cc10347af9ea8ff5f5037357c7c48f07a2eeee16924965e2655f88c04a902cca27e65bf3f91304a5062020a5556397157fa4f6cef0be91e5b57c262c554c50de6d3eab67b443bba6105e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c10ae870d3479e04121537dcc2c3634c8cf8b5ebbaeacb0ad7c4ed921d3a152c1b74709ad5e71afe4c779434ad3fa2a2b20ac5d55575d618775931bc6dabd3dce25406a038083f3f93f96847c14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103c8576ee89a6223a5cc237819bb8bd6d98b6e8435d3d5b0c5a2bd6cf62b400e626ea59220586062472dbb5952c61812a4481e35b8ea2fbce847c688f3995db024728f3e03329bb34677107817ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e3fbad11173f9a696830aeefdf2edddbf5425ec3676e499ddde0c06f091d753e68c055cd54b8e0085cab7c432e9e00a6f268bd9c47742906166d4e3b6d0df3a92cd207b1f9fba16c517fbd52a8b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab0ff131b027fbe9a253c8f9e5918468a9298897e41fedd2464cf48d74b0a0e9b310f2d5214a02f4615351e759dbb46a3e613ecedfab472b148074dfeff3ae55595903641db40fe4d1237349e039;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166f3d79fa119225e2e8bf4bcf67cf5698c601303f41925bc6a687d4e112343b8f043109f4eb03f1578e18c73e5e2e0e4145e058753a80df97f5975d9a85480583181aa468215e14d923c18a1b848;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37bdd5226efb7589c34da5e1ff3ea1c2f90000ab080cb9dd00defe0573befab79aaf2c9819326d7cfee277850504139af9d5819fc84b71ea35456acf519e30b2a9fd56ef4ce4c6ba5515e6598ab4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d59a4fd8a8954056061495cdce437d594a57dbc65c96d7d92d844a1a247e6ff1b01934e26e0c71b69e6088e70f512e8a443fddda1d2e919912f2167f4acd8ba4342ba49210aa3c2fc9c136baa78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb09c14f92be01111ee378239844a7baa4094716b2be6d79ebed4199f71b1e120f1402a287b8e84bff21a570098de82d84fa3cb659800f039f3317bb641aa594679702aba6bdd5fc83159597fa09a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1853c341923210de2f890f4c139eb40ec14a644354e1b0ca5adc4d35bee46492bf6472ded8094dd13946b3878bce6de92f21d1cdc59a3d62fd3f08d6caef7205b38aab7d581217ff82f9ce9425ecf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1cfa1397d4c111e9d1984cf4c66a0638b176ece89e01a31da0eae5b8eeacff03ae3271c84d7cfa6df7450771eb10ab2a2dd9824b965e0d636d4abcb76bb497a984fe0e04ae6216a02531d1dc88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6110be655abe43fc6851974ed8069ef465d7d44f5b62cd72e6184b5e9c2ed2d20b2d517eb9a57ef3b50b464a2d622315fa8afd143f55de56c5a409c995bbb918d7ab3f64cbfc0c13b5fc7cb0e6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd59423bad4ff38d7919a9b26e274c456606a9bf05e0e2eed90c6de010216dbbd595a51ac670d7b8a7d721efb9f127bef6daa03d59187b78712a6e49283268d32d079b40e8b2a35fcbd4ace218690;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2e90858d2fe6784e55b40ed47f24cc651b9e4691fe6ab443ac4ffae5cf468f2807a5f42f30e837b8f8b0be5fa167f05174a19b4de2d23b381b5752669a9a7d6106f70f852fc004072bedaf1a93c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd048982f67122bc49137ef2413cdfa64e6dc1a0764ac8e53a8565c3e46ebb924a69654da1e4bda82408199b2cb5114abbd8394e26c922c768fe953924be96979f1543377f90ca44391996659cbd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b26a6953424eeebaca5dce0c769382dbf21ea9ca991690b2062900d4f0f27039c1a6178c94c0f7bbe153b7f5e2fcffcc198d1dc322b879ccaac069485426b2ae517595882f46c2947c16b995d196;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4891fc108bb64f58b8a704dda29619ab501fcd36ee1eb07c30b8223055ec965916d67325b5154bc3c8f421c5f9d5725e2276f434a67e4ba393f8f1fb0ff8e01b2cc97a3acb6ca3ef814dcd9826a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91f1cd75cd8684fe73c91e76d69335fb5b140e53fb95ba38a19a210d04ca26b374cd88c5e11f941a7c0b1c733a804eadd36410de8d16c805ff358a6d8f7769ab18a3e08cfc169170d378e2a8ab19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h546bc3547dae126e5481fc516f8cd4f4578ff94bd55dff81034732b9f3c4b710354c9a19fef1bd0c57dd5ca88d12f4ec346a410e5e5787440c7cff2570fe9d5a09ac1999a178ff6a3fe99671ff70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h881c3e17fa470b3b7b29785fcc18b2627ffdeb170f443ee620ec7e61921d17f2762bb5c51b8d5f1fad306bec9360297c08f9d9bd7f7ce5f31ed4cd5c32818f0bc7135e13b7b3f8c207d1dfc196e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e9756609f73973c818a2fde8286d7f74206db1ec7151a135de776b493f5c587d10c1391d623b1961d4826e4211c02a7b662c13ace1bf2215e3e60bb1dcde1af4a885b04a340aa55245d7e638c97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4520ad6d9884f7c687940929b5580e47048ac451d7494f5a9a919ebb8b672d4e6e4ceed80a497020b8d063a0d363b4bbae7be8b862561a22ea1c3aad990692f11738267c92de5a42e7a1e3f1e78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1695164f0f3cda565b7e219420d083b797cc4b9748b71550d1c0e2735329055cdf47a6f8da0ab88765ba2b109725ccdba38907e071e6fffcd1519e3100674a54aa43c98e22d7b629dbdc45c4d1091;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adc6922dd91c9a176956a4b5693ec17dcfe633ddffb691129d5b50ed371b7ffaeb82ff0e023b7ae1b2ef87d5a1dbb72a4aadecdc444118b0df032091fd155ef23cc4e5b486ae8946f279a284aeb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf1ca35c7d4e0a2572ac64014d13434d53410cadc64b30a3823ba09c3c0c5df174fcf668f6ffedb59c57dde5803084c71bf2d57684912a7596f05dd77d7e7d334332b75ce6fd198484edf389776cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7aecbf17b8ba667937f7d60038aef0162281f436c6c2d987c16e36051f26724c5ea75d49da1ec9924fb4dd9ce7f513696af5a9bf6a245c13dca4b84860d0141547ae385f13e7773d0ebf1f7d778d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he146eebd092cbdd8f5a6481f2dfa4fc5815205b97ade6f9227354368c5e012a8db8357b50b86d2682d894bea6981e5d2df3a0dcc6f9de07bd56e0d2c6aefcbbc700e2b897b5f4fa10612807fdaac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180a5345fec0247a6d00511294e8e3e7f6f501cb84111025b1dda409cdf6e5f0e33e4ce709aaeab0e362055c6e201252fd07de790a2beaa599c6a56c4b9b6b7f2140d6a51cca229a1f91cddbdf64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0307296131ca34f89c789759c6f23dfb1f47ef74bbedede307b5b193f5a2a8f4606b338d9ca0dcdc5eb35af35f3d1cc9de60970ea496c4f9dde7f95853d1805cb281192e497e6a15666d45a20b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0269a6abf5477ede6899c32ce282070f9e0b86092ff7359b71c06fced892ed79d68c1f354e5d2b62d94b1208e276579e049728aef9d44074f3c77d0028e12c2dea176458426c462894edcd29bb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6dd9e13e1e7413d4064f952f926307619df7b6814cc81769e69be35f8ce63db99f23d42f30ef076a611ace22f9143fb6736bc9b38a95be9a4f29f4e0b5c23417b389f796844402ade4b6d93b2c63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ea60ecb5c9e8916fcdbb7f9aecaf793199d8db8dd49100c67294949259faebc28f1d79bc18eb371725724cd4cfd37ad8b1275b150b1e1539513cfc645f2c7f925b1c7a5499bfd0ac43231a98e97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1477ab5e3031f27248b8ec3b2b3e2b2075d7174edb5b175739609d9d1114c8f5f1a5aafe25222a402b6df4ced68e632ddee99e76b19348be9dfd7c7fb248ab1f31449f8aab5d5ecabc840d0aabb65;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e9353dc6926a41e5f27b1c1e75d32ca4b3ba775d4bbc3b222bf48b02ed6d61d4160ce76ea90b6d045dedeb52082fc251fece053c5fe0c01c46b9d7cd4b1451df4b5a00d6baf7d5af176dfe3555a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h585d2269114093310478d91b95695c45058bacbaad68d6ffbd99c7b137a04ce4b9fe467e115e118ba5e1dbb1b741d36ea9b480a1761ebf656bd5a3b939aa1f2e19ebd7df3b4d57733bdf0ff8296f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0a53bd5f1edd90cfe33a13229d4f4117182004f368d31a4bdf7496718966b6b8ba71b333103231a891584c42ae8c1d077e1bace0abe830c80d400d7177434e633e5575e6c2f9de57fe7987cf09c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1746724224d344e3735e2e2be48763ff8741f3353d41f808a0ecfc90bc7431c8194567de9b7cd905156c1c8032004162ba673edb2a51cc09780113ebd21cc788ba8350b3e8d2741659a9c08f3f586;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd61f1b0c556f5db039846402f028fafefcf336363216696ef1f8a48491941b7670d316363911db3d8ef4e04b38b6ba7ad9085b3a73cd8bc58ddab7801753d09aaa10424bc12b30e513f1d9fcf410;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6592493cb27da7af880d4166160a934430ed7a83841e8da34edc4a1043b57fd7b7d4704779eecb219a81770536325461098f5eae61758e8cbc30ab70bb57c9737494f733b33bb2e063a20f89b77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27b1c2dd9e84b7af0f814d30e6182df40ef006103c87d19adcb0411b9b74952eb1bb650c549482f6499e1d4b0784496f98cffc8e5514ca794a5b63418902fa58b4250baf52bf21e718d0249709dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31e1ddb3faef4b3fed5a1b2ad24aa6ccbd5ab2acd9cc8b8385da3838d09ef2dbfe5eae2ee012d09ca0f20f5f3e20cb96735b35aa120812f46c07d97517444944fcc94f46e917568ccce3088ebdb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7879f90941c2307c007455c1eaf317af1d1d3b818b20e1b907a0352581fb5e70ef80bce11893f93e5e06658c5a74d634168efdf1cf2920c9b5e92b7b9570b111965105ae4659800801a961b4204;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cdb11c8d884bff9805fb26467218b1e80a130d725584734e310b9ef8c85f1208ed4d8af2dc203dcb95a0643b0b32e99ea289e749cbede4850e6901d17e76942fa2b7ff7795e9442b4e8016d6318;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5fcffa7e94a4645fc71144bec6ddc0ead2ed6591ff92a712b5b417784105442454ce4ee9d466aa0f0f741ca927597f54e55d4162f42b4a6531674baea7f147644dcc8fc3451107a21eee79da869;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc20c8148d3356ae1dff50c87a960815bda0994d646868777c32488a6ce67d4df2a691d788eb9909e80708cedba26e5d81b5b18138f321b608988a927c04dd84d586fc9100fd82578c96314b7295;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c38e1a5ad25fc0f8b4ae80938a69076dad1e114c9c6d5d0cafe0b3691a5e323922ca22aba19ae2698c69ff7cfdb2eec6c4ef4eec94909fb7d370edb91e2f6dcc33cc20bea27b2b9a756d9c6412d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf06e47f9700b617616cd57b06dfc73fde81ad91fb5b88b20a2325d1159ecb5c65d3d250860f0206cc26879334efdc172c22f426331fb8916ef292ff3a1b28f863d1164dc9215886864ee438cb00f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f39f19a8522847d55bb6a151420513f3de970d3ad68d7308fa61e7c0bde2f436c763bb96e331c02cce89f9abef17a4eaeb12cb49217dfac0308fe2ad15ae724f5d73f011fc05504abd777b77bbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154adf7a4147e215712374c6e0197aa60adf8604169b7abdbf155e88aa8dde3881dac3ade0113b5fe9fd2dcaf9da3bafaedc2f7400213685d93c7b594caa0bc4c6c18010fbeadf987430764ccc0c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137403c077f83e736552812f6ec07683a79a52863164dc985b718c42dd5ead95b7a64c740c93fe72a0d4d48a65a2079c327cf35b016c917a31e4c15636059ef50c9106f77b3b440f0af6bd23f88c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca52b88c1bcfa39d703f00d93116a778e45037d0f26721a5cbb5d62c32d7523a6bdd6ce7d7440f1483da7f9cef0dbc991159a59ba62b4e08c0c238746984b740c3d0cb0e49dd4838f847f3ca7b31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88f7c2b1ebc763f680f31b4fddcd6338c348d56440caa509e78eff915f2734c32e75cb15fcabc27fb65a39dabaf7e4bed1804f75ea42b89fa974027ac0a966ba6e1e0b9ce5e38ea677ca9fe0e3c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6a66b07a62507d1294cde20381cb94482f822d23a511843867fb513ff377d7b3e8879b78fc46aef27289bfca17d9e87fd1e48d04befeeabd5f8a4e614bfcfe7bef7befc15956d531e91ae5bbad1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4012911610688021d2e618efdfe509a079d90e71b3670933f0891d692f3d49a14bf0728f5ef78a156818180a724a9fce92da8451783f44ff09c449a17b50c54d0a135b8aff662acf9bf6eca2d194;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ad1225b4ff4ac4682ad13717af095481d717698c8ff1189e64ba18f43e4d647ae61570a47c49481e96387af6674a5a9d3b76dd8a3a1b2105b5078bcca3bf7fbf175477a4becea760549a7d3b09b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18561bc02167033e5f7b35cd4c8e8e477c3b6495770f31b3d58a31b0b92a0d1aeb9e8b23257f5e9d98487ccf13a2c66d811cc15265ff52cde2006639142efc2695e777b256cb1e4f13a3a08699ef7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52d0591d14c95064aa5ab639ef165e005c6ce1d48b94ef190a8dd5e85ab1e6ceb21139450ab614c264565654e24c59bba5f1dcdcb8fa5730959a659ffadf6d2dd4b4882399da972fa0ed7c49043d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45eb798ac53619fe786f9dbe5879c526b158ef78f8ffd357c38e5d16724b36c8dc395bf941a50d4ce0ee53af109ddf535b0ee895647f5b163535c369c66e5d3b69aa0f2b229ea79d1208aac93e48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f8a89c7335aa3e85211ad9a0dd54220883fc0d42c1ba933739a6a1a17eb3678d4f747df6eb952551d091d612dee690bc447c0e4f8d87593cf58e66c25dfb9d6e080df1f617b99729fc8510339ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ba6dce146c23cf28ead77829d8605850bb0e505574aaf34b2de923a662bc74ecdf64487fb50c633afe29a7d930ae0a369efc3eb040c2cc49ef886cb8f9d226eb4eb1c7503832beab86f3086ac7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcb99e7811e6a3132772ee4989cd738237c2241384f8d9cdc6c13e20bb0763d0661db2ca5cd7b1756320c091b1fec88d31956c44c4a53aaaf824196c93e9a5d48aa682e099b4fe5e866bc3802ed8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198c5b3807b870195beaeea0d6ae1308ab760d95460b2f123e746e1e904ada6df80a9415d698731c857358f3ab22f10d9af790c35f3ebc532d7871f013e0f2e67ba38496ad1b6ed5900bc6209c10d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1128026a42571acaa249658216549fc1cd858f61b8b0fb07cd76bfb9500e12b5bd529856bda66c080c420db2b0f94545242864ecea573c095baab22b9cc26da3752bec1ff97620a8289b26383dfaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6fc8e15dd6a5901e9f6fe58d0edd619959c84da886320d7c444259aa6662389c494f9f136079e938f7684880b011728f16b5b15b922576c6f2fa884bac8236f9db09ef5e2098881b35659e663fe7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0431aa3839837b689bff45ac8cd7d7340f9cfd0c8aaf0186d4743b09ea63712a7af346860750d1996039588732556b767309d7f1a267a792c75928bcd72c5acf5dd1f19895e26f1ebe0f05ffebf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c74432eace826276ad922fcca8933670805dc42f11a67868f871079a45cc570bd0ffbd2dde513d08db66c7df25014aae27bd3429d76a33b44e1f210ab06205d1e8752ced9c248c1e86d6f6573abb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb610acbe1c3b59bb694d9ca8df3b7f83a9dfba529adf539746a6e0b7f96dbdd1aa0fc675680507ed88d5810f179eab851bd8c7435be698ec3a8cf0cb5c153019354daf26b82ea7747da8b55a697;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179342011a32f4ede5a0dd638584a2e54a399da54e693eafc3df8be90996f4299e8a894d02f6320d0b460f7108cfef704b455b8134ae55ba3071fcd71c8b68345a4795e25fac481db8999def0f596;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1544a675fddf2e4535fed4b78ac744ce7987f852b30f5dcb51664b789e1610c1b68550596f9bd2762644ca44676c1027d9ad61b1410c26a5d4049342dd137d77592f5489ee61b4b4397c2fcfc8bdc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120ea3bbd86eb30214ad32abe16509f8d35b6d5a7caa1d52de575352bc91210b6f39fc51191fe6a4abf3bd724c09a23c6171a89076e8e27e7d3112987481476ec653fe97c41c772cfb106c170d26a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1362dd2e001e71f99158f217eda7101295ea3134c17b6a0c1bc37340121c64e3811d5e4c32779593e2b9519bf19786b572f72eded9538d3d2673412830053ba1108127ffdbeee251547d145450c5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e8171b9fb0396ce7676d0a52de7768a13326cc3ec9059b17b14f2b3fa9b59ec20ec9e93d82066b0483a114b470b8474b9c149ed4d4d5c47a091fa18274777d760e03be6a0e74444ac59f5688573;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h920e6a7823a808a6c564750c7059809c7c6e2976d4d078d250323d69a0c40f8c44c3870391cdb7ac18121e1c44ccbc65d8defacc1e93ac3e6485173b9057dcf81a75066ae3bee84b639108504f64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3877e8501581e9409a7102b1d67a4f1eadf37c558a7f2b3e6f9b5f287558f2f54f531887f203147f85fc3d41b8695a37e363954e28a305c7c36d0836ff2816cd8ec2d929a23e60772d412dfd156;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h343748bb66126eb1e366b44f765a558572905a05dedb329109a97190b7414718365d4209ae277f66e6222abe17cf4beec38f36fd8a010269144d39324f0ec146879fbfabbe5580b39bc1f4823e63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88891715bd408d464d5f29081fbb418e88e8e53993e0ca48ca16dd04da0db65cc607f627745fa492082a8303b9996468827af5a5490ea757b8fab9c777fdbdfe73c958863b1079c2d33e3e09d2e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97f0f20beae30671602ffbca3101f44157d7609e23e1ab85f128d2db79605b3a9d5022c41878c50eb5aa5be24eaf994b708404855a122c11c0ec64de020cc636b05a8e2eecd598269fd10a5fb66c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10aa6ae6004aaee5e548a908e61fe29ea7db895ee3d29adf9f401bb3077ec28819cdfc9dd6c7c299e59a04dbe59901df59800079cd4473491130ad5d028bf918b77eb331846bed018fa3939d4ac18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55e8b82a51e06b8f01a75be067885775bb09421c285856eb5807a8c5ff6e8c0c00525b48574453c6b8fad8c4140a2892ce4b9e2b5506180cdfa0c074a25396214d77269057c0983ff3cddedfc73f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h758dbe389d8594d92be2b31c9b0bb35eb5acd2a5fad6a52334162abf4426f31e717facfcaa072baf001f9291b75c8356b2ab832934f8d6d2f641ac86d91407c6f80281f521d7310021fdb1531631;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d211e2e6c6c28b465547fa1abd7ad4f2833185991e84969a232c42274827a53332fc924447e8a19d8e7fb8c5bbe0f8df7d2e1795f3504333f133fbce75ff679cbd532ae086a6a5b66346b4c2f9d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63951ed4e94a51df0c09d2451c4962d0d0466ef4126ea1f26aeb53772a77830529b0775f11ec0622bb2c230dd62e721cbcc0c9a72bf0cbd41f5cb1d80e238ebe89cf30e71cf5d43e039cf140ab1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fe10de74941081efff43ece203e4c4352d9c249f5550f8babbed7def18e4166fd6e96d8878ccf9c1da7fb905c9149a3f870be10f9f3acfa9d4fc9d5eb910f15fc3cd001b041842b6c8a341ef1b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1839c7c75094568ce0b99b2e2bc8ce2b205fb32350791ee5ddc6f59d6e90a1183efda6a75e8fdf64a710cb4438038ecd1adf90097650daa92a5b6768b180d9e6f6e9676ca50295a69fcac92734b4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bdd30009b80ef3435a8e7bdfbc8aaa74afa3d1d22252ab1bf0193691568b63d9ea58529f55f39e2f796fc3854faf573bfa6d7732d8ff5b7e79f8e857aa410e4fdd90b96caeec4e1300d3a0abf7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h217ae783498d8a4254b4d30deaadde9bffb54086e2a987746e43a0b358a939c2dc11726df31cb6ae506690d3bef7111f26c2bef8a068ed910e49acab7bfe1765c37e6220480b3ce12a4ebab72599;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124b5937c31348f9c53de8099242c2726ddbfef76ab7cadd64526fcbd99f933fb1ed793315a44993ad68863af8e77bc3375f7cee0b40f5f12768e9d9d4c323553a13da6cc55a97c1b89cc3dc686a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123f2fc3e551f62b9d2e46096656d2f09fb9c83f2c51a6d7bce9fabcf9b7a1409a804b58b4ec30f92e99a102b42a8b4cd6b3899e0b69e308d00e038b32d403d15ffda226efe2df7989fc3f7ce0cf8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h982b35770367f2971adc4a22d0f7cc27f98561dea21a1af62685247d839432de088ffe23a679566ce1cad00431cf470f5c6c9f98555ae4875127f71726a98aa2f27fa0f9c6022e8aeb07c1faa22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ae724ca977444036998ba8c38389000f17f0e8d9f193b9d281c6e9c3a562e6709ca83078e71adcc79eaa3a18c0414f0ba028bd5b4c4ac961b4b45fb8e4a1e9834dc2e741c7abc3d278b058bb73f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0b806fe099d4f4f579e9373ac6039a21ae7dbe10a7859014841a388cbff1648cbcd918fafe17b53438bd6bb6a2634cf7f366442898497d6e82b68306ac868518945af077a68e180705fec982203;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173bb185a9fbf28db6898cd460ae1dcc3894e8cea79d756e34cea2e0346e0a235001f4924be058a8fb7509a07ef1e64415e458303367af15dadff20664b2627e6ec75702e34a21ce6d927f6e9978e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7527d101f83514180d6312875672c4c04d7ce801f75de87987bdfc29ada08f73e3bdddde0656b758d84ba5f9ba7f8d79c94cbe279af808f4165011c42adb5432a9c2d374c9fe8d035985e4dcf66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h853b4c79c917c87869ef83093cb3bb11b31c687b5af41630344b978530ce2ee4899cece595ec3c79a5fb300f0d0bcddbcbbd0c5e0780496b70c0728a6b1f3fd3182edeccf967a70ede1530071a75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b9c6a34b46e0a374084438fd5c92c484e718e048a70a030f329d962afd814798c45273893dde2cf2f4206483acb8f38770ed64f742405bca784fde4d994c9d56ac51dcfac58987f1b36f9d53c75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141b043ca60a6e586371bdf232ccd6cdc2a48e8e480665884fbbb047b0a39779d9cf993868ed2bcd761876f52d4fee8632d7731bccda92141ccf5daefc2d5b862cb7a3defbed715bd0c34d147eba6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f399faf2b0f2fb6aceab6dcbcef9c3006df02dc186b9bd22216cd92fa28ad992c0e448af4e9326c71d1cf223256d897f9abde4de51069560623c1e9479381e88a2b5a2ee97a43353f31a97952f8b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc21de69d9bd3cc264a92cd4c6f3257c060582ae83e1fb5ea5f3c5ba295230a0e5b24f5e65b0e4f656875715f48ac4060aa86a4d3df7cd25f402a3660e92c9a8359a10c593c73090b67d65326166;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddb9a898b6cbc06282405b8df16a65408f2dc149135fd7f2ca0a7257561d757751fb9478ca7e78ee5d59457634a09c8f0f8de89e74a31f8bcb7b2a5922488c259ee0392740d1e6ea926a3caa55e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b43f1c854d656e34276b41a6df7c8a0fa67b4ffeb23fcd28071e32ba6c23271e94e817edd28e5bab81a1e2a3ee670722166048766a89b064e5692e065cfd754087e98a408076d96605e53c9e35cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47be92055f17c61cf76daa731fc0083197ebddf427dc81d3346bf49f31b4870283683cc962e0d20e5704e56aa7ef80e6519e3b181c6706cc43b822ffbaa6f3f24d26953d59ffe19bac97f4e52d45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcc36cea6c5d0decccc0eb71eab3a84a2efbb7da59e8d0d925edbdb13609d6a39ab47e117fffb76ebd904c444f639acfa063b19322c8255f7c8b56b03ddd439d412109ab32ffd1d068a0533864cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1d3c65dcacf223845cc9afd9e81cba278150944f4e69c92ab1ef9a32dc1d11e8bc86489398cf93879f895f181184b3ba9bf08ab8fe5e92bd7268f2e6c17012697920ad33494e6f73cc01dfcbb79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15aa2521920351978695897bcc85879ce635151c9d5627f71bae5de85072ecb498a79cf16b412ab25e509997b699a8ddff39e8ac4ed1b9bc81c8d5ce07b8440a64e219013e3f7b7f4ca8bc80aad99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15dcbc2cfee8ef5f55d62a873507ac12487fa3ab1819942d636a850242b732bf12ea71b6a606f0c16afaadf7b96499633b1d8d300478bc2240fda50793f2e3c7dcbf643fcc656563a82a9a21ab603;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce6af5de56809b34f4f8e8a5787272ec85acd55cf40ea20e066e07528e7ee022b3b6ec82d5af3ee2fa082a3f4ef84a3be21470214559752cfe96ed79e4766284219f5965c2aecd1ffc5174ca9dfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h788430d7abeee1cc8e8e3f25cdbe95c79a084552b78dae2034017da423aeb52696f2dbc7248ed157b1205a6ec9ef61bcaa7be0a43bc0e6789c40238ecec38d275c4568f3dc450d0ff91e1933bec2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afbccff178c1bf96d4fcae20a1098149d6ace02dce1d71cef061caf4294f6cccc7b4cd9512d2f796b66979d8c767572531acba963ab4dce657ede4c9feb77a246b867eee793fcc1d730132450e58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bee24ad871bec29f4a9544982cdf6f9254b4e7f746ea8f6120739ca1d05349782a77cab406836301703ddf3f5ce1ebc84acb1fde49194ff7e40ed5a50be7eec2f812608756e15c0d9da77e6e5ef6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78a235aae3cd06efbee54b437f2e3e13d12d06fd141dad53e447846c80841967d2680f04adeee8a1ae2cd1cafd782f973341dbfd81398562a4eb3822c34b4f2cbe4828c177e6f0855e1a1ab9c6de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172da4a678c2eb6bfd3ef316fe9d7ce7fa4169670d99ae37589bc1d1bf427aafec10bca4a1ade3aa10ac3ef6b3930b2eac4a140ffe98ccd3622ba85a7a8db890041bd00c76aca754ddb6ce7c92c1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd04d2f7fa47e5d200b7da024fb6c4522928a798a43670e9e43edd85a9057d69f535f3ca820ce6919bf803f12dde2cd2b6990df21b4df8b4d94f27ccf5cb13b0e20ec8ead6bf3a238bfb61fd45050;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc56d1e7b1af332d74f0939264a773d632069bda4b4ec889aa42c4c0224a05fdcf7dac3aed34085b57be17231bb2f6e7fdc7318dc980dc6ee91849c50e6a2f50bea27b6a1d44d749788ad9f2dade;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b77687409018adb36784390773309d3585cdbbc6181f90de657314d958cef25ffe0a27c5da0e68cbb602809b81e53f0232f13416df28c8800ecfd98b0a1a3dc8600b7825e881b3a57bf36cb5e3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11fb22f37c6236ad893a68b41a3a606bfbe5e8c755a40dd0c22270460e73ffe2075e59cb0471cdad65117dc1eaa32073603ee950a62b553fcd823140c4992a4a44c9253da836d8f313db028082e5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h793e613e5f4d9e415ce6799d25ac41fc8eb58911b6fdce68937c4394e555cf10bc9d88392bd7e765451f31a36f96117a3962a9940b252ab53d7df66356e66d2a23dbb1c936a078eaeecbd6b3c31e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b7e8cc52431e24af364df320fccd1bb1165c1ae9c1f059e5b0ff8ed084d93bc9ec40998ca9518de38593afef24a4b592e2359ccaa57a6d3f88c56d071d1373adbc8687f4344168750f9e938dea6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2277c785aca64bbb0617e0543cd9317b7ef6b3352caf7fa6f3e86a124b171a3c2dfacf242c303f67e401e9a2e089848eb09a9bc3cad07b72548f6169bb92c2c3d058a4043233e349f084cd46d257;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54ea5eb3dcca37487490b022777c148ae49ddf850e1e6fcd2ab534886f5bac90f81a41f61afadcc9a72bc62c0e76adcdb9e67177d2f03e9869e506b07722b9e0b6da14e07e835fc2d3e458582d1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2193d4c7d12e1a5e888754cf726d184123e677be52110fab1a0caf7961b28ec39b429e99a15ce15cb1e217ea67b213d7a07777ae17406cfe9869527097c5f53bcde160645af510795e5cf234b0c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c1bb8e16754df7de581ffd61565322aa775fe57a4afd4372fe2fb4fa0b65caa21a65af1cd7ea5c4df4eb541975e705a933bc73672f2a354ae98c0d7d548f950182c4172cef981aa73ae660ca168;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4be68dd6b7e675c80318ca625961ba06d92db9c34924a587d1ee65816e43ff5156546b90adfbcb273f932e87f5e8bd0293c6a3de4cae271fb8a83806de9aeb71f5cfb65ae498a41bbe0434e1e666;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24e4870015e46539d38df506389883b314af4cdc9a97692487e94843689ebddddd8ac75348cabecf073d31621aba27a15f8da80754024efdac0a275c6a6cef26ba68fde87d9210ba4e61720e0e95;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2017fd712a9d2a9dfeabecd0d9a4f7bfa6228ff0deeaeed82800f4c07fb5a7ed82f4aff4cd6432a08c126614d8fba2b2646fed1d77ac76d22c83bc0deb68d3f6baec960e7cd01d045e15ea5b009c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7dad2f7838282ca0643d454f9e3998009368359884f50d5b843d0d96191625dc5736542af120983db7bb153b6d6325bc8a5428c100e0d11ff068a6c6ad796c87486ca00cdb040355ebe68cad5e1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac3450bfc44bb981d6b62a2738ac4e5f3ffe386b54a83010ff0940a01f7eea8e9e4e0cbba25fd097166e6a865c2109273b93c1964137f70bb186071723bb99f2b48cde823e77ff94997caefa4211;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9451d71c668cbabd033a2ce4a088dbef56832898fb844d35bdaf50b7abdd46071109ee5b8d881e10a33871284c044291c61868c7399f41f154426c11b83fcc8d4727bdf954a3da061d4f833bb29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d896db87bb49a6d6d16896b81851141a982fae76cd2eccb939859b55e190f7768dd54702473e0120b844ba8d4af1fd6e1544aaadef9032ef0e648baa413426424b7d1972cc20b85ab748a1ff2c60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c5b593e9e59d45bf781ce9fc2a6b30a8061325161d8f958b0dffa8f74656df9d1f3e35def31c65032bdfd525c7cf00f3415b8fa26d26df83a6499aa282b9621942aee6da79b6ac5913e8dd9f805;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3481a7c90956b053b0cd6b890be4f856c0a1087dbee9c8ab582408f4ce96bccb286523486380a6a2a41c9d9a650508b7569661a3a5f6e8bfa3b4fff69f7735a1955e11535a66a53bd7d4669d5f37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1918ebed820a5de5ca153d8d18325c920835558b03bbae9e8da818a5c2f3012744d83d497adc71848822329479b17b2b0c74c9fa49f62d32840bfa11b5dfb3892d079a527f8cea4ada68e6bed6a93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b46c6e28251afd6a3569dd112706b9b8597c7d69d03adeab2220da2507badb81f1c4966c1dd397192bc22ae5804c05cb243f4cc78448c6756ecb7ed6c1d11a458b6b9cb494604dc005948911a5a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae1e69f2797882022192e623f3be54b6e3db828d581d3381f32a6bb334186b296bc318436e6a0d1adfe9f7ea2293515a9a0160616a1371d1c1344a5614ef212ca5537e7ad9c1fd58bb12c0e3c451;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he30e946281d5ba5a93230aa44cd5ebefe91a647174110c9837fefbde8a83e46a85e29580f81b75c58abdc71bd14f952cf61e4cb09137d7a2608cb3783fac170b8333cfe7e9853f749a0e70ae9bf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1282928a49f36f3d551708dd986cdf6d0b693e84da8d6c99f318b973ee1c394f94146358242b2953ebccdc2cd5f0f2748602a8b2c9db7aad74b6048171e3f6be2b1ccb20716d2f366d61e2d210c57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26fe36f62e98a85bfd71a38687a8cedf2129a2ad7fcc5defff1732872085f47456810e8cade4c921f67b24f0790449283df3f22e71e061486979d5024d2d23fe0e7a9bda061e904652367195265f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e7b4861e58a016fc3cb3e6810d94e8da8be553a394798e22a5754a0d87eb104b5f7fd5597b4414562479d5e7a70fb7f2a2269470cb54f99193ee1b71cc86f156096d400db65326f73adf343b2bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14092a59ea11d09a579c18c1f375ab4f29a73c473c6aed5058764e7b1afd6571118d6c96897e5c2cba673913e171e0c151e0165a013af72dadab95355a7b80315362d28f0f735864122f47aef343;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8a4e4a72a478912f6ba9f1130b5a524dba26b175d335df77ff2e4cd8980f3cb1c13dcfc1e90838b1ac69dbdb917070cc4e97100b68cabb050006c6951b3df9f6c879a9965db99500b3056b63988;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a8d27c5519a3b0ef0a0c91824dd0f23f919f19b7218cc0c62dee3485f67c83b30c4dc384591edee564176eb60d814b9cb9eafa588d41e7b287d116d0416ebd435189fa5e9bfa2c03350cb5675d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157bf8ec439e39aa99fff1a7e4965f36e951548b8d86c646ac64b9ef22e35fe1d3d64284c7c76f1751606c45b559409df0a6a9df7af099db849ccdf6342fec769622016694b76d2cffd58a6aff55c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a9919cc277e68a1c2ee58a39e96997ba56181422c172c47186a3a61b20345500d4d3e380383e7ca0cee80a5de65f74eb6b10956b9a8503682865a8e7d39346b7746827ae94ccf0a011441ff2c13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8d1a4349f9b5ca04cb1ea95cec487f5388c294f858d064b989f051bdb628ab7ebb3e07eeac4eb11faf7b2b1dcd6583c8eeb2a197334be28f14b744952283209b5ee902ce95b945c7301e2e87d4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35ae2e93d004be5180d4d32a6f5126c4ed5261f8ee15f83acc6c8b360dfe5f1528cb63229af28b4db8e7ca1280b70bd19ad62ba2b0b7847f3dd88975be0d121b97d00859bd057f3dfcb1d32fdcb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e312c9c7e22813d2971e125c12da89988a0a2d657eaa9e3e932e7902ad0ceac0232a4d218bf3d563b0c1b7db279bcfb2b23b4c6530b307377a81e05943928a6910567f9123eb5e2b3a8e5050f284;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a11eda87e7f6e7ad109ad2244fa55ee73d1dd9ec2018c66784c82368c58f119ca11641e8b20c1cd09d6d9c604936a0c8c3762d7ab5e95af65ec8303195d830e67438aa0f79745cde34ba70a8266f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbffb93bcb986d06cc77373687f3f55238ff51c68f84a1428efc7338512efb04b4ab60d27aec6c5735a2d2e12668e639b61c81bf548c9bdadff9e2df9ef43ed275349af9f7d72827d9fd311839c56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2dde608d648d40e4d0827b89101163a671683b03545f8ea843eca04640f7c5bf685effe67150d899526ff512824f847eac114a9bbff5dca4e410e6bc273d8891953975b619583edefeb7b72d04d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9291268ebdb0e79f324e4668f30ccfb3df529a8b6defb2371beb638ecc8e8762245732391abb89db23df48e18024b55c72e004b4c4c90d8f16c3ee7810d946370e268ecb1ca66417d68508598287;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31d94d50ef669d2c9ea964b14bbde16e22f85cf0cf9748ce62be29835dacb2526d969a932144e5e415321c964f876f84ebbb11b8d74a5c138f4509b196cccdc72f3d3160e97ec1c3fc3d803d57be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha23db6f3b335b7df83fe5172f00b60fb7cc62d0a7cfeb8976ca625f959e88cc3940cc8c6a660f397bba52725798927739f89baf0c3dd1bd81c5cc452a8dbd9712f5df095f6a0edcb962386ee1d82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e81f71ce7bfd26e295d38eaab6fe4b176123b394f18f7468f422cee10056d4c5abd8592ba83f6d0d9bfd3bbed4803704cab216348ea0817ddff2330c65146160be5f3c69a30828c07f832ad74bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea8b2b2ad5ff781e1a8090566558af0d066444aba68fee6cae28ef2273f62320df7c2c877ab5e152dd9e4159990eb8951a409eb4b2d0fc53d40465ee9b7784480f3f5dda5a9f1ce1158d59b7ca7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afd0a34addc4010e3c13fef9dbaa4a7cd5ef519060c79702c349c76c53f056095302a2eae718d4e7fa6951a7158512f3567ec27af5f5f6c912aa756ebd3fd18956a335a659797edc431b78765f05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137e877b0083cd89925e8a030933c44bf202d7ec4e0e39b4a4f0984d787acb63c0f68fb34a99a5ab179adacf25a63bebddafaa876b104ea55fd2b15ec6fa3eeabe79179d964034d08fced7d3352ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f2be2ef704a326cee06078b81f1b8ee4fa1161a65f415987ee6e9b978d0ec9f355d701e15ea7bf4d08d757501200e67537ad1e5989c397f53a4607fc96493a84a61e0d3ce5046f7c5b9070cb36d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182824dbfa2af40232b0711d42edfb868b338e516ec83324c4e53d96c9d055ffd4ba3a9f1441be19a479d413a28c48b5a7c9a28dcb5b678b7a6128efb82190ba27d6b0369249c1c36dab03290a379;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76451572666de10d90c799e691a6fe060f365ec03134d606580eedba0de6ff427b0923841f52c9ccb63a964dd356a4048304c21a4757bc0549130465269386141aea61d47eb3f2b5e61145fd39c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4b663b5c90a51ee5e71a390a4a9879aaa78ade5f519b558ed1fd3a1e20dd21e1695e09bec41bc3426b8a727f8d425bdf2a34a500384d9ef0fa7db7d4c9b8b8f41e985ceddc9c0eae5fa6731ec10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a5091ee72491c3f7db888ab666543e301faaf8faa2a68195ae4f87c0e42902510de79f8262f47685355990b5eab4e4a848cc5dc186215e76cdd6e768a7eef1505f5817860b18b26a1cdf44e3b4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18801505330f11246727ca487adffe728c09add3fddbb906bb00332cc9ae4b00470a90445cb6e063ae23de78b7643885912c76d74c412744d2610200714c9c59b8ccc4e5c2e66f3c69e71582d2eaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20120b7fc7e5d7cc70ccd1dc6f8c158500c50d329a25c87639dce0907972d8cad4b47d41412e25253ae928fb6186684b63cdd2948f8b62fb3a0c946e3fb73dd811d320230fdb3f4d60956d424c91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28cf22b249ac60860c2ce997eb54ff7ad2d27bd9108cf8e2988671208d34782feb170393aec436625acb5da215bfc1c760f24721321073bae1493621217436833e09840d11c099c4c437e7752aec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9d89d7c6e5400f345f39702eb5421246b0d4bded6e96d1be6890117a4cbdbb734063a235155ca84bcfd8bfd0a786f496b51afca63254ebe88ad63395272b2555cd355e98c6eea90826a6f7016e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6c48075bfa5953a3a470b9f53786ece66de1f7675afd3e538b46ffa36c904596969d52658b1ec74427a286e12ba1a5d7c2e0ac7924ad342e928d6fe53b8335286000b329a00c3fad3cc86dd978a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7aca03648405177c50f8a81af24dcbb11ba727ff13f39098904bf2e0808811f1d40ea3b3cdebc210492187016e6c85c764343d2e09efd8171dc0c4ed37005cc5bb18afc806292e559f7d944c792d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b56d38d94ca364f996152c65a80df8f62b3347ff27d3420eebe16403c27a61290a11d101556b7c0f752ef64844e89fcf702c7a11e31972042b1a5f3246aacdd886d9c62021e0251f3c450d570a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ddf4e0cd4f8ccd78cf99f8737bde37e1abec4bc3d34f37fed2b618310c7b8ca9ed36cac3b3acaf57274604987f68c8b53db7d5ea4cb24553cad743ec8fa96aa9993c541cbfd55517cd7970972ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173a2f469f571ee70f236caee1a1906ef1d95f05a472e1dc7fbe2bac9010fb95d3052def21fc8287c0f54e244cd28189e1cf88e159fe4a7da1587b56cffb6c0a28ea046deb7e766bee9861225b440;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13161245ad4c6f22762d5add590150f432877a684090953096e9610fb74495e7888610bb8d2f9a476a2171480f91b0452e1925dc4b811b680e6ba2af8b9862cc2157d795087f2ccbe78f4bc82d4ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haadcec1b83f7975882cba9fd734160a4cd36a595dad2034964c6a328880a9f26de3f8a83206353a020099008555c8ae0459942eb33114059f98a286ee438ee34419f02ef87ac151d385b332dad20;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123066f2af3d09a9b4bea0c95fe7d200b3950bcf209b6f1e2aeb70e7b2b348fc445f2e5c4d0d69d3ca42ee9fa513cbaf1bffa60cf736d6dfd7477765cdb858da7439dd16683421a4c14d027878432;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4add29971bf8782adffabb7cf3867320750d361eeffc7ff373ae42608d5391e34a2e995c058c9a49cd65c5d244641b4af9a24380d6e4c6b2d91482dd19bcd474c8a232eb0b108e110dd8d58d17cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1145a77234a41a3fb06225b5074af0712a85195714fef95669ed65bb899f117faf5b538774e9f8825a5958e403b67a2bba9679cc11e0c958dcd6d51f8b013c5c711154300a95ce0e5dbc09d39da13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1756a4f1bc70d4b8d3c0bae9c34c23c54ecb5f0afe38d8d1f5136878c05e1e5fa8c90ec2ed3ef050eaa918ee18c06c48c944cf9094ae94018c1e9e73c87b6776002d0f9d6ed5398af616aad9022c0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10aebded526404eb994c996336667c6a37540813bcd5677b309406e1d12c37d793b154b932aa8b4f85ef9decae801db1e18f275335d16af42824bc0bfa95c250764312c4a24d8b1ecca792110f8ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8ae5ed09df41e87bb7c2c8fae2ef4da0b524387f2e3d67fc0a517ee9de36943de0099c80ebed39f339ab0be210902aafb13fde74831efea42f00f51a8983cff63ff9e22ea9e2eda2d57306ba2a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab1cf28eb0250771edffa82e122f382665c26dad15c2be829edbc91c99b6b704ad3e4e252adcb501b2346c8c2d904a7f8fffaa79b6e4a462556c70c79bc6f74d3eb82a334f0f186b127cadc97fb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11068732c4aef99c6b0123ac3e8861b94ae438e73320a8817410acf9866081d1c2f3b68391fe3a5b087aec0cd64ffa79eb4abba3da939af39413b5658242a8a315abf781579550ac9f1c0e2b013fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h734b2b2279500695da40655b38797c009a4fe47b4b3d46693dddd32b29a616fcfcc6579e015112d7dc06db1a930c89c55ce74ce65138c9908876e9055d023aaa3a81bcadd99ad683d3858e97d9a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h453447d84b51b303460f6a9cbab245d37af86fb8c2f8f4d20f9c0861e512107520aa5c09fc215bfd57131b021009e8d67654bffd30872e56ee5abb6a123eab76905c0012fc8c031b2db031681bf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ce82a3286253ea1958016b1df3ec78dd280df45c65894893523b97ddf5c7b1687ef5a39fd092b7ede3516005577b7c90e72ed316e5734e961945ad01dad9288005592cb23d14910338b907b6faa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5088371ce298be79bd33adf5d735d9dfaafd9a9a0883836d13ee89f13b9af6fe9741ca7da01246b7982ec08d1c9e37961fa5a0fe6c22aef7f413bed5d43147fb495f78e59b69abb25bfac452ac14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5cd7936117da26e6ae1dc5dade23671ad164172c13a4ffe1ef00ddfe286b8fffe84c1c41fc9029432a06e6e4a30d39759a8d85551c9d6a24fe01d9fbc013b923427c07542a9a37d8c752b3f7fe49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f31937e39c391eabccaa73d4743f94cc98175d64213df4933d97f3c05064ca6babcd5c0d2b98d142aef34b4fae33ab55b7d8aab73ee1a87047612865bbe6636c8f2d6114f04217ddcc5a928f30c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c226c7151aeafd6047fd7900478a5ab913dd9906313a89be128772767c9c861792da5fb317ba70d8961463e6b78b6382775883c926de9e967ae8c2e3def44c940f001017d6c446e86fad0bb9bee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf713402060665ae8d65fb0cfe40902220256ae75655885e5762ba12dcb0b7c0302a592efb90c48cdbdb5d0a43d37ec55284dba366b1763ccf98cd17b411c9af3b80e141f721ce07054b39ae34c77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c4c802efa1424c44523573f9d317f4d5801526c6d28f5392fbf5a6b63cd609f3ec887a58c96eb73d0b1831097079056f0bd3a123c4c00332ee09eea271b8e74a6378cfd9a054215a62ba8a9698b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6721c5c71c1278310bb8d609675f1817b5b5d21d84a8df70818b9a0010a0db6aa346d96190d6746a433eba03381c0b746ad4d2ae7d88bd6b81ebe0d1a6fa160846030b03730f70d9e83d2221ccd9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9bc6fa205558e8ab9b9794b3031a143a23945e349f353cf48d2de8f2968eb79d2127fbff6fe95f3c46f35fcdb81ae43c55b92e53ddeee687a085196472fb5c45d5c6f15e9faebacba625f54012e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e5f8cc97443867226c55081ed9e2b5a269299a9918df30b13462cc1e9b86c33c43f6aae2fd1e7f12baf597613091d8824236957e13509567ee60f9f3dabea3aed7966ad8505138cfcd6ef6cf2c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57c769c36128ab3d49fbd16cb6a4ed96bff4b6531bef5308b96e545759a66d1946ea51385bc2b2ad65e6180f94fbb554d6ed454f1d68cf9137eec1e1f5b2e5dda8a14e21886d4b66993846241053;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f1ade0f338b234f771337f2db41e5a443755bdcbee9d5e1dd75fd7bdfe0569d285a27d9626ea04ce192390189ac5c1208bd65d89385935ae866c3ded3ae3bb4546b69e29f4e1ceb1823a2e8c8df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196cc23bd6ffa74cb525ff2b8dd8dd80e9c1fd3806178204dbe96d0e64f241f3a64224a75321b4883edca158f765e4c19562c5dd254e6394a37ed279d4a151b95366000897d7d27485c569929827e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e80fdc1c12f7c00accd1f64892821614cfe808bb3798d1ab94a3765bf4d44ff39aabcd95e6540651a2e6e17fef6e09108d679ce5e75731cf346d0caf09c3a335ced93e8e80b2ebabf20b63fe6ea8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c610f8e8ab25dc7b334457a6f1f447ce4133d95504e99fd0e5252dea2d092dd9c35a713fa68d3fc186dd0598fc9c5d4d7476c39ecebf0ad1c87f67be7c2bfe80f91d6867ab48fd81e88c293db780;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164ff67aefa76476ee7303319b4d99571e3f0b067453b5ccd5f9594c9f26986f868c9ba985d6b37d91c324d9bca3a3bf6604e1d078f1b4804bd215d498b820e941dd230e274c9d8e1b4a80cbd5bbc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2eb8014588e26888cb827a51e3c8bdfa69a5450ef618f248d1703e0c0d6fb2f6e56a194f09ae415f78cab1991b5470dbcca857712424f861be8b55593aeb9e8c78a626c60bf02b2c84f94274c19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132fbffbbb6c525849a372bbb8a833b3800e4db5cc974a414d4af16169f51b56f356685aca412bed29a47882be3da8337d14e6fe4c386cb9efc1bc9eeb4a241afca430007c0b55e72b6e27760ae4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe7df64001e299edb1a11395fc302adeeb17e7d26c9f72be0b0d828535e751f7ec00ffcaae4d0b1a544cc58ed814467103c2a0156b239ea8f6596ef7cc280a9266b66f1f366a8900b22084705b61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18293ca1b3538fa6eb603539addef9415662fceb9504dcbc543d6b82148ad6f21a046c9f4109ab48aae56a3a3a58acaa5c44e3665763ca43a695e9179bbbe0973b7f8a2c2679a6b4b965fb604b462;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f58ea90b6d4e51d0d74c746955851200f6f368dea4d9c725f71c19ddb9d71883d8bae5859d934dbf461a42be167212edd8efa9a01c3d608a9e6a522270233b5f05d2b4a6e564fce73524cdbfb58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d5a72aa7df6ea4674fb96e633a361c39a4495263127dc24176c6c73a76d1b09f6dbc8e23d9359622822bb20d2f72a314be72244ed140331f8995198da42a87ca654975db3dc07a4726d4d952875;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h266e8ffb294acd6ca0bfc115eaf07cc0df4a19d9fff5fb553a7a714404166e7f4627a14b477608febee67d3813dea94d0e4c1d07a6a9ed508a6cab77dc2192ee94adce9602052a60bb63bcd034fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb17133d2bdb6a82fb0629aac9d88e7e0583a2d7b05c46b8f9f7d725fd05593fcafb163923c89f39f64e5fa229fe353aaa6a69dcd70dc0a3291e6640ad585fd77e0848f20df62e15d5912be65b28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49f6010c09971e5bd95c2121a206ac19a987fc06faebb9e381d5721514a8a7917151b0463704e0fc7c81889e06cf9ec0b6fbf247ffd75d6b11725db8dff28cc328cd03cb74d8641741de7f7f5c6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185266bd0e3525f547dd0a5348d9ff57568912c5c2b5e9a0af86793ce3d72ad8835fa54d8184be6e73ce9fe7a368d554993339cbf7aec8acf744b2a3a13fd0b67f45a5ebaaa52abf1f0132f36de11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h373c25a2480917d19f64b5bacfd953ae751b7495a292860a4c146c70ead47c7b6f5f09ec79104aa9d00555ee4123d63f450cbc64f817ccc80dcc2087441c1abe1a75f640dd5d281955aea71e0254;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25d235b9f0e47655891e2df644cb6920c229531340ef52f89fd3a5afc280dfaf3cc7db151cac7b928f67393b0e71ca0570dbf2464a7b7cb3f41ec6a1667e53b1333293dab30b7150293b2f8a0d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e59337bb44f7d6349e30002c35f66afea1f1031d263f9d24cd819eb8b5f79fad4b901c4d4d4511d2154f302b8eb796f9604fc6a25a9accc27efec52f3cb5f90dabda2ac640195e7d1fe8f1f3d69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1540d4370768467d410001789bc7cf8912c736e9b3859204383ce21ecce92afc322a7157977cc05c625a7c1e7227985b2b355ca0c7353ae7adc8ef2d3db729ee63b56c6581892b70fc766708df06a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183f80f9816e0898dc567d572b4824e910fd3aafcc5aed4e108cff67a02cdba6b6d95bb9a787eaffdd7f2d4fbef44e98a93aa6c9a57b2587822f31d31a0cf00709e0ccfbb7b5ad005956d08cb7af2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4c7f0ded9d90748999c722a7b354264a554ea6b11f5bdb5d65883484467dac88eb843db50b124dc48848da0ddc3f2d22ad52d78c88cb3391b8564660a215ca9032a200b4885f90fbd1c45fadd58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175350a1a456ebffee4aca120022b0e638093a5aa252ebb8a9bf405377dc34292f05cd145d1fda981b4d4761a3b258401b6e251e098f7db2eed073cabb5e4b844ceb0ea05cf24ddb3fee9a82af2e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67f4d7fdc6872126bce212f55ce97064e8a02222d4cfe33375af393f7551e38012d59bce82c6d91e522794ae7741c17e46fd61f5dc8f40da5f3bf6088c98972fdca6584b17bb64a61be73bf1652f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a2fdf3a9d535a185afcb5e9f98086720dae63801c74ee11073fcff2de723689003e70fdb8e4744a79690659044075fab488dd04f59fb1d3ff322c0d52feddbc83e1e59f1c7c6bd159def02f84ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138cb0daaa10a7c91843faa891d0933c13ddb56c394b5769d6700cf8a3d881b30a2d654aacf0bded9cc05fd90ad8c69798d48965237b691116ffa5b79dc7e8f1a14463387a20f6bb2090e39a57fd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194f731a015cfba9d89308f12eb8f21ba1e7f516bf838e220ae1c832b2ec3ecce5d364138d8804a3c47623d9c1419abc1c42502febdfb438e9995751283a6298b0828770e1542eeae12cb12f613ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab4c7c8202c1588e97398f598970288cb54439a35cede46d43b2f8360b14b6821e3429859bb928e8741efefe5d1fcee1a18f134bb664285f8e8dc7a595f8c049815ed7f479733d56250137190c75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185dd9e47d8f56e39c643ac74a3b906d581e76ba6a2490679cd8cdb0c23c90a3d37cb1c834d0226d0a17ee711b7e30f7757ce4dc7bcd8e68ed9c37460e288ddec5d00701ce3527a0aaeb10abf01e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64d58f116ac8a4f37091acddeb5d2a7cc496b80fae74e8d648289cdfb6d79709bd44b0b77b43e881b2382aa002f8af14355355345aa414ba45590fab4ad0c2290b12b941fde010bd28f3557c8a0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef15b6538c305c4c966479770e94cb901c49773a6dfeeb12803c64c00fae2d5c71a3db6d0c22b638776fbb565293558ae95cdb5803978221c998cefd3c9a6fbccaf1b2adfd6d0652117460a63e9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15df86206f1a23d12e16bed0419fa0d08a6d1d0d9ee92838e2139e0a4a14228c860d9cd976692478173a3191c88c8983847658ff3a9473e23ffc4c095040a9938da9db66100262b2836f531ee4fd2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7141c6f725e2e1149165aff6d2ec4d981fd94cc3bfaf670ba8ecdaa0ad73e7c632b731715cfe2fb6006d99007e90bd4499b49f9680d35bb952164282999e411956077ad6ff88d03ec9c65ba5732;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b569ef08812681dd223071c0fe4e0b83113b575efd534a243c1a79f7b4e15e9583a027bdd778f7cb996c423a1298dee91a7862592228824662ce32778082381fa953f3be9b1c661991a14e253b44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132e091faf978fec8547b615fcff2caba4c223f0229fcc8fa2fa1a4d5ace2a232073e29293f5b27b3e15d7b5752df00120b6a587c4d6fb84f45418b401a4cf114d272c6580d2ada7928f0d7894c13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11318892a3284f5e44d2e4fe8b2c34c12f95c366bf003dc38f6e92bc1467c00f4ba85e597142e3b925be9022ec51a9e9e71a2897d61ad2df5e4bdfd9b8b62748c33eed99550a31c2c14ba45d22155;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f708484958d56d77ba558bffcf53338096e856bff742dbb825386adcb4ea42f7397ed11c7cf8b6ddab7f9df00e6db3c341ada7c3d13c707d106ff791df164605a5ebdd54f8719c9f1f9a46e03c21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd81a2b1f15262f2e88e8a55cd15ec28fbe8cfbd863bbea00845687fde68c7674a505bd18bd3b9c5cc78e7fc88901682bead13852f168b97ebd6ebffb6c5db7996cfd08c3e22f29b8975e3ad38dab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce8864fc71dd1180e533c7b55dfa551168bedd30628b62b36e34c3ec33ab3f622abe185a66a7977aa5d7cb5a465bf58b617e1572e77727b94c28659b573e59dc724d3be1e8f9bef3a300c6fef0d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee53ffc877f384a765824cf13efbc5cd130084d25b70113a60eb05a8c3d50a85301e62f46bd6d3ea4d26f9e780f21d769838f38f53c3f01b4ab72d50d92a6be6e1876167303253ee792650a8abbc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habe2abe219fc3ae77ca151c319be65f8464aee0c4103009ea183b49331e6d90329906a58dacb5829c200194b5b18d87c1c3754e47386b133e0cfe7b94395bb2c8ccbcfe02926d105e4f8c59d9378;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d8c36d1334e072665c01a97a69ef4b31eebfa53ad038111ff24cfa72d489a77d7cf5398fad2d41dc932f81716790bb1215b3590c38899081170c64c22369f0ee251e4efddd941b7d09186c7d5c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69caeccf06940b5e805e191cabe14d2ee1747b5eeb4a5ab29a780e2d18359b36a48a4b444fb05a3a1afdeb5a36a5effaaaa19746c162c497a9b09857a4a13da8f84d55ec889e27ffe7c1b1159aa1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79d3d5e8c2df64a5d852ea2ae05ac07623055c3e35b8e1d039e21d10aafcdc93e0d263f8ae5c3dbc2d0a3d3ee12567cade438ec45e645106864190bc3819cce7929ec4db71cc5eee7c55dfec6716;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f04a07ea7720e6eee4962b7066676593b25b89d3fc36ee2d0307aa2fc3a9cd803837295325a71d334574634408983c2adb81d7cf1cf62f12162aab8199e403ed4123f2e4e6ac42e887a4205a07da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd1bb04508a727046bb1544ecdeba4c7a3cf5d68a58a7ab186b7bd040d588c0a62b2ec255d4b6258f960df46b32ac624e88146ff82f9692c5cbfcc43e19cd565e59356570e9ae738c18a51aa4ead;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0abded0c645e22de353d3f84a413532cfa78d4186fb5beccc214869b333789a8f89d0f70404ec695bfadef2f420c094eba9a2ed3a6bba8020d51158aab3210aa2611b47c138f3345d9d5500f26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8425c3a5554f974687bc90035d5c744a048f4f7c56b139c2619832596c43baa0f8405d40932c6ef2d44bc73fa5b91c9a8bbe6778310eae08298837ca90c072e7f74da08f23ceb402f9e695219e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7ef075a92af36b730a172a1024adaf2adc28e9a5d01780fab1fe3e51daca8355730d97026ceecb511339c5594e3e600f2e830f325bd7c0f7d08fd4b6b550a37a5343407575407e6f134be2e9cbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c9ea4f633d65f10f8d7d30bf10ba6c37185dd1572f022d8924d4dfc12746ee2313cb9f92b196854c03bbcc915c89c904126b82df165238ed2655e0bf795e2b0daefc1f7e41fb4073f9e484c8621;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae02cc6f4f8fd489eea8aaa9d41179d7c87009b04a5eba8643cce613fbd396f934df7fc85ee684a9fd3983d3dd110baff1500ccc02155c97882571929c2acd0a059c80a6332f42a9fd13a8fd1b8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b534668300e82bcb3f2bb5aa5260449e6c1538227af17094260491b1bfe1409510b00c04d2c8a7051723530359a07ece083e8ac4745fd1b856cd3d37880bb84fdb9e63f22368448cbda9486da6b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69a448f5af8f0d606e84f13d4c7db8d1f9a36d9069a7ac9e62691820fde0bc10af5f452864efa7906dd3e7125939b2a1aa2555ec5ecc658c5aa47462bffab2a240b5ab979f11900ee658d376434;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd06f17fe544b1092915bf4fbdfe89ff1e42d6e07bf6f27700d312d28056b994659c0315920fea3898db54bd4b155b32d9109f0eb11b97e8ab99b4b42b8178bdc7fc00b7f1d27553a6c0dc28d987;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18439cd40d62036b6f509058b825ec6933575e39937af219ddd3029799b317232ed0acfce82ed4bfa5084e5d65380fb35954d91dbbd62073c71e3065df282ea325f7082d73a2d19f5494a012ac0a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7870a472538acfa5336a8587d88db15ab1a10f18a344ebda6071e4c200f134c1a79929144c5e29dd8d6facb97a5b1bf7c398629dc5aea299dbd22f2d064c0621daa956d3a92ba46ca7692a769fd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158702b5ee9c2977d20f74b009677309cb0b2120aa621f580a92210c24b1a5910a2c2711b42de4b46740f3f7a0c54f05c9ad1c2108d0407087101048e602d3da6d82a0e86384d9aa7a78dc7ec67fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111d6a8a399ece5ad13cf90f507eed26fab291351fab62eb897486fb8744a317824add4269bdbbd625366154c4556442e9da64eca4b96fa830757717bd7813b1e0c50064ed535bd9032b956e245c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h881e3971c433feb847a398fef70066dca7d261cf720528391f6f7523a9d2e450d008b0bdc8936c57413abd008897d59637b2db8457ed04725d75ecd6fb77f81fce3fdd5b6e5ac74b01a5d58e2565;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc7de59c002dc86c4e3492b7d49e900e20356dfd9c413245bfe26a237e3f55d3fc144250a6ab014091cee7dd09cc91c1da11513d48a5899c7b37ba0f7a0dcc0a20684e60f5497e51334861aa2f07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d192a7885b9fad3d9342024ad1809c119da0d1813db5c1defbbd4359418ac3c904bebbd297bd07086d3c802d2da20b2e8257e37d45f5b3fcf6ac35d65df73a96b0abbdb50badb78cf8c261951565;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c45bce22d77cd5ca1f0f9d2cce9f1762045add57940638e6fc5a946a23e6fe74ae575eaf024ada1264627de95cbbcbfc03f05ccfbcdf825168faddb9195b3d6be9e29503932b41d7c88a5f607ab3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d43290fd91d328e70f2521f1e9cb4c17677a7c64a7d7cbabb644e5ece4caf8db80a98c49898b105ef8e87ef4d9d2237b8665ba024ee1f95bfadd344d1843294b0dc215ae393fa8fbbef7151cd8d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e6ba2e61075660f548b6fc0f84093ab83052b3355bf62066c6cf9014271980c49a748bbf844b3952cc3e7c860a3e886e19bab83a8552dd2700bb880976739bb9f41146d8957d2bf14d304f59e5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7526ba792ec844899e5201ae7592a1b04d7c283d1d2ae90147b94ffc9daf2280cb096997328b5e69953b357fa8cd7d9e8100b6d36de8032468f69c0c3bac650dcce4070dc6a0fa5e41543cdf091f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b150c8869373e5591e4e1d201514bdb9ff05c4292e3d12a1d9154e8e690d575b8cd3507537f25112260c6059d4062be429018d0652ab9fad3c952f71a66a138a8660b24907848ea1ad7b3e93a732;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163f203dcbc257a75b9fe5bd77eb850245a9a314e597c187d268380ddc3ad8470754186afa4115db45d41a2c94755102c14590f519803804966d6040c9e1b3a70e86d7341bd31257b59685706482b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44ad3bc24ac99d506eb399aad82178ca26b8cb06c13c3ac9522162f814cca0b9c974e5af6543c3ac4b4add0572786897ee39d93d9bab67b3d4dc54659ceff617d208321023c4d4a8ff8f26fb01b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b96683eae8445556e1dd4e5dbb39d1770c221e69697e31b1ec77a6e61a7c38e97da2f795e6a88ec91d3dd988b0fdbb4154333ab2ca4fad5efedb45c0e8f0821500a6cb3630dc7f0caaf6ce731e07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4471e576e3b5b425488b17a3035dc6e553a07617ea0b0f9a4fb18f3a82f765b7d49b68d192881f99a9c06dfd9ffbdecfa5545ae1742049911c5f61653843a9646bec92da8c1ac3dc5b5bdc36e00e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8fc7c9c92484229200211b269296bf6a80c396323a851d6f5220f7a164e7d804b1efdb0b15218ed34c47b9365087bb18accc3587d96b52cf56fd48f1bd239216d45853cfda75fbbc83b23a8aabe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8aebac72c7f5419265a9d4ddd20228a60eef4a6fc92e9a43920735f0c0fb09b5007ea103885816bdabe69ba428d522d8bd01b5a9dc68995e4fd2b2ff031f1dfa5a5d515958bc588c8b519657ada;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heaf6d5c1285e7862536178a1f22b34025ad75a96786a315ff89e3b044f8cad8345d48e4f75c0d6fa66ccb96e71ccf76b14b228a9758f7c3da4ea145ec6e3a3a4d1964a43a7d51140874b9a20f396;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b18b32350cb4999927d249f92d1e064011d721acad584e7930548a3eaebae7a66c3b1481e482cca9fd6bf433704290a79570a66a2707d965eba747d2cc277711b7deb0367892c7193f323cd12ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185c03abcd55ef9cbfdabf6099b088eaca967e51e71e908e67b990469f5e0f1d7573732f488276e2bf415d681f3499af31c45bcf99dfd04e989e5b57cbf545223de4c1e8f2bd0fca2916db15f6d08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdf01b7e1813a0b8b67c33e49cdea13eba3ded082762583aafa8137f0ed4f48b643fe069d0117114faa054c326c0bae71a6ce9e7e75fd89d89771e2722b944e82c1f91f4bee104f04a2f8585b9d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee884cf3243bfade71e04c3cd0dad86d9ba14ee447c78deb443be77228e4f83c61c0dc16f83feb29b8133f317c6879861833da53d94bb353d79b874b916b7c88d5c240a885497993d707c6c55211;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33038f008b5bbb7b73b15a990dc62decd599657f57b3e1cf4cbe208713b4c2c697b6828ee95acf5a803bc21705603096a932f6a295115b0567ab5b70f358cd991686b5c439fd7fde477718671f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34a4cd56b0c03bd939be958e43960e61dd6de3e6597eb6aa32f15d96a1d67235dd9495c4f3ea04cf29932f7cf921e423759faf4cad0e974089d8ab18ac3de401533deb7c2d2f8ce65e72d9696ca7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a5ae524a4cb889ae5ebee206159aaab790ed5c610e6f7edf42c47bf606f516368605171c2317060a840e2af048caee8b420213d499dd92b7063721c47158ea351379b2862a8e496c5cce1b8ff2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8d624ff05e8b01f3065565c72e8811265b1a6a8755ed338fd6e46f7197bf10832348d48cdb37430103f96c5d9f82c112ed50c8d270e23ff84481754ecc60a44580c607f5429fe4d91d60d1425ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4f88f278bc391ba6714436a7fae90b008f1a55ffe2c3e780e272dc3f6e0bf3d4bee6f7d7d8b578b3a05ebb9114dd931ebbdd3e942ee3c176c46036e4c6090ef29fd471447315b217aa1a22a647;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137182fb8546fc68e4ef4203b882acd5083f9970541df2074c91d9d785b3d0523eccb1b69957a35b3aa4f915ac3ad039a7ff14d7c629c3b5d6a760fc4e24dfa99c08128e9147d078f03088e24fc5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c139a26e1492d316aaa039d38b4e1f4909839e4cc72890ff15372cfe824bbabdb523f3019617503d52a82911bdd732138493c0de1cf1020a2dbcb1444357c444e9587cacf974668989c653080ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb898ddf2db148a8bd8e11d686cff26cfe2e2059bf8b6b8ba48fdabffb3e883646da000b17edfcdd1cce35dbd73892f380a68d9e3bb29e9f6b12990f166d4ace6333adc38dbf9a5fa9123ca0026c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b889f4373857e9986335ac52dfafdc2241b3a3fd963a1a492a3ef789c0c9ef74204fe385049592894f66870cc8a0908197b82f5d60385f00dc4118ffa9327e0e0b32ed764df990dfcdf418f441e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heda136f9fa44938ebb4ab8d5f546cd25b7a458aa4f7ef5a44bb4840fd592741bc2cf491438c56ed32b256a0b5dd7c0dabc964998b33c2cb0c0da7247b4bfbfd9310d7d192f70d9bb29b50d50188c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h917bfcf6effc2427245483f5f48f4204dc974b13a0da35d09ad1d976e65466055f97e3f7b3ae820b19584861174ae8b6faebe538b74f438e9ac644c24f4e5a8c7dd3fede74ff00fe3e5f6dc724df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ce23b3de278b7b95e93bfcc149cf189a045e0cb2f95a4e03e46faa7666addae40ed5015c0da4f16724c22e10b82d8a7b7a067185c927d51aa5c8c959745f7c1fa01409afef9e20211dcf0a4b3c0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6ce86ba30718d5c41475f6614fcff082fa9d531cb5499dbb60560a553d771d719b1283f62788a7c511d17360efe4f492e6a20a79d74560bb9e6b8901f32cacd43939e9ba4ac0f99d2ca4859155c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82acaf3be0dc513d39aeee826e76144fe3c98bb851089e2eefe53134a952abd22fedadae080715f870f56403b2998d5091b430aa4c591aa392d2e79743f328a6f39b66ffd0789fa53ca8118ee52f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfaf0c37b732b43cec7b7554701d1a51fd917c20b770107901e5aaaff6b6c1324c92ddb38e9e5071393368231111908a779e38e5bbce1c7d94c2e88cbd2e7672e4b97553417d527a079606bdb873;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109e92f5b2f6b53bf1e47422bd22bcbc3630784f4d3727a7d1bb1f15bb6b51c713d714463decde8a21c5054a45e9036e83a505bbc6fcab4e7577a4a1ffcf8dc9072b146924248946868105506a490;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175a269ab4f0b341d57a316a1c59d61c4a0f664292dbdde79c6105f06c4b2981a571eca06d8995c149881fa736cf7b19896e4b878c2e025bbdda3ab26bf86af722d0f3a8bc7517f695f054cddcba1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfda1498192a5d76a9b79241aca10edab64fc39bc31fce87227132707029b616b3960bc7468f047eccf69790c3ef3d5daa787c9eb69924b5b8c625b7a9d8f747701065cc26e9568dc7e6490dc0af9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef9a8f816c4605fcf84bbe397f01c24018f84a414eeed8bcb682b9db3502c0a80ba9b0f080eeb2646fe2340991bbb20b80adabb815852ee51a77df405d21fcf7d691bfbdb10a3fd9513acf027074;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf75018185dc62806835be95354153e6405aad0efb4f0731fe5c0913de558b6ed244f8b08f1f21ae65d3b5805238fe64efcd1e20e23c1e8d490e865b27f5ea1fa81797a98d73bad3c79a8f4231b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1907278bc0e7057a6ffdc8dd5e1dce3d63e4f2d6e84ff453e566401803761c71cb70201788f7a5dfe9555c81bbd3793316acf0609a3873a3098bc9aa2043cd5f175630241f7fe4cdf8d191ac3e849;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f55433733fdb42a2cd3ad52766501d776d26fac2e2545b5df5371621e060d05528609a2a204e35ecee2d0c77916c232dfb5cf5c378817849b66b83df618f32842c7c5ce663255f1c5253607af54;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db0cae885cfd1cf9892e5f919c14cc81525b7c2e6b7491055f72ee03683fa94125d3f920e9dd5b9f836d4e34192ec93751adfae8a7d4b4ee023fe46bfd6d3a9e579e2a30fea9b4593fa745f95eee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9b283f8f69720018d9a352bf3311f05e1a98b3d04d057ce942291bab2816bbc720a81c5ded3785e1c0d9a5c35c0337c4adaa56873ade59ec962837a40467b164e74d67cd44b56a242b5833eef93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbb8c13aeee4e13171fcad6ee49c3a5f6098ff9ef5754510c4ec67e1980d5760bb2fbf30fcdb052279ac8699c5a47179a483e9dcd301ef83dcc178e0c4bfbb5cd6af19b3bd0d06c144d1b04aa62f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6f3f7ca6d5131b1fae0622618d4e26060a9b334d74c3cd059ea5f93e05ea2266021ca8dc1ef489e6c61ca82349b8703f0de76eb4d793f30af5fce7502e7f8e42c81a8881a5c52254ef92907291f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c87f9291b7b77176ff43c20af60ebc498b05e9de757899d9dafaa04867ff744c691d43c53b3b3ea1150c01ec247d9f8459befdd0a3926050b19cc0e05cf0617b6f1a3e3d4f38ee2274eeb5ed8e28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171ab34b42818752053d908591e31bee2c043efdb1ced6a4a3279bfcb3f58dff4074d100fb964282e693b419d5041a3ffc09aa3aebb9c0d980021196df1fca3af53c4c0f6d417019cb2d4416f0cb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b4b2488c299a41c56e6187430870260348d9d0525c8731ebcfb2b78420b6ef9ac8af85401094a12808c0780c65d65e21a72a525761c219e21b56a816ace4d70b9047e0ecf3a03ff708363e70db4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3338f096cd9ebaa5e2e9a42ce0d3ced4c31ac7d377b306642e1318f2117f5df29bcad39936bd15cecfe8eef61f80990a513e9f382737dbbaee47093e7b625e9d6599510d4839590db6c2ef9a4904;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e4050039b36e9d6d38debfcbb93536a6e654edddab8c5379415eaadba2addd14fb8a3cdf8c65de581076db503bd405c1d7b6e52cfcb16ab7a0766a12c9052a5b7a6b6d4ce6a91ee50b88cc677d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44187d72206234e74111b747b0950baebf530ab8aa5a35c35f992b5481256ca7277010ac5b1ffa6b570bf699da56feea7c34b7c5eaef5609478414df109ec70ba1998517bcf89908dfb3a3f8f1c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf9555c9092bf5626d76ac1dd095229e228332ba152001c07ce4c76e1b538d1a83d25b6419a5553d4afd1764c8109d5085e061d6eb60cc70b97e784adcd789892b59aaf9c2130555bddcf3030777;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191ed436869e190ae043935e9653e076d8ab30389e3687aa92da4e1641100cbe2249370d8f68e0156b60d5b30ed98ad87c00dd5fcb38af122e5a406dd91f5edf84a8bd4e01eb0f6c6cc2595c70f97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b589c88b83cafb03c1279f87da961a84a1ae1eb0d1426f1edb53f34101197562bb9df7a42690a214a2a525f14c8a27bfe77141f898004cba1b8d94e1ec79356345a369e230adda232e58b69378b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7eeed0bb3638eebfdfad91a8e98f9cd7603aabf19efe8188f92ac48f653da361104f6b9e33668322af600641e7510c4f991cb91a8d93bdc872cee6adbe88fbf005366fd7cd451f67f5a785227f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a40f502f63f5015acee00239c44b925bca14618534163f980977a91fe934d67f7661d44f7b797ad1fa75bd5af4dc7302ed96773438a13f8fd91eda08f5c4206a590ea18ce5f4dc8b6f11cae6f806;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h293ab5dd5f0c51c6dbb3fca32aa321ce5c85632b64139a3e7d04f510310189f1ed1f152ef37645975de3d98ceee2906741d599811e961c2331f5a35774ccfd0544001e62356ee7d893c3853ce6bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b30f3e41515c9722c66dac531cb79f966a6d458af220c1bd816ed3d03be0133d8f0c77a7bcc43a6b5fa3a2a4f434c34c3fb73cd994ae7fd99acb7575c8c89bdf6155eb8a794158fcaedeeb3f454e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d2db1cd2da28d4bb16fef2e2aacb8e18c626e71bbd395ef51e68cdee1a5c2345d5c5a18d20c02e49491861ef4294aeb08eac91cc4d7b299a6bec6a93dbea8a26b15eb70edbb5e7210e9d5f80a50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc55814d4f51c0f8474d8f6bd2c37910fcde8e5a11f7798ac44537e826059458263e7c0a3df2570fff42347e9dba6e5255f0cdd64c9de04e1850e4f5022dbaeb7725d04497c7b88f658c893d0a1c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9118d8b16c4d3b551a07bc17935932637107682d25aded6d29b97a72bffb0b5f098423f11156692610c92aa515bcc6b7437a9ef93505318a7ccefcb9482ff757709629425cc7099a48b4a1f9a8e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fd3ba83531b907d833a85d8573382a742744c08cb5660903947aa4e026e8f780335fe389c9402b257639758f427bd65d595673b1e1c04ddd70f83e297c441d7ee72067fbe0e305ab857ee654505;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h531cfcc69f993fba02bd6e5b3f7a494213eda09e239205306902d29308b578a81e3300d94dfe8e5bc4f4315f87e86bae18f93d23c5e368ada7b8591c65e708b553d5726cd51f3b885acb8331b2c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haddfd1ba90c1f516f1b648a306f106709829327abedeb84f8724cca64c0fa21d002f4d1e11e39b96a14214b8ce4166e1cc9039d9b456fca2c3ef44eb5d0393df30c28cd8f68cee07c9d18c06f988;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf13a08fc10c245710fe9e9b69f69153e2db000fd208d93ce8d1258402c289a096a1bde150bd63bf51d0d602afb68e1286d73a210d24577f3eac4a2c12d3eeff42d79278698f892f8cd62631a368f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h667b10d006a5704cfa20c5bbd10464a3daa7ba7cf0f21ede72a9ff42b52a4decb8d785c15da3abf7a8cf28daa821904c8639d3cb6583348586d86ff63c01357c1385fb4bfb3c11f53e6e1749af32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc131639a93dc197def988a151311f1fa53a128e96cbe3baf3353dcca7e80bb73f01c71399fc8b90d2821c20cd3787f60d9efe3675d5821c12974dbaeca15ee8b52369c1285be92f33c3f6ccdecef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfad6f73486722abe9a4f50683a0f990026bc5f77e003fa966b78fa006fd12dedb30e038f615a259d72710466f31aac017bafe4c1a792a87775fb84c4353e2569f53552ea49273bb257b70f0f8b05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbf523d8d8f120f973a42c18ac27fa615ccea275d9c08cd566942a418dd10972ce63231135269ac1a2f7304f9a8621e5d04f23f70f5f5c7e974b635a79361fe6d9103e47813198a039b4be097a09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1add24de8bdc3b06635f7aa929c5b9edf9fdfd9418a4fe0aac97013410aa5f8a773e03466d648cfb45854c22deec7f3d54f141ccd0ff20f7028429ef3b0bbe9d0ff7620364e44bf629c674e8579e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1a07ad78212919d7879d6c418f01c8ff852fa8d36ecdb1be7e96650839f5ea44113aa9dedfef6075af58b4b818db039a533eac4267d714d6ebcf6cab07bc1ac78de4836ed13121d3c44dce8233;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4748ccc71edb26bcb47e3ebee8ceba2c3af2266b3b35725ca5a39be9f2ccaaf0c0ad36bd2e7c4d2b75df53e2b05e93e5f0f0a1ce1aad7f0f14949e1eb5e92731a47d6ff854b6051da1ef2744d32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afa18f2649ba68fefa35fd6dab4e4d43b0efc9664b0076ed93bf933574ac914e18d241af1af99abcda00b078997e2b360ada14fae04f5f23e06a0f9c53146357a2dd08bbb0159de8f7571152f28d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76f256b0b0cfa0037664808b8959572735a94dd5f3c0bb0dbfa729b67b374c9182ea86e2a87a0aaef28830220946e6f01570a24b868e3bb99be5524d55da338ca0639d246cd3ba5562ee490bb55b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6ded9eb19a57552408975d35082c8b9a62549041326f6a1e37e57c6c17954bf3e38a1d775897fa8439c9e54465a477aa98d3850711d9825ed526ab3336e8b3e07d4c7a088ca43788044b8cd5d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha375d62e8957b3e1d30e14ad3be46745801c4a39bc9c1f013f9e5f0209c2f3c54e2aac5c53cdc7f74bc70788c54c60afcea3ccaf7d1e5181ba76941bb1b40029fced71d5455a50d49c4c9017c4d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h585a40d897abab581203b230471261c9355ba5de52c98a448b4a0ac565bb371a4633046bce7af68ec38c0615634e29b19cf8c867abf68da7257d269781b86d37d2c05c811d76deb4b4be017322be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1293d32a9ecdd4eada5e0f7d1cdeb865e85eb989351763fa64071a9e528238b715b1e18502f89643e135df3328e34e54b2ccc85d63750412cbb1031873f1b54f4e42f8bee9fa04154632019553bf1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8195684ba2874b1b72ed866d49bf9e67ceb9a004839d553b548a000e3adc78c458c1dc0033f153300fce1a89342a5dbfacb39ddebe8723dfa768aebd229d2af1b3e45c6f4eebfaa97c4137208c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h476df222066ce4906d9a36f1484260267dbd614e8142dc1c1dbde53c4a5afe9404a8f0cb3788d7063a07a9f3e2f6df78c3cc2de511a2a0c1e2a871d0c687b7712b9e79ad5738f19b3b6ccec08d63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140f0d77b6023b15d52fec54ec162ac7bd6a214db9bc7a7591e1f9616c8fdca54f047dc620f9cb6c48ab1ed1197f168988d0d651f0caead822f6465b9a75ca64820bd06f1931636c75bc12685fbac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa6abf183d97b2e6f0e35c3aa9501a0857e68202af99c8e747071edc80540b1145cc16e7cffece853ea2368c9f9ba42ac263038a8f68d64a12395dd2840264841fd7ee665d72ee0169246a36a58e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32a3ae9c2dbe19046608b84ac43ec11a651c010ac6f5edb2404213034f24e6f67d56b8ed5ecddeffaf68aa3b7a15c487c86c7ce87113c7cdea2ffd99929bcf6da2a3cd3272e454b77dba922f924f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129baf2e806ad71745ed3f943ffa62f0ddae853701cdee89d45b95cbee2d847aa82b4bfba07f8aa8acba517b9069e407e7a0d7df9dbc6b2fb6e56f5c41ba34953da3475db166bad7180091b9aaf01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5144c020f3420ad8c85ddd8e8a1cb86427f6b63d5d600c70499d318a352d545104240cd054afbd25847a9c73c20e039aa470036596f57c4c45b6e372ae7cbfd6e05e5140112774613156f0f9d398;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a17f1e807b51d86a852c7d372b20146f7c7e007111be1a612580c41de7a4b8e1f53b5ba550dc10d87a45e954f3443ece653cf0b635d789491b264b841abb120974274bbf02b3b8e085da630693d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfff0886b562f91ac6906b4f05ae5a42df1dabf17632574bedf1d6c7068af1f8f9b64571363ad1e26ca5f5aa331f5b898a6545d005b3bfef6734febf96593abc9f9ecc0be46e848c26a7f63850db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182250ddada34acd4b6e0353c73f09a9c9ca67b3c72522d8d140f7ffe92d19fdeb18c1364c8a333f0525dfc089bce6a7585448b697098d9796a8e10f782f9cc4aa441324b68c5adc3baa40e0c6316;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfbb87e4e09ef66bf8b1021873bb028c6080832a9e9b070ee479de966e39190e42d7f18f194d8d2f730d3a85154a13bd3f4c1e074201fb3674c6609dd9973d57b887c007e6af3abddb6d2b54c388;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12241d7455301ea320738e1def7e075ac6669a22740f8c30e5ed983ad3485ddfce0d883bdb6577d4f091d054c51d344110be754da3bf6e3eddd12c875608179e26dcf6377eed90b970058849b82cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32556a0727c63757f065c8db2d8ca8c4ab77051fbc6f799f84ca9ae9d3521f6c5511fb10d36f88c4782b91f60d26f36d647fc57f53be407ef37c96cb713707964f97a55fd916e3b6323feebb2b69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f1480ca6d91f047dcdd0e493b836db261e2a60d35317e49d7adfddc9723dbb54769eb164dde9ab61e0c0ca32c52a29bb78a43cfeb4b214fa3777d8b9fb6859233800e8b71c0ddea8c7e3cc4cd52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b43934bc724a95fbe8e2b4e01799951f5b929a88e52a06b92dd2735155720036ea7a9321eb5569e148e1659346b1b2fc42ece44f2eadeb8a4618e75afe687cde5db318ee1be0624002235f833d96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86dee4487fb78d4863a7e1801af5bf883c3b6dcf09184b61c686e164b0b0779e8b23dc4959babf67b5df61d0b454c7408954631b718744a5bbd42932e919ed1a59caa05fa3a685d6b6f67e8d8477;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1958b88512379cf7458407252c37ff05da9fc02efa0f94da598ee2adae61e8299078e5752c1484fb479a8c18c7cddfab91f50bc7cd2cfe0541559d0bfa798c5d6dfd1241212f1ee2e8ee18d4f96ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee6518fda23e078c18503310a57967bdd1bd9556b59a0534498ba8f64656642c98529eaaaaea412b3e1482ce102db5d3f2d8b50ca75a6299dac5f0f0857616dd3896dce10365bee941552f1c9840;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f05b89cd5309790af7eabc62b8d3fafa912b2c2cf5a27c3ce5c3637d0ca472780911acdbf97111fef886513b6451b7ab504336405598d40738c07a1288d0d07ef6c3d0a1b51d38a4a4589f6d9a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1299f27b3d9bf9faa9a7a3374883621f25ba93d26e224bc0eae4998784a2af82ad30cc0b1a4bce878631b579e81667ba083ecb4eefbaeb69cb317ff9b900b431c2769db5cba4022399fcab790ef32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b2054bc315151cd6a70b62d1478524f636d137044a316fbbd617a73c83420d3c0b43dbe4dd22a5d05b0a04abf5baa4d29c6cb41f4bf8bf1c979e00fe15d17e61024c8f4faf4ac15800cac8fd5175;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9329dc87e77950a9f45fb21f5d323a698a5edadf569716f647041e4e49e825e1fadd036574f28fbdbd64c50ebd97f13f4aee6b6212860f22c1893b4dbeb70f53f4c7cb03d0ae0ab0027eaf3d76d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ffe856c209ebdceedbfa7a60f7aaa49b0853ee18eda5b6bd59daa270d66fbc45b9ca846dae88c29828b9fb46d0e7626480b373ebd189c5acf8978c8d97e483b7c94b8a0f3cb9dcb450af0d8d208;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82f80ec0a38c013e71bfb38e93dae96a91b9b27fc139898adbe1d9e6d141795b0e5a8f7e7430081e5ad69c227635724523256a2f8feedf9f2ab008d7788d771d1e58dda42d541433e489c3d24ae2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195fcb8ec440e027bff6e6d59ac033a94dc7cae5e5d718900126c479abbf87c0924f8b16956012d7b21bc34ab2f1d6c80e1effd29101300c0452a233bc40d5c161f5447aa1ef461740088462bcc1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a39434bf50192618dada52d45537d0f38baf3ffaca05767c0a00d9cb1a391735eaf38c17845c336d7e8c777b413b49434b2793a044b70c08d8786df7856988b0c08b36a7ab800edfb003d3fbce3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3926881c898fb2542a8c8e7f996be72dd8b89d7b355f6ead72305e6b481d2972699b497135b5b3683bd7e397ecaac93a2a6e135dbd67185c9f65b4f7723a1acb5937611275e8ac4bc2959ae08ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1daaa950ca4a07a8d47d65dbcfc65c04d7c839ef7cc6f712c4ed8fafdb8d3abb2d6088d93fbceb8a742476629a697dded0943fe18b96230af99e9c80adc37f347f69559b82b15627d28b125792cf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d41a7d5e8f118a8750762b225032598a8df4acb3c1d5b4228120ba5697352c1112c61f20abcaac27cb762f3cd3aa32723c28ea3397d3c4015db4dbe693d4d4cdf350cdb9db5c7eba6986d58cf338;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196a86fa5de7d59cf96c0b20495ebca478fcf976742822011b5ece45238ee5a410302734a015e9f7bbccea9091f1b6528239171186f9e7de6d8b4112bf6f2f36e7c978b5f45769239f5c2c66bab7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6be3c304ee705e72d711f1288454add7dd0f757ae2a93d2b5fe974dd2f8a6a8fe97c2f88455b33535b02afd51894afb325f1bce78bd4ecf82d6be27a4675095469d2385dfead12b7d203bc90503;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e335110b56a09514a9fd95c08b69e56c0297737a44d04fbb2a6c5a4a56c5f0da18e247014e1e960192b75b1c421ede9e9cdf33b6d57f842c12aca910d32530c4799e30b0127e8fb3cc2454252d57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca332874e8a85d8dd2633f2c788828cc96699bfc245203745f5f8b821ae6fe8240bd1ebe103f9f1e9c64b8488545a0db86e179c2cd40588d4cb2e53a2aeadbfe4bbdb70a4864517bf8864e72db7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4af2e4305453e444d3e224fac2398e655ac7f867ff60b425b955aad687677aae50b802034bd8e0c3e4b57bef829e1dc617e9052b2bdf532e13d0d05ee6d2064d1de35b86a7bf0a6da9715adec04e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50620b5aa39e21ac6134aefd6d375999f54f452c8058f689f15bb9f7773c27c8b9d7656b7b155bbfef746fbf36b6b9d2da7bff5f55659e287caa6091ba0dcdb6402879900ebfe18aefb0f60f819d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de103a99088e3faa56f213e8a595521e3f08e5dd844eaedc1074778cc6783bd2ae2f87322c60b5e08c4e5f1a143b043d6579a1e659d61ca34096284d0a49cd5fbf817d2de43d067515141322be28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfeb604e85f84b3289520c029813f184c556b1e36ecad901fc616b3d04422bc4781e3207bf64b9b1611563b933f6ac8167045fa38b7d47a541bddfdee89a0ade7072735aacaf62baa9dea38cdcf69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1164a5d94fe1220885e54ced2c088aba05bdf8bd623f3f581246fc6e7961d70c5aa3aac9bd41afa2e5cdc2391a9da0638e924280379094664f15fb16a75cd202e697f873776397af5c1dea110a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf934306a876d1d13ad4af3d9fd1be26c00930cb74d0002e91a8151a35ce1af41c32de493bb1aba8a19e1b664fbbfec4b4b1fba4c8a594755ff508ae0a0073dd588f7a7d75d81719e46f391b1d931;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a6d0ef35e5b82b392d7e60e6a6e491deb4d2ac926a17d4324f464939663a2f0175b86adaba05ec6117a666c894b5a26474a2c6fc9e3d792a0e35d1365c48c671ee580fc5cebd966db49e4d06e3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1524bb51b3480c85b5fafef58d26828941c66c4a3276df1846dd2f580fecbdadede9eadd282fa0ee5a821eed28f3e07d6e61433dc0b0109d92ca21971760dcbe0785db96ec6d7cc63a74727905552;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0bb233dff1b7e40d30d96f453b2b4a7aa5d34f71c6067f3f187d5a1a0d44dd5c8885e0b43a06ecd046479cd4f2875fb376e3ae2cce28a883c19036ce485d1073786d555db085402a7c242cda3a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a77fa3c5d3d4a09dec76bd148f19e9ca238f47a7de51bff2a056c5a8d05d99be4165d7d8b97e1410124536e144e7e35032ee4d0f9d9a0a7851582eb54fa91939284633f2e680f46707a9769bb08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hecf1e8ad1bd114d6705a4014c0a68e4e887c43b0cc88441bca270686e4fd6fee617b6652650cf16b707175a30f1248134a857bae40d5a7908fd330a0317cf8f0c144716ac0e4c88b5708f39bd159;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144eb3e179a54a05da8da370b2b97e3d16b14a631b8fc1e21ffe66a858c9c20ffe312775923ba795d89cf6835f3ddf569e3ef35cfcaeb9148532b62e4ba13332e515c0f22bfca7ecd0595fb8097e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148565dcaf653b3da7c8af452ce89f6035b5e703b57705c6c175e615da3f006967082b3f192a7334ece68d3262417006f908f44c7df91f1ea2adb3e9322e3579d41b84e112d720598b280cc54fbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hccec35246e65cd79ec8c7925698e060bb7aef5e8e8a70b7497d355ad96d4541e86256ff482409e32ee55c0f17227bad3b54327d44af4f82b1139d7ac1be7c8b223c8874acc3dfee282d2ae5fba57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5d98ec7a3c5fd7aaf0045cde24e411010dcb0f80be09b092088b568c796c73a5e7acc299d0a0b039b54c8734d40394cf8775d2b2598f39b0bf9bc7efb003960c7dfecc510035d7a8df1753ae056;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ac969e828baed0738321b1d7d11832ebcf5831720f6695ea989fc156879d2258f2f589bb5a7ecbb948822c552ed378c75af96ae42a29f6ca2cf5eadea7e7a269a9c8d942593517ff2e56ef652ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b319e221f1c2328cd11d21d7ec4d72a88f6a66d3d680387b590f9222784af7caa9a90ed1e82d2b0b12c29790e7bd73a13e4decdf82b9ba0087581098e1c7603eb7b88a4cf791ee2a68a72d4b8f7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6df7835125c69978ad9948e7cbf4767481e2b8e18862e41c2e0c56d3f5d4d077330d1b8dd50400a5f613674720adefa2d9551a13e2181fb9c42d5b2e4af36e7e9a83128ebf5811a18880086badf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b31d46fcd2909f3c76d0ab449abb944b2283f4cb42d9b049a843f872fb39571a16be0a8e212e0c7fd7e871fc29469631ccc37d7552edce35021986707e7f8864c67e4df72cad7afb0f275943115b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5cc6e653aa0351ce1752f44f1819af5ae330e5711deb991aa3796d7467f16a3c3c4a663057e4d0d60b3a4e7cee75d7875376b2f42d59957ce1e99f108f95bc12fab0d0c808455d70efbe3590bcc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7742ced1016b2fde717e16e118055657daf0baa26ea6d1e4033ba371629dc07befd575087ff11fd0fdbf76147ab2fc58a5c5383cbc61064d2d868fc89849611205133ada4c4be01d4c7ff11fff1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec3de1334439006067702fb7301a248807f8d94dc546660dff5582f122a8b16e4a420d437e072a5e8fcd3ea3c164be240ca1d37cd3444cc8a80b08e4d7cd5920799e4c89871adad0245f62ce272b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d66beb22de128ad288a578a7c5e91fa8fbe0024dced829ef0f7be606fbeac133da46b753b54af51386cdbe9da89f5057264787a643848d0b3e1559c02830baeed52f33c82000b2dbd3e192bcec11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3b8e2f0c45045752f4eba1fb321b5fa9a3e0d5731762a8ed67f431c1d929c4ba5a18c335a694eadaf29334b552bcdae9b215aa72787a89c415a692ae8b057e7896fc9f35c6d8c255041cf817e4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170e6a4e49efa2bbfe22834982a881ad5e249c1ea2ec20801be7de8a73c3ae380c056a5be9da10754effa854ba3935b05c9e325c869bae4172e40529627df3bc16bb2180a38e19cb4255ee03933f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6db36206dcf32af858ced22cd0de4fa628d76e79c97156e6deb9c1cc966f76101c81c6e0b5886776cea030e8aa1deeee5c2b809a908455ace8782e1a62f18e2242a44af43990dd6b0b283a8c92e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8dd97ca6a8c0f07fd5f0cbaa874e374bf0093d6765ee7ad37f19d27220691ef052a0328b816e62e20b4c377858c99de46134b02290e61a0996679bd869cdb5d531ed6e913513b71730f1c3bc28ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e8626fcc58bc12a0e1f8e18ff83507efed608d6fe5063216cb87122e4a1fa0dd8d948c378260596228a22f37ae16814b55f97ed7dabdc5cfcfa4541bd74461872a619eef66b115040df5a02a6c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158b914e1859029b2a26a8d877168aaed9267bf9d99ee2a8edb71efc0b12d4b1c5b294d86f2159c5c749c59f04b30402a7afc451b2e0c107e2e11d0fc0649f5002eab0889178e15ab275355509d12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1228500ec21455cd2fd0c73f8a60bd463d738908a2eacf12a20d2cf7d61a55d815e45bcc484e40e59525c26e2736ed5285b6d1049f93896b77c63437901d5b3fbb28d7b4d84967934ce14d7e63348;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3e37eef812862758be46714bc1c596345a408819482b551cfe02ffbcb2c0cf6bcbb493ecd6a39761cf04027cde960beafbc2470b2d7eabb195674aac56a02bc2477b80ea22bda6f83b7275e411f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1067115ba6857224d630cf4593031455f6d6d99d9e1a952ecd063e0c70698df731273c2564d1f9fbc0f4da6aa9e28ab435e7d52e67a3ad3d60de97c91cf8b243eb90911b721f000e70e4d3f70e92e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h299c985b3209b768338e7de53e9e43b08cccff1c9e089cb6f6690e874dad38e5bd665c38ea5efd2169a537a22f770865235394bc09a57ea0bb5104eaf8db38647f60d91f1ebad75710ada65b434f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2105c5106143b58106e9a7d940ebad339549a56bf89247366a009c23c4fa1482227a1f457264971c9cd1e505985daa0d9e9db68983b3b9791aab0ed6f1bc8d018ce0396b0816b6f116100797ef13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf41f0d52963fef194ef030f3d6e1dd70dd2ba07c92d07a8985774bd329b7b0b00f7dbc446b45b071208dac27aa5ae843382a3b81ed0d7196ef0601e34aab7db3afd0b0dab024e8a0316ccf23be66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16adcab8a87f7421427ddca53e02073ac6976497c64d08573a5a2bef1bdae9272270f4400178d63f44492191447eaf7cebb692eeb14dbf94b5673a3182a0785dd953c462aa084274b055379c983ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfaaf9ee4961851485064b1fd583c6e3e811792c34d951f57fcc0717aa42813194296163b409d2f371e16da9ef78f778b0545987e4b7f33cdcfe9f7e0d519ab8908fb670aafa0eeb86bce5dba4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6a61803c44926ae80dbb91b76428cb7d49c6da2eb767049b51f0662a32ab8b359cf7237028cc0f20c86db9d34372454b16ac9341088e2c1d08bcba99743278b08e2cc8aaef3460052acd8ae6c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2bdee6ec218258f4f6b2b9607f06f0389cb15a4ee170f011aec1e9ee49b0d9e19fb1c838f1091f7ef3b5615ceb907327de2415709eb1e080b92a68a62c0ac114496c73bd93570128cca96d14f83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a8c5d4cc6d7de1652361784b1188d9dc7750ccdde5c89da5f4180ca0602b4fe80bdd29f51514537c982e449a39bb7ee94f22a764222ae006c9009b94db29ad9d5518cd1b6b10ccaa0d95ccbad55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ef5191c5d4e9b46a2bd9fcf8019c3f0ae31c213d6db1c84e456c1fcdce434621fe0dc1747f695cdd28a7caf2ad614837c5679c33cba982aa5dd3167ef3a72715d5c9d66c68c7eed0ef379d02b38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16eeb31274ff5d609d2eeb0a2c803bcf06b4e12a8f58775c5fd62ad736495f5c85076d9f76105d6d94df68d6debb0e9986821c7991c22b0dd2ec9fccda29d1a385e68326e610a37119d59a4b09500;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1694db4f812da6d275c44dc0047fe05e7ed4149eb571af8f6acbe8073bfd4649441b654583d5e7f94ca993cea9d747d7291a300ee3858e504868f442f0a86401bb1cba30f1bffb792f5578c6a0c0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1868a81689931945a8348e16804d08fd17ac69f8d35fc664ec158e4ff9fc6500e81e05b508bd073a54f68b7e36c9a5b600115ba955f816817ba3a54f6ecbea822f5d74324d31735dbd2ae07f2408b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a2011a31ae323f4de64d864c050b40965859ad854b08f38715b3a1fce167188dad1a9679728f9ed6da5370c8ab920d36f4b060b13738d044bd1f03321aedff2217861045451d49c24fd8fbe9b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d29d6b478ee5517fd61b834e00a92f44cbf59aa11cebf570fbc7cc6b437f51352a273a752e5ed9493c7cc84f39ea72173d246aaa88c651dc083bd57f9fbbc2a710e5c53830101ad35502a7ff762;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f16f1ef79f7e3430369b05aef0320f6e2268cbd275d99f5a570937600ffc844f2d84ffe6c2950987c49eb9ae8dfd19232733a196563bd8b1411d4dad3a8fabda0edda49b579a6ce055898edb9fe5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe03e24f407ee62aada73d56d041ee0bbac67fa3c0259ab3f9e334ae3f47f73d76ca7618adeedd20062cc5e646c4a0cf9abf61eee5cb907d1ab858448a5c4a7b04ba695926b99d5584f8d7c4e06d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0e94d815c57cfc09dadfe01e23a7e29f363f516355c53d8b98462d69091d82d00f937f92a8de331e6f1834b328f15200c7994c74fd9e006e0771243ba5dbcc86ae3e3ac0e21661734f593701ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6960bc28e228dcb1da1d7998bbb1597cd1d86369cd07de55562f6b8b0fffed7bb872da2429a9f7ce7e353ccd6b04a260d9b5986aa2cf78fa4766ef5a76a188f8fd41d3f7fd1524164e0cb294855d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0a1e45bcb42a2d22a1f5148f1136420e19f63f2f247ad0a7007fa0b654eba2f9905a3582e06628224037611fc87f178700a75cd4759578bcece1c32cd1cd4618ba0b4bcfc6f489b30efaab660d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9052c3231face8f1085c524fd0cb678f3ef1697dbc4515d8b3c48ba958190a7dc5632977f11efdb25409353e05d67910a827fbdeac9bd36c11145ee04e316d30e5dfa1405d6b62f32d6d7486ca53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b19b7847f83d3fdaa900400b6ca9a257479c0485949a288d59c8560db1eba076bfbbc57dc78de1d0c86ece5bc56655ef9e89241e7ab52d59b1ceee35cf80c75d23f317359fde1e3ae3008711cd3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe939d379fd772250d6003421b6701c5724b5b7b7af549ef5c6b47da79bbaeec721afa6df13d0923cdd29c87e9e47c46c1529452ac241c8bb13be0755c50cdd7193891368e94686a9d50511e059;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f8cc638106804edf572cd8e9c92fc4240643f60d043297942c24dd7721c4302fa28031e5917bef6c94e33751d8235ccc86afe2a91dc7cb93908bb106695ba5fc039646bd763704effdf9eec5bf0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a077c671c16f3defe77aba21fddbb499b7ae852a9dc45205bbeb78d41a477519ba0ecd83928d12d0bad26f372cc08c7a785fc29343441369c4ca41150b4d2e96bc9113eaffe4a0f64d7e03c2c43e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13be8b3b677ece04765148107d1f553f535bde436ec8063aadd6468153f12f1812eddbc71b05d97c028ac3bb2a478c40aa613d385e7e356c283789f9af8865efaa80b0a43d152e5c0f53a0068cb16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74072c2da731f604bfe175105ba7f32cf2b5d88355a5127c7382f63f269a1a7e8d856ff03d16800fa95816ba324518e6f08dd37913e68ca1f4437c89648553437dae64aa725a04cbe35f06fbf694;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117fdaf3b4674338fd5c8a4f445ef5a678ac4994450631c387098e8aeb70d133e7d2c312b44d17b07756a1fe3cd116e3aeeb8739812ca7a21e5720e71842cedf5adaf892a1d524d290c3dbec8109f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16561a23aaf9b01b8bc08ee2e5ce35397d1cd612b092c6d811f2fe99ea468216f54de9233709b6373b2d43596051d44aed4bdd526b04f4505038d947a93afcbe174a659395c1f875507d514004164;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2ec63a788c7d1c181740f1ce7fe931061e5cbf9bb33a5f5b2f824a77beb740de859e62a21d7a1ba180aacbfcb747c951b2bb8ca67cd5e1a6648f7c9824bf123d8de57031103f9f51e83dfd0274c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17af77c7d9a48fc4bc117402519618f99cfb43464879ce654ffddb0f25c84a365a5afb858dd8bb51cc7cd544b64ebf8766636aadef42635dbd9f4847aef09d9fde8db684a7849775b98c1c8ee5eba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fca2596df6f0a8fb7540ce9831ac1d1f95004e397aa36aefe7ac48be1456c5214bf0244d4ddd69b909609881cdc8116e579b50b0fee2d06f51777180e0943d6ada05675a0a6130153dbb6022b306;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca8ed59166566d6ead3422e068c06226a178fb3a2a236697da3444287dd1f62e776c695f04738ff2e7624e280781f54c261f61241d7d8062c55b34e24c5d36fce427cab46778060c489d0c391b63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2b5f031afc5ab7034aa1feb11e86db7386315109076504c14bc3bf9b23fe3024e5713c7cf0125cb32367e73e73dc9a834732eface4b3cacc18752f8c3e3a926260610ca6b18c565ef504b74237c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fec16c5c5bc0148980da9b14b518f8ce4d16fde345e5e53cc9dc7c276f461e82e1b08aa7b3d0b841cb88580af3dda2d7a095cf3da3ac75024f5b438957d10dc90600a7f71d3923ace619caaa01b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b34bcd3135e70ade1f8986ecef169832a75f362dba605fc880ad89c13615acc0ecd07007bc0eeaed68ef56508b840b8236f01c1e315318e8332b56a9b3e64ffab9d138c15f79d3a986a4f9ce9b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b37c02a30de3853758981ef5490b2721c44dd7e8f0935dc5caf413dbb2c495ec09fe216af82ca57948ca9c494275f1119daf05cb81a3eee934c48cae2c7bfd08f324e0c2287a6e51fa7752c87aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b6a3e276f28357f48788d96f7ca4ae00b4015d80b79c309b7c204e94aefd36b7e6cc66b6ca2650f28f88bf8edd5e4f546196ab9f68566a0be3dfb82958e49e12dc70d7822413bfa6095cf56c913;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bb93ac91266538d8c9182a65444089573eab5e3b19152f28a19ff42aae0a6a34468850b07a09aa4836375060ec50560c7f6b5985506516003c18ff5db2690f3cfcbe256259071fadbb98b11eab4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd73f35bc5733f681509b7e7b509ae5c3f7a507049ed28d069252320ac182e7c2c6a53e84cea65b0b7f6063e9c9eed04f78556bac82834be33d52c45663310530e65e327e0f58baa69674a5271325;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32855756a8785961629b5cb40feee6ef173748c754a2d2aba347046cb43b65c9c7cc4eedebf5f093eb9294ef1489aeccbdec3b1ba84b2f422e97a7d84680aa1a6610d08c96058438e60204c4d4d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5c4ee1fc5212f87d1967d91b904d36113df744ee855ce0e35e83c9ef7347b2f42611588d31a58878bd2c8dccd73f778b4a7ddc36a1cd9211f8cbf03311150b04a6428dcea40935b1084c4bcbe5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e903ddfef0b81bdde2e07973f5af59866d9a04def21f56d6edb68b31b1987391012d03d1b1d002b698960f886e654e05150f2610d211c21f37aad7d92a79745b60fb8e13aca2a0706f0cc437a2db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58b9b1b9d9cf281475a3500635396c1d885dc667a1fd99aeea50e87ca5cf58192bb9105037a5669b4a7102536321fdb823595865a8e3bdb2e582f0317383072fc646371c4c81f363c1629885d237;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186e5398ea0391ba43c44329cdb1cecb64b48e2509b0790701ec064c48a023154b01e785642a2da970bc0a09e9dbb49981625e68412e6aa334b9934227daa0f027a594bdea19240d78f8c1a157309;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7a6a9943874a4ca97f2ebf40923785804f249ebdd983eec1e6593e84de327c3745b50107bbf8908353cc9b9bbf2583834afbdc67fbf720b34d2536ca4747fdf42fcce642326f123148c8eace5fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbc9dde8f5ba5243c6fdf09d94da3efa9bf53d31e5f40174c7d9a2245d707c8f5981c9a24519e89c72689eb0cdc1d3f2c9d53c0b581c9d8641c57d24655218df07cd4f03339539a82abd1f5defc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h874b13c5ec26ce92f92c669276ba2f70da3628220a1ff3f176775cf1cebee60d87d1f586e856f8c20cb4805a72ea790094c276892522f676474112c8de392dceea822aeba9306f9dc16a41fe519;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122fba8e29d65198d6674c3b0ce79bebc2cef8e018a0c815ba141ab0cf8eabe03fd7a095eadb805618d7de25c12a87c110e8369436dd39f8d482dcfbaafd06d8886302373a034c9351d56e02bba34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d04990684671ba7a0fed662eacd6d7f244275c2af6ae5efbeefefeef027cc1d6d2c3d2c4b4111863c18831041508b674553368bfa742a975fc3e35a713e95a7eac63a89c6accbe13253ebfe5006;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c0fe01d9df13204518d3f6df6116d78e8237d9b77c18bf1ed6355e9d36f77dd42c2fc407e145c08f2f181eb8cf3f067eb81d716fed8bff45691d374deb603bb76287ccb6ac282184476cd2d3d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd39b004b1fe820e3fd5f87ee1d3aea5c31104ee47fcb2717e67edcd06b1270bafe02cb620a4ee17741797af2fe4d3947ad4003a47a4dc31fbd75b2536786c46f4934c14722a839e6cfdc010d2edb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a9628a381cef98bac472dd2dcef030af6ce93b915f9056d729a649b69597021825968076cb7806f1ad17688f3e296947ec0875db264b323a3824de202cec034d01fb21f7594b6a4d6b4d7341c1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he52a686d7377106fa0565abc9a3e6b8bee0c43679ee852ea9c2601a8084cb37e4587ed0d520096cc9f5da854a016a4c28de5dac593bbb3b05c15941693e1c6a9192e93c27d86821a4bcdfa86022;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7d2fdc4c4efdf0c8047162abe737c5b8e28cfaa09f2b1283900a4fca844385b9de28fce1ace57b7033606b4178c8a4b911502212a77530bd6d03e2db520c847552e715124614c3e5aa0e5cd40ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4772044e71650d5383caa32ef0ffe6b2f159084663967ea6162ac3c53791d0e1515e3b3a5321cbd7ab8b005ecb21e75c538a36e7b147602100a5231449b8b04bde36a70187b8256903501a914a63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7c11e0b1c5b48383557542862550c3e4e0e93df8a2d8dc59fca8b909923b4691f7fc6c7297ec7a727cb1dbda33cb5ff10c7782cbbb480fc34b4110a1944d61f179f6c4372933a64f3202b697a9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1895a07ab05fd78a89f0dfecad2020b7d75430def65fcf9dedf7842931c8d6a47818d34670b7a8f8b2f76f8865415c41b90d4569a337d1b2eb80726056ad7d61b39e3d948f0634c8f44ce5fb1d548;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c26bbc40902530921588e14f3122928d13f52ef303f2af635bee1ef490029aeaa32140ffba5e695e867d2938459d7cac9202878824933d2c82a417f9596f213c3735d1ae4ff6d86cce7968de1c3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146ff0118561edd2aeb017e61ef341347788ac03298f0c0f20e43c1badd01a473c044c9833dc149c7fd4bc2efce818a82c23f669a27dc864f4536898cb703b67607e4f32becf508b7b99b0876c870;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c51cc592cabf3d62310bb886867759374c81e36781ab85ff0c0c932295751269f4b6c8a6b7d333061879e119a438f1d5c1451f8570852cc2c42df101453949026c4d585f97d61759bda79043bd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ca5e75e4c36546121a285d4b8e143d18fb4b5c4a6f305bd857eb38a5e249219728d9c273c2922a33e55d8db4d4374a26c45488ef87c09e0d996f947624984a15925bb63d50c6c14b7f91f46d3c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4c936b1f64f47ac297295c24edd6473f77fee36b0fde37f215c621ebe30f47c2441fb74f8ac6bdcd866eaf715f379ab222e6ae03e4d7b2c06baf2646c15dcceb6ff900fe120ca0a12448fc52733;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3a209c2536bd053af45755b8afcbe51f6a55472220879040da871a237a73321050d64648a8224d6d8fa30890af73f8d36444934d8c77fb6546e2c85e3c90335fe5676750f45389658fe64a51fbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d6c7c392a07c76dd3473fabe217e1692805ba823cd2a79bbc0ce1454633ac14994992205852b6e7b6f81afb395613b9544afc66012f28cb1c8d34435eadedb63602672157423f020a60e777093d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f5998cafa47cba134723b529f53074918c208d09cb5d46d31dd6d63a863412f29a53caf522fc3cf8ecdeb00595b31b79b04022f80d0a557977d79d28eec4b0963ab86723d1de336a0e9189e0397;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaaf19ff85c04e68b6ae624afd6c37d774741a4d1b413d20211696df475a27eb1c2ce1662f11eb3bec877e256a9268dc1a7f21e2a5a1ba6754f25b693a791ff558439b9a478b710cc0ab4daa4d9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb1679667cffb84ef259ff1dcfa465c55d2760b41d1a06c72b674387e9da7df868f04b53860e1a7a6343588775ba95255b681f049bb2490dcea84feb11c3344fbfee09116fc93f5cb5376ec449de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6f5ba7f4d03fc98346d6b34fd2d7ba6ea1f922db963c49e747d96dd1398ef2fc1703b6e731ebe37c44b5ce01eebad6b9ae4e0916acefd2647a4835a8ca1984409b5cba23bb43eff27be2e7489c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8bb904f51af259fd67b254198019c1a84db9f1bdf725f4f77edfe96c59483631ce24542a18881c468cdbed768e270b837f0cc4e16c5af68e863b29964abd3d9c05abd086b781ad3a65f42f5be92;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c7dfab4d98d1b3e3c01d5c99a0b0cdbcef9b13b33a907cc3a59f72d20a9e391452f634718983cd31418bb32d88e7cc9fea9f9f7364e79927a257df8de649a83483303d3fd093276d92c72f5464f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac922318d19fee2aa76934646f21d1ff93bf65d7ca8765e2c118163242cc00d5c45c9601ad5a878be1ec0b9e1a8769ca8922924bf4653d5a9fabe6bac98be63e7494b76ae4260f775f1553f4e9e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd0951840e09f51a16439ad46f361c6f7e1fec3e8c65e1fe4c4b5f55e254eb96f49eeb628db938f71c873a70c43b2b8c601d302c8e88a2325fc809e826c22b1d3a481b72355bc5dd13890f5f736c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a6d7fad2dd9b58b956df60f85ecd55ebc3c7d9f951908f80e8fb37acb9e4efd29593d2843f75a96ae690803ced28419b585aa79a7eefce3d0eceb70da55cd5aad9975414facf3de4cd8d41fdd89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbcd1c0956573999b392025bcdc08202b50fb8677d9a3f929ec59192274b5bd482b8586b5de01fc011d176d2dbedcb93ca6b96c676db0762dfcf793f54bdc5ba4f6b4c7c5c00141e56ad28c45d3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b445b00b7af09f35306374531b792e3f6c11cbcddb1710f1c47b6bd38da93bdeab096b29c920febeeab9677a800418bd92ff2eb6b889d429254594b3d8191eb2ebc98187c10d74b8c24f25212bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154ed9a573031886150fc05e49f868dd8c653258d9195559addf3e7f8856e70b59ebe8c4c9a3a2085319a4f90a9e4a37f91feb621e294d36eb081fd9b7ee822839329ed8307c79524b55ca75b47af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ad7e7bf77f2ba99522a1a7a82bb98a3429de73f230038ab7027b6399e695c567231d3120ded715458b20f77e2a1de88c212dbf48d8e85065fe66c60f7eec34633109ee8a089e55779cdb021fffb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7688fc16bcfb7bfa9bf46e316e86b5284662d2d88dd1414c4171e5152722b471b08e99856e83917cbb7e18548d84ddc36e5aea423039267e9432a2bcbc33ecd7d2c6e2f42f58fb69fac183ef9009;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c8e75822df9642b83ebe1d48422f7b1baec8fb88334bd74867a6d1c2fe2474db15bd3d8bedc8eb8e36d3cffc158aefafac9eac79d599b2a8a465d38eafe6fbd5c0bb4e3d32b45a9cafa2072ba7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20ed3cb22571d11f55a33baf6e16bb9334fcb233c8ff2c51506217b05a8bc4e626da2224db17184303f78d0f6fec433cbf849ae8d3dfb0fb907fb80fae54d3b429945af3b9e7f578446f030ef656;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cdaf574fb564d188898485b22dd910e298ef8bb03e8dfeb8469f3b2481f0d879331aba2833a41ed50e22c5ea7c8cb355fe57856dc36dd5b93a530226e3d25fda02330ae79a0feb8d5afd5da2b651;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb835d05bc8f9b2137488af24ff294faea3f41959f0343706798efb7e1c0d8a78cc20c62a592332ae39affe347f132cbca0a76393f35d48e68ecd0185542bd6c3d1e8676ceee24f3add3fa167647a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5c37e4cf183de4eeabcf1ede8b179cd1338848b5c97ef8de539e628171a6169cbe0c4a4a0c14b2f4cee037140e21529d8d1907d14b226b2c0a2ba4bdbd19aa065b41e9292c7c3e2667b6ee3fbb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc65f4a341772abdfa22a63053acfe8c7a41ff3f37e8f3751cdae32cff79403031e7e791b83ca45846cbf0ded3cc7e2775229d01a09a5977422115f55564464450b3fd47ce219cfa80ba1233e977;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2aaf60eed8de6188dfc86b62515ee2c214a99159d47cfb607c588563deee5535b50a841068fe3b5ad49d507b356187d01cb8d905060e4270ba96d9431f6d4d911b2adfcfbf1dc24f625f2536f86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11dd289e7cfe371c4b60ad50815e6e123b6da6cd60c19f426ec4a42d98c92d32f879ceb62c31ed025f1f5ad170e7819b1b408ae230f0231fee2df799172f00e5ae478ab4ea18d749368db8b5bda6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b93306ac508aadd31d9022c3f1c46b4490b66b674115a3ecb07d3b6a72c5f6c4b59ebbff985c381a06634dd4e308d07a9b766eb64a11ffd1b51ebb559b99f6ed18303ea6dc1114efd927afae2618;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h877117a31721118ab69e745b16dfd4e96af741a2b3ca7c4ce5b2141272aea9f27bef335889bc0961f9ce53823d7782e963c192773516a7ceffaaf1e61583638c34329aaebe282b87308f65b7a134;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42a59f330ee08871ca05e0d2e6a3b15981bf9ff11dffaa006840a78ae5b97a04503784b85db844e80c0c93db77543a6f928edcfb94d42b8b760a2aae101badb38635e1ed0048baeb2caaecabc3c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d52e0eac37eab4c9fa15fc5cf20756c0780b6a95bf2d37e30ccf16629967951d1a5569350546d7c766310dc5753d8b7f15f1de7e2942389717a63b2dd0d5b5686868966911db1a12cecdaa6b554;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf306be73cb043af47b8d20cd1de120d40631122ed8191c3f26e3fdbbebd9f258e8e5a832d38a982d0859dd6eae175fe4fddd533cc04d7c2183c96f5e5f5611503e92a480233050e948dd2d4cac0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4acb8ca913f8199852b2c1677728e150b2dbad471aefb7cb3e464616e52cc600d495ba3bfe72056c839768edbb001a378e3e4ff3b897f65520773419ed7b460ef5180816c0dda8a0139341d9a44f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcaa2ad52a471f774144817b9d6337054b4f918bf40a6c16d648ffca47819171909878d6dfab092ddce72053d39e967a926a44895223dc19487bd60fed55190b097f16faee7a3d28047b91037ac0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a287fb7dad6b849cd40af4d00837cd564e3a21cae566cff16743b14553dcda1c959201d12b6db44e782ff9143e0048e048dd4a24ecfdefac644ae809852e1c8d6aafb693034c972e9731976e6a11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c7b571eee633e14e4a6a9a350f4d26f96e5421c0762c9a8b7574cb65eec78507a93032333a20707ee0e8639febecb9bb886ae434be2c444ff424237d9732734d4e28cc2ee8babfd454c8b857f89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3a199dc3484f7da5ad0fd97d26865401c81cf6329b557336f2077dc6f65134564bfaf57a1e90eb8386f09b33b5547cec9b99a75869813a2ca07f93b9fe57dccc490596515a12e16783678acc7e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a965132a2fc5248d26cfc3e4383020bbc58b496dffba0659270e6ca7670c5e874e45069039647926ec83044e86b9410d6bde0b85445f4a36a5b00e84778cb020bc05b52e736c3372aa01db95915;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d08e1e004dd183b25ff163e5e7eb1e2c3025db080fc6e4cc81f6d25cf40a927df9ad0d1051c9f4c2c3abe9de41f77a60bd417c602b7493416e1c45789694a941f1264eedcef4423af73ddb10eec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158c91e93f548164108782fd8a1cbe17ade16d15c703e90f34f2abacfc274f5707326eff7e990591437364dcd6c635bb438bc9e8f2fcbd9d1f9a2c6d73148223f39cbb6b7048c6940168d9ff98b6a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7d335032bdb1bf2851739e67d9318f2c69fb3f69643f61b79045b92147b395f821a06853e387828cd93f742009720013db122071111b222ba84ac41658e488ac7695938d36e4fd7f2ee8a54d3f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4523c9a139fb75920085479b9a74815f05fb290cdf309b1c31eedf7233ff6fe9745035c1553815534769c35d241e09f4f7122568bc2571472b7f4de3fb90299decc2c0695921cb5c893fc15aec14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b3277931dfb7021299ec4b0d3d0c55695b9bf93110136a678a04530aafeef7a9edab89b979e5d1eeba81115195e9292e074e91f1305aff8951720f3b8b63b753d44d98b4a2ddf3c3d6cfafc124f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a9242e6b8be7328debee5eb10af2676639987619cd9c032038629feb20baad2b89d1ccf2a3ae5b442173f2a1860ee9726a7881e521e405d6c23ca8bc1df02e26fc5b6dc7db3eca8d0e3590f7164;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5531842f4b566a327f38263108858c004502e1b477aaef0e1c92a62441515e2addbe82ee8f475508a8cc7a4d194af67313c30a95c0f2572b387fe822561a445d9a03f34c2bf4ae1c5fcc3502849;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e076898fade82170f1f1e3a35cdb4464c4ea98bd2be3ba4909599b5c0333b818f319954940d114df57f504e08a2957b73ca6fdbd1dc83270cc410f2da4cf23b4428fb55659c606da93632d75ca5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b31f4588534babc2ce2e45b1c4db99a22d3189b83e1d3a19acbf5669299b308c9078cd5acd762e900877b7d8357bb69c5e89439048e40d90297a2392a17d0923fbad2595af1ef6bfdbe8f90e3b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b9804eb3ea65f5cdd3497f568303de3c2688f2dfe198ddb1406210fbaf4074e8ecec77e1a69fc7fd98903ac3b7acf6f3f2512a324bfe1a45de6874f4404746f3b93e61a68560a93a5ad346d668f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e2fd543fc667ab78291951c9066f508426f0f58a810daa75bc23fa5bb7319b997455c9dfd07110ab99d719dd4c8a92a35308a2c3ba8a86879d40b0ea25bde10f40495e7a442d5e6329bbe17af4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d76e101d464947802bece0840806c3f8966c8ddea515aae46b9edd5f1c8b0808abc030feda290a09166e32eccb7b4ee2d912c37e9d8a1bb85137474699cd920e1185e3278ab54252f14b3da8f8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ac41229b919ba1a1935f94a3b5e681fde3213bff3aabfff419305f65a5501a8e9a29b00bd0feca0b096124c996dc4fb9411882156eb61ea92f997dea375ddd0de4bc0d68479629139726d3f7642;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6f47b902f020c1e627faff5bb66c6042a1497c1690de196acc8f54efb45c28c91a14d9e3f8d6d810d326c6c4fbda519a73fcb1eb0d167e1bb1e9eec7ab1b11c5f560b9aee79989e12b9f9681d1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172fae7526c36c2e3189470a100a639203fdcea2bf22da30f0c49061ed8cd68f28e96073687ec01dcbc4fd745a4b0f36f9c33e978ef895a2fdc6ead9fffe4d87d27a1fb1bd6c3162c0654ee5b5ca8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0e040f61700541fa3764968b87e0051999b90286baf3288eaa378c450ef5acc8a506514a91075eea0184593a9b4bf532571abc426e629fba6b8ee298fd8ea48ee6bdcd5349dde04db27baf3316b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea1e2e4af8359a3c5922edddc3b1daec105dea601819644fa43421a9154dbf19f814dbfdab713659b8273b9fd8664b3eba426e9c9259aec35ce42a009b8b61a363d8aa3562a956faa4164fdda5e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2321e854475e4916bb9f4e0eb4cd6978350c80cd684c5e472243eec38a03540d369a5eecd75eed26d56bd68f4122c0850012ffe93a109d9a77401085db8edb43cd2edea310b157ebb15a787504a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196ba531532b9f6bddd09136d21002374790fa937aa0989b3fdf6c8088e24d3b1dc4a75cf40450ea44f69d9c0cac9343e67f0be24eaccd95764874aef3b93b510561273bb4793964baab21d7e0782;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f97adbe39718c757be279a92349eb258de675fab24d9cdbeff16ec61d6c04cfc8dcfd43d518a317bbf6186c209367db6dc6fcf608c6991f773dbb43f4a694ae19db46debc03cc9581dab4996aa1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23edd221df1944b6c6a0ef5a796aef1cb03d805f189defc27e075eb825eede8689eee078d19d668dd5e1acf8b7f24a9939c1aa7f4ee670483081de58348ced94e4ba0f0d30c507fdf704b01b9b59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10202e5dd2cef683b3786c2e0456cc6a7da68740e8bbd98c7a6231b3b276419223021b09c441a111af4ddebcc8257067db8c6460de76e7af140cc096b36ec769b31f09ada50d282ee6392aa9a63d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a29d5f8360799f526c8df8986229754e1b6df0f51ace323cb1271a1391d450ae64c277d9f8413e3f719d8c0f303594914335f02ded210e8f700a26b748b13bc1187fd4f29bc1444f96c9d7c0233a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb5226cfbf18def0b3a852707ef034f9560c4a7626f4ea94d1bcb397315a8b5dcf2fc3f32400b9599d56e07d1e00f8ddb59205221610403089b772d9b07894453c1d19008867e86d11a7f42068ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c32eace69ab5d674962c0bcd6964af7f2ddfad03cc7d364cea4b558ab60e35996de23584f19873b662cbed64158625292eeabeba9baf1415a81cac5b49481008b0f25b4d1eba66ae6792c28aeb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf4f46c578a53ec26ca301ea025c2dd68a769d5cdf760f175fee35d34b171d4a93b4ca5f71b38d9046cb664daecf82334815095b9878bf4e66774dee64ff2454411c24d902f1d5bf5111c5c2d709;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f3f65bb7ddb8fa9a3f9dbf3d695b0e63fe2b2660a0627e0aede1a799e82849f4b2c229e89d9dea2c44bc9e17d04d7a9b927dc03db65c58872b7ef0522dd6a4b86ce828546b977d401d6c215e760;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16679e01cf197a18062fb81c2c3015e1b230dfa26993629454857495efd0d95a0d926f58427dec496c45aea08534539702bfc78aaeb04ad11536ed00f9878312aa7792f355111da7cddb75485cc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15740cf469a32290202a6fb48ee92872aef32ff1fea6c695995dd92ff813d0ffe3da17565d36c29c835c9e52f1592a773d5186d43a318e49c746f5504610258a15ccb3583dc8c8f09b2536fa14848;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2d0dfabe12bd03f8c6dc2e8ae315dce9017f904ac57a16b10bb4632a74bb8dadf3db64f1fd8bbf79a55507b5fbc089b08d94514fb4c31a18df1438fbb049f2e705c7f677a9883fecd81ab25a03c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab9c7cc99159c1094f853efba3e18bcd6a122ca65f8482b468d5001caced846f5700c16bfca909226441c69b667bfa24c3427705420f1bb92cfde008715c541f382e728659dc5f29c98df05aba87;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe3546785b90c38ae813afc8dc176bc5bd6c1effc5534231f1d080e14494d58a81cc33a768c26aaf9b2e5b5e4f9ad4d94eaf65c62f91a03be303cc6420529ba58215144df83037644571303b0e2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hedd910c7ac6bbf3ba0ed2a4d84d924edff06a77deed1017ed3dd5a1b66227dcf923105e16edba9bc2f75085249eb75bf216f99508f3d1854c238b416648783ce5e0ee3f22f5af3e7fba80d20c262;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56c54b4b3f34b45d615c8cd6fa00dc039a5a07a38ad8eaac75cbdf36ae2be4fe71003062e480d553cae3f880db5967b85158340e2d438fae4313310eb73b02ce4eef59292f9dd707ecd2b16d9ee8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a4014eea57330a1a097b20acf556cf0c0256e564737f14d42cbc2e45c6f05baff707db72d19a5212a5091d547f8f3f154a8127d81f19679a620f26ac756a43ec6748110a71add8e6d8a84b129a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3e42047b3679d99063b475e378849758c485fe40f9ac930663129b5ddcae1e2868a9d0e2d758a3fbc1fae6f9ee105bb215649a1dda47ea80d04815284a64dbb8759f58c7a4ab439bb42aaa0e600;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5d378aa6b6c915ef13605596bd60ade7c1c48368dbf20448f3f9a4c485339de9b396b090d23cce34e06c30c9bb1433e482e5a9ff9a5e4c534276ba8a28a1279ea713823dac86a92bc1894db47cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43ed1f91f2ce4522d25401c00e7a7d8cb9d2ffe0717cbba78c6b8bcd22104d7b2cf152b3d04946eb7c3f6f4710100054fcb41812491f2c3bf4795d6a8262f4027d7c5e50635fe904843a8d2b3bae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae92716ed5e61909ec00d43b25e3a51862a3f7ae1d14180d1cf504f8d3f19a4e548650a11d86b385ad08784517bf8f00e8aca90cb1193b736c6483532ea3e298b45092a9250a216c39460a7ba351;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f5887a4622678ea823caa56e385a48ef5faf8cf1676aae42b67298ce3f47c361b91c924a42036eb207c97e15cd35b35ade28b3e4d64d5ad1cea83d74134bef327c8d9ab3217000658f2b6f559cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1a62df45abb03925c091fb1208faaec9ce92b2e8976a2c9f8c7c381938e0762290f4674a7bcc872e6f5ec9264b7217abc171693d9976637389cfbc64311d949c2ee06c5b7a2eff8f2804dcf4e97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92fc3597779215c3876ed4647722b77690c2c3e171fa8de302534f24b7ea464248b049dd1a903e871744a9880246719d9b8944a353a04a9985dfd775612970203a17a46108eb9a874ca26d6b1ca9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e34406fcfd84fe08661329e123cbd65c74262377d87554f8a153aa30580c00ce2fa5eae258a5de50ba3a2abbfd876a5a746496f8052188c9acfc9d04b26d7afaf541288950d7dc963ba2c55c3f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ffdffbd76723c3559a6866ffbefa0b31e40e14e9d2fe7e86f7b22b976c7668e8a92110da418d7bbe8c9ca3bbc5a1b6f9249d3fa82f34f28192c8e7c65343643d004782065e0a33e034ce30dad1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1724c90b7c53fe7a940b2494703d4c192937e3e33ae82d8f771609365f75ad482fc961e2add542d554e88bcfec75c50436447bd96c6326be83f9ba07928ae0abead42afc5f73172c219b7a8ae5458;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1486a7cc8ebb6afe3961a7a53c88083f461364ce9d317015cad48e5da0e08ad6b8b3415335f2ee96ff4f638043668756143bd0d90b5250619466f5c70ab8cf7144b6a1956dbe6e089b9dea19f3e50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e65636a6a4b1ceec782c56d092c1814da715435a26fa1946a0872e71508be2e2c421c33d3620c75e31486b1e8550d6ca57a66c3482c851424f7bdfa30b5a8955f6262091fa2691bc04270d82c16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9f021cb98aed8ab8d0fab79f8081e4855e20314bee4ccc8f397e808dab69078012ed4c0a10ec9828be9a6eee4a6e0d80df7e6e5390d4e760134c4dd99d48e6514fa0d22b90dc1fa36fe9671c600;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176a35aff0baa77fa39c18d62a805f49c2401941c583ade7fb16403e4053b78c8c09fd554fdfb0c9673e6808befed369a3a5c5c28ae2f7f605e182c584d1bfc09ec999596d0391dc3c83de117d317;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf95130e52f7c65c84778fa382b1d339ff0cf5221d42b3ec4d1acc7f0fa8501c2ad832ce2bf006888ed7cf7262b85c5085e7df81476d8230b9de9c7b18a3b8a29f4d9422c6843abb58e72e2f06cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1672c13b698e5bdde393366ae71702325a08aa181d461e17f9f0b3d6695c13b2850ab3c7ab2b06069274691759b5f77f7103ea5821d1c6099572ef24d81e49d0e4b5aa33fb320bf2b13190ba2e6e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0c8f3a014751a5260744f4b61742284974532efb8de5cd23bbad6881a14265aabdf106fdd9a86c4e5d57dbca135d89437d6c0261baf682804d0ecd5b14a941b7ce93dc7ff99c465d9ee60480b59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19897b050b44861fb04cf372311a03bb41f3bec12b7941527f7449fad16293d115223184d92c2eb524c5738d7602dbdc5342a778d00c3927f1292e6be9da8029b90b7885427a606a600eb83834969;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e42a7fa1c180544a65c348507205c1006b5118887d88cbbe4ff6067e4d8f5d7488cf85182bac004b88fa624a33d0504608346e4c05824eccb9c69121c26be9c57657b635b1b4c4bbc7bcc431b60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faaddbb2d9f8ceb1731a1c39c175b7d67b062aa0d809c7805478fa7df52c646e51ca7918ed3663c3de6ecf8d5329c02aaffdbe3fb1bd9bc569b593d504d42965a17081d6543b2d26583e312ce723;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4679d29e9d08935dee5eb9c762917b17ea15c1754039af0a16db71a08602377bf31a6e5e97898366ce3653e972e83c15d153fce594c3d810e397b09f7481e2e64eaafa0e6732c83749839747b14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb51770bc38735467b824ce3aaffe137c9124ba49d15f582262908d576442221da891d6efc877b497796c09582a9b5fe17903e271d80e44df328357ea10594bda63a9c580c7bde966a86333a33674;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcab7b27958cfaa0f0acf0ec0f9566d407cd10cad419276b56993c900d532d6d095d7d0863737adeb6380d525eb7647fdee56522c31ad982f42458df7b34fa0d84a530c33d9a85dd4f79cad0f9ce7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1332cd6dd2a8a9ef134c8ad1487e979de38d35703b9742b230131f44fd2f5aff5c5c41e6a27fbbfac5e4de83f8d3c7f01a8e101de379f6be716091945fd098cad61036533ec5633edd403800794e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ccee252fd558f82291013990058e351d653ee2b2242abd16114e7103f196a1cb2505008c6675075b409923cba63605d68f2bceb507fb2f2e23787e812698e84a6f3d0a2159af668bd7e28ef9bb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4d4952bbb28bfbb5dff41823019404431e05045f562b53736a776446fddd1bc647a68a3ce6732501dc8df681371c95b818841d9312d01cb3a46fa4436179540c6c52e7d8deb00db62640ce338a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150c96184e619b7e47ef918a316a6879c1cd7a5b33a7358b7b47b3a068f1f62b4801c9f422f8bd5f1418792b0041d380f23fdb90bdf6d8d96fb920a6786495268b0cf45affa3c2cf3d4457d54d11f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e64b44a1d2be7876929f68f7fadf9af9235298293df5152a9ec5d9c5b889dfed423b4f6fd6ccd1cdc31de4c879afc2a8ae8741d5f228ec228420cb2edbef6d0d5a48849f88b3226ac8a4bf9403e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c0e00736b683f6ef11e562dbc5875c37faddae29afdf021df7645b659d709fe6333087922dc3daa98ea6261c7b7e47372e6f0da0bcd2b7ebb01d0455a70770c104689c93848edd2474e12954f44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d9d8e1c1fe30ee209feb93c6c77ac56b0173246073fad2c466cb32799c0a0761c49cd8a25e829c472e4da877cbf16c514eb0fef46be92ca283a030f284c999117f475a6ead521f9fcfd8c70d5bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f200b84fad60934b44adcfd2b6c9f513e57ea905e097c6435231405d1fda9b991e40c63cca9c926a7e4117ddc4bcedaaeacbe559ea1fd8b61f3a11972978475046e2ad12202cf4a03a06c7acaaf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e7113c9e88a3182e063ae11b0f172d775387c86bfd41d17a5ab3fe2344e4211bcac0e6c9f805410d0660e11ba6fbee659377f0462b33aa26c2fcf3fcd59f9e043a653b613ee94429d4d806cb9e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3385d296b075f13539a3d5702bbce571100ae284affef15f077b9b70d34bb794252fa576d1e8bc054f0f9e1e3e31b0451d8b164aad1a52df845bec3f46ab0cb27573ce726b39bd95e4c10bf31f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbda053b753c9386b8526a610c19c0e77e2f0942bb970adb58f032087f30e0c2b19a6856007a789b1bc5cf20bf8a234d932db8614f1317cd68aafe8af45dcc11e61698203f808cd0d26e5fdb9a573;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f0225542fcd2b0c896c797831dd646b08db5f7fb70580e85ee9c726e14347999bbbebe849b550d7dc7e1e7793194d88920ad6bc001c41bea6f1b035f1cd12a7d3695ae311cb1264756bfeb3ab5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188189b23e12df17502331e56ea5040d6a87667b9f2112c2b0c4d7ab504035d9921e2b8375265d3c0777f23b10294cc0b9d704c6ae0b69f78a7dcc66d065a276f101fdef69da9bf241f7ac7baafaf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcaca3238629618ffe2f37f6876e03ebcf9ae7e84694204210b5f5ab5914211f0a4e399d48ca111b3e937cf698395d0599fe13fe6878651dd19919cd2332da4d14fa576fe0215c1070e4256b7c500;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b6ee0a56ff848a8a07d5fbca4220479e87a659bb5a2d7367ad61647b0ca36475a245b121a0b009bb7a31d2fc37f148ae682386963b2344d96ae44b64a8482aea94a7d37b76eb1a0c6adabea81e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he82e3f8c754a9a51a8328e83f545e65c3e5641784da4ed1788557b92c281e8fd79e5d949911caa1f5e75049da7741caf9ce61e378e13f6bb8b3b80a096e334c03a6309e7a268a5699c924a4a010a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fcf91501891698555bccedc4ca5de1604d55fc9aeec5cac24412a68ef42d43cca2442955761699f62c01f5c922a425d3645158a45d9cabf3b660b9e2f97b75eb73dfe1362ec3f8531b56bc8e9fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b1081d0474aabe9091017fde8b2462226786ee59e20986dad78ca9947255795c6a6e4b39904cd28d564eeac871d3b65d3c9f76b7eff206fe4ea7546b31da9f5bd43fcc8619ff0902ac6b608818c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha05f376c05255fa0cd122ab5b754c7cc99e3e62956085976721a80f18e52fd29b8c4a6bf4481be81fc655751d15376ba392ac0d78b492cbe5335b81bb858398fa10c755c912e6308825ed246e855;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h507c02334fe4953eec00ce066681fb89d5ac566a22629884c8f502ddbefec0deb05650abe943b3cbba08db9ec6b1b19555ab4bf7895a11ecdd0f09a5276a166a3c149666141086edcbc98e338d50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a6df56afd5df398bc6ac79d7ad1cf142f9313d53e6504d877a1d6f0b5fd546854ad7ae773069f9f9658768f4a95d0b5222cd720fad284eb7ff5217be702fc91334ada59c80ec7d6823b57c6d714;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fdae6112f6949a038bf2d2249a4ccd5e13d51546b16ec19d618b6fa7da4099cbe3e3a1f2166346e316986588009571057b6824ec59edaff7fd8f536d5a0b06c385a6f878a710970833725422aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a46df43b938400856b3522680b988a65b02d1270dcf9816b71cc0722c348aeaa7965ba68677fe93b7bf8945c00bdc7d32d03b16e2b174f669862ced5b8c176c88be8ca899799517226e5d7a22a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce23e18c1eb19d4799b5cdf628c7fe1af36f8c7b74513e2dc2c2a49f4c136b7a1269f6eeb86ede210ddf46c2d61abf5ddef28f8bf46fcd1caf99703e4c3f71c616ba9e68449df07bfda9762fa599;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bfff27c6f9fe79721d8696223b2794607e2df0aec86f6adecba7fa1efe6f472b397197fc11ff1309a425d611c08e1b35c19333e9481ca0e570e18d8dbc1104d2b32e28a1330c5f9b6eea8430064;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a10e80354a415feac1e52805e553ffdefdf72682dcd88bc90228754f0af789abe8825c338bb3c3b2d7efaadae023e81d7aded598ed10fb99c1b41bbe66fa6a2ac242673e3f1a7563d5b4f50abb58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b2342473cb365daa5545608c60f00c351c2ff15f92bd61806ba8954266e42f14ed1af4aa04dac73b810c25982a69456b9baf144b8175ca61cb876bf874f1ede85c0657a5b612ff735ec3ef7452e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2964e32235b7efc16b169745e0a2a8c19113bd91deb40c25038ef4aeade3574052f8879dacf74b5644fd615ca6668a01491cd4f8582c4bd8a338fa31f8d7807b40f3caaf01ab96c5ff6471cff9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c613c12614a1ab6b3d3c7252b7204c4996fe3b18572216c7f1af070e85e9362d7ddcd2a37128a40ecdb14c441a992b7bc30b377cc2198fda959309396ae6025e517d93d0fb78ab000839bbd0fb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc981ef0decf2482ae45fa608c84def0f43c3dfa1140aad4de0f21835e04f2a1bd5d472b2c931202e4b25bd8000c31bab6a8281baa7297f6a1800bec220a6f215cdab81400d3e8ce2e248fd135cf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c7b5bb6e06382bda0937e0cc4fe2a72f3551ba89ec728be4061527445414e37c5ac5cebd1a1cf590c931594c0453f84f7487403af1c6455872b4f831003bdca1de980243ef2d81d4a5bbfe19a73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b45192cbaf219ef7559fe9b65a98760098913400d2668c4c79ed30ed4c61986508a04fa9adb46dea58eced7bada1afd9501778dee0d19bd3d6610c01cb6af36c31d3bad2c8eac28587e2afac1d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f95e6a4d9b2ee2307bd8964a4cc8bfe6533486c0dc23df4518feb10e6c3cba97f3cb0f6ceaa9964a2b6cee07f816e461bb19044535d73bb67930b907005fc7ee9626d3ea6c868ad65d959682793;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fb4888a7b9950ff4696bf09f164ddea4fab17b1bce960e0c8115516412f83671d6f3f5eb7163d8c8342e93a25342a032295ed241813a35db2d1ed1224dec1b4471a7ff3cec03edf4d813ddac195;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h569a40a4085efee1cf3eda408fbbfbfce546a4a0c500d617a19e4d8574f672046e7b5787323d5fa65cd1cc5698acbd0c05e32fa233faf56a9a8272070fcb3b1ed2238ac4247e529c951e4e35941b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1094ee675aa95bdf2257662491f1aac4d9911749566368a06bc4d15584c9da0e9ff1ac578922f6b7418d32d4e33dedb86c5b2f5b217a7bdf509ae08439ce154b9afb1c3bc97827cdb422cfb526e8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106be3638140de6962671cb4c4fb9be5365b9e005e6fe93d5eb3f0a0c9933f7d17ff106b6d1beda9d3553b6b5b18b64fc582457c3a546580ec353cb237ff634db30427ad0e0abcdc70fa86fefec30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e8ee0b1e6c1d38bdf02e7889d63d8436b3b1099943baaffcb04327d4f61aa2d615dd9ef557d06a4f422862fb9671f31c60af6e47a85c7d181ac5e5c53f0060a8ad7de71144817c83016dbc4471b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42059a8df0ae63a55856ff49f3d326f744435a9affef378fa7695277970b12437e96d06167874b07e6958487312a1c5369bc716faad6e24624be723740080b172656f7245ea81f9b5e08482d0322;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc47eabdb296955a655b49c72351b19cc769ea4f03d5051a979da3f08eb738ce76ad1ac95000ecd8c48dfe748fa4e89af926194e38ba843909fcd61fc0e6bea779354e3d24db76cd400bcdde0978;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ed3c5591a6797e303fdc8945ca3a030bd372b03e391aeea5ab3d501ee867719735b1599026d80e27c02c315b6291720ee22fce731f0eee38cbff04e49e4b04655ea6094187652abf030ace68ec9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adcb3d939a4b890fdfccb574106e18ce1d4e7631795540f49551b0c8c046dc842dd837ab5742e669867acc3f492037d8180facf8cc26591b7cd1fbd545a442639f2aaddfc783cdcc16b15c1a0f25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141118f81afcba5a1119401863ceeec7c040e1766414fa62920fd5478648652105f3664ed59208a2df6c27f00b44cb6cae19e17c04f850e388b55c5b23b3d33eeb8c104a5bd2979131739f04cbdd1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e22cb10a65ac2e564e19ba69fca7c81d5115586dcb5be44dcfd4b3aeaf7c0366dd26c4a098428976f657506e59260d2dd59699a5f3147d6fd9a45f69bfede4fc12e9bc59cba4cdb1a9ee2f354492;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e3acdd96fd9b0eef89abe25ddd7f83046363737d5445a097f7bf73ce2f6da66b4762ebf6457096d3b145931dbbfa2f2004bc87c4e73603277f0a845a37ac38368ebf6b8dab8d64cc03eca447d33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b03ac01d17109361f34c26d9fac3c72c2429e4cf354deb6b072efc3e89cb935028d28bc3079aafaa26c2016e968b921cd8b232f9abc26d074a5fe206bcdd4af6f03335ff168a67ef0092d1aacf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ccc3fe481760cff1b019ec26e5e21919f01389ee5b6deab0b4d4e20b7f79005bcbc36faab660a8268b348ced11a35c1b0ed4c2c2906d5e3ed35df450d67e02ae543d86d2cebf4d056943070660b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he946665b32da2189e449b829806e2fdf74707098335d0b079df93cc8b275d41ef261530352c96e6b02af5f8e5c570741b410472018ded496e91aada8c8910efb0ca7f88786fa00d888cba1b0b19f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41132f24bef12e023b5cc006240fde73cac28fa9c9484445032e11c6e34604b04470e4c2730f6dfda4c18657a8b0a8e5c2ef58bbe66d926ad21702cf5705ac5288e82378158c8c3fdb8912643f86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6f55b12457d4c992b595026feafd06f4b3b969125f78abfc2cca88ca99d8ee6c553fd1b969060f24ff9c84908ebd14ffa067f5b79e9c69ada0bf7260188fe1ed269e84c53c2431501abd82f6bab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1255fa9f4307481d3ab37ab5e954699184c8a98a086eaf123d9f3fc1db02a3141690fc3ef2ca9098de93541cd297ffe0ee8e5ca182244154d14118b3b24db15fc18dcabaf3c7ebaba16537295bdf0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72e9b45f5ad9b0f7eff70c541d4d51805d98e2c123f2a58241bedbe92f5aca42d3c5aea0d7fc11a8b642f388348bffc088d8699679d5535a2003cc5f122142e7feb725a4a4f4c5e063b6a73e1216;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14badc66b4fbca3a4491390f96a5c82f58e1375922dcc9a1615309ab4d54263c193a04a9b95d7a7f36bac6f2402a1aceaadbbb11cc4b5b912b8a124de1eef0d2e6cf80bcc23c65c3048d003b94d4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f6bda88936ccdd144c2be0f5019bc7cca8d57a2a3f4e3610e9f69bf3719bd8dc8cdcc0f96409ea078f4e56e4231ac4661879479bec460e979c4592d1a73646a640b5123a153cded6638a6381d0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b20afe680a151a9e1d55ffcaa7768e27e787e0712d0a8996ec4f01463c165918a4f8b214c1a64bf2e5c08aa906b32294178b7614406895812b9b02e3976310ea3b3a7ba15186ab480824b5ff9b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3d8cab028e29812098eed3129c280cda34f136eb7a481035b859b22be79aef7f9e5eb1287c614f74581651d32f97ce783e58d33903dfbf3fde0c6e2b821da901f20c95a9749554703f6d9782377;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6f6c091cf0c3663f10bbf8c8bac9ff4d486d67236da3601ac03168dafe7661067d1083392a170e71fbb16f0c72703baa8711a5b95d6de68ea7d5a91917bc186fcf26bd0f59b9c1953c89202d82f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9839af69b7c46f6a5c3933d6ccb14bcc63e90bfa2aaa3b7ed9e37e1b397073f51524c105c489900abe0b8fe6a5404a57554ac6cc5660a357b869db2cd3b859f1b9f256de215b1d3241d87f7816a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ed0ff1f74ebde9b23e4b9424ed863d869ad137aeb02dc0b5e049e34983c1a1c926bd24167270d312f881be6c4944573e63fc514fd18b6eb8170e7901964d7b1d49e5dd7f16217ba1be91ea6d25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h84a8ef3ff29222b44813526aebb030bccd9ea5304da653a962cfbcec08300824890412bac3e7f7cbd8fda326bee6415d2ef7eba6cdad836fde72bd5ff156c9196e16722de3d7bcb5ad9f20fc4e22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77a9fac1a531eead924b054a3f251c40c6571ad723d4aaaa7216d11ad18f21c0e0df5118d16e0cfdcb660ca73d1907c594621ffd8d514d993f23f3baf5bb44ee99adb7ab9e332708e7caa68911a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f15c73b0b38a9e5705b8594ad43ef29d88c82ffc100ae4a91a3416b25460319390a613116e370230956d9c3ff6524fece683aeff35ce0e9740d290c2ad293859f36a5a8a457a6ed8d6ac7712706;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196c9178593508c70cccc469f37dd675ad216f8d4c91c4a3c93779919a849a33d45ad800797cd6f02aba6c023550ad0a3f2e1d2bf9abe9b7f2dce86414a10a2f9e65d1e73144a58834e81a9c2653c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf34c28bbfc9f42d4feaa28673b3bc1317fd3eb8f661109769c8cd49b89960ba1ba98de74d1a35ce1f8731c483abdf6b02c42dbbf0c4736555c571abd85b4ac5c1abca5f01819048dd820db560a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0a245864f8fc005e38044ef490fa7a2bf13d4a4c401eabfa43e723dec6420c5ef42cf73e6b1408e804362dd48d8054427496115de4c6e26500d9bb74726a7c71b33f92e859792b2dde4bb054352;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h38db6526a91a9f323fc558dbdf8078f611948441b16967052d0c4a656fc80264f5b8f8b17067905b1f5ef69709ce01fc302eefb3918464eff8ad928f3fe657b9f65de5eb727230892fac71869d72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1205756f3668768648ec414d75c00119a9b16ce7a2eeb6b2c365a378d4b589c709919a6cae79758bc000100c59ec9a3d3c99c7298890da0f5395e2a14dee9400f1f8d5df6a31849174a97a4c2522a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173c111e84a4d5f09c38587134273f5ba16b39390d2503d08d666e2991e66e657c20b068e100751ab1dd641840c775f68a1797c08a583906fb2ce98057b6be31ed97b4506627a881675a122906e39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24670054da12cba4c01a6dddc25296f7d0d2b3d78ebc9fc2ca46ab6189b62c254c92fa78e454723a4458856cbca72764b792b3d15dd6bc66796c247c12b9ba7f325067c12445557f2ff8df6d0732;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5dafdc2fa63fee8e859ce2aa9957fef1c374b7c9d38cf1e1bcbc4a07a72d5dc609c5e7e58d255a79da848a4421b38827b6a3654a0fe46adc86dc7d76b01a7941158b9e3fcc142f80fd5e85ddb73d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fb11566cc952deede48cf34872a53c2c19e6d4099abc9258471368c3f7e08c078a9d8456b0e111b12bc9ca2d92bcfc844ba8db8de418849ab30376f9fd01c20c2ea33bcdba004230f10def3a420;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b679d1482a9476864a1e2e3ad1aef4dc501dfa87aeb0e72650a2d8329be07fe711d9447cb371c93f969a1f98ec05720327714257d036a8647564d71f1eb78b797b1ffd2e9bf178b3731df60eb462;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h444697c4673a9b5e061559dfe1e024b262ce358c8dea7a104a69cceb06a14f3d1b70a46eccbcf76fbf8f7b5598c4d297e92fefe862661db214c52d647a837047aee458672ec44f6c0c6fc4cf46a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd66c755ba5d93e71fe4ca6e0a5116cc0f8dc5d90024248e2409304845b3d58f61411e2f340cfd1a152562aacf2e67f89979c1369e324429082638090741e4382dcf8925058a40429c8b848cd524;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c3bae51d040fa2a4ad14a952cb33ae0ed41f7e7bd9a5ccf1249e7687678bcda0b1a97df65f6eadcbd62bcf48f3229983ceb50d17a57c46410a9199b9868b86314132b7ee105455f358682060a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17650a6c347d2fe447ad0b1949bb3c73db8bf0c93fe9142f3b16b1e5056e4b79d47f9c1f292f002823a32ceeba4f9e41e32454a0050470c3fc4d3c784d9b0727d8b4166bd61dafa6a1140d7afb911;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1629ea7b2725143b3691ea1af85c620231ed92ad751f0a06cc94401bb499469d4139c1884f1f66eaacfa241b2195a6f3a695b224a5f13e665c8f49e9c1fa38f6fbd5140fd14d5ae1524237bad0c0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0322fbab539353e045ef11548b2476eeaf1c5c194c05a1ff0ab08d0063006a3aab7f7aa33971b462658b8f0940554534b89d081c68a35439dcf5154fd84abbaebb95ee434df65f24f3329a076dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b4b24b75aff7685fc9f0e369cf337637c57ee5837eb6ff8886b9afd190409916e420a08b0eaebf6fa1f9677c216c0ebe5e898dde5ded9bb12611798e92eecca05752ae9220700a09a2de59f2466;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75df7ffb12f9769253a89a0c410a44c76da2e98d783f41e5238101ea5f02f3ba838805881f55b66d40e5cc6b58efc8e91a5824b849e5d0b5dd967ebc889f838baae66951185b4e40a895d0b01df8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5a2bd8de775342cfb78d6fa5e5f75aa7dbc09c4e483a3e50ecaeeda69ac71a59fb2118645b0fd8ef4f68cd208018052570e25b8ad043684ef0c25ea2f9c964089167892e3348eed4c84aaca0299;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfecf7d10b73919cb19e0ef3a784dfd40d1606e420a95cc54089c2f4bf54c634ce4df6242aac6b2a2e1251dee1d6763d782bc744af2554c07f4de593f8c1b6877270dc857abe892f941c14700447;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7bde2a88cf2f8c6eb4a3f86ee886b327767f43ba3ee814ef8eb0f264e9f66609025f5237cafce4c1e584c9368888618b66a600801d7ae3d292b4d49d578c36e1ee1ed6748658f4d590847d4e3c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3352e26a65cc12b3af25cbfaa99652d02020feded084f31de206d681c485c6ea7e821513bc196ab9e3ba03fe82c906758dc9dbd2087cb4dd12cb81aebb0fcb836f8fe506e3863cccc9dffe5e92d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166f9151100bed6264f65a6d832045fa10ce8a3eb107b986f460fdf5970382fe2e238bee552df1fc712c58134930ecd84140ee9a7ba9169d4582483746ed24331a304d454350608b85200a5ee9694;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf285ea597fbcb5bbca0c6ea1177c9160a0f06fcec7e2cde90c0b1c9be71c140905d11e86d6da769ee2a2a7cfb6bd27f952e38a8b084384b94f5bdaffe05a24bb17aa16f0705fe33c05a9d92f4809;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca26ebf8c8bb43e7f5a1ea75aeb45df7107d9edf45a4fd38b26475544a72b62d1dc5efa9d0d6aab210d6d307592c2f7b5650d2083b86d40d424412ab455490900444c095fc01b2cde1725bc0f7a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3571e5b9e66d0e566cf7fa21b831a0ed2257170cbdf6923a9ce92376e35cc892f10dc6eae49378777d85c60bf3897a454cb54729de284781552a7fb6b1ee1fbef1916f875a4653d337f51faf57d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h914a3865a75fd06005b180070e094e9d9dbf5a2ba3d26c283b845b3b4b86d415f1a073e8ff78d9b9fbfe4d8a599fb51969cccd84b10801e6faaf78e589142fe3ed153c768a9947a46f50316d0f03;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb578cd889a24c2b7f1cc4a793cdf28e233903de645a32051ff9fe5455c061c14855ccbf75ac45ccf8f82aeb0822f02e7f5fb05a4b7238bef8ed5364658832e85e2b589ae09d377122408406f999;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fb6f8e385756e36c1a111ad46249505a754176d93bf146589baafa3ce77c6b1c12a6ad35079d04b8771cbbec3c9041b8ab6688902b480533c917ec172426f39a8458f7d63e401e8d41c8ab097f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e5ae969916b715f1c2f1f8e4495023b91879471c042e4662f94f33f73072a0cc102e536ed00708c0948ec40609fdef7552ae5ea2dfac8a1411724b35a501e74694970752e8d1317670124c773b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be786d4d62b65816647167b63aa079eff705c1a656c6c0468fa500a52b71ad60ad6da819238088abc095d968a1b38aefce4706317eba73b059b95a8575a1338f479bd4613018f56f6bfce340d8e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a8e4e06fa2ca5a532f5075b2cc01c39bb9edd9a430a0f3915d1b2d31fffc1b10d787cdcbf477621652ea1cabb744941bb03c28d602f6e9b5f3b8061979e222ef3ceffe58f8478f100eafe2155e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90a4a16d4a62d54e8957d17503274291875edf2396a0c9fa96a529821c12115d0e2390422381f709000e2b6dfb0a1820d8251db868c9b67235b74658ec1192a12a12a58885cb6f40a0c0178c37ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef5382cfc3ebf562c2077c4599112abe8d712d38e7c0454c8aaf48037a490150d19743c721e39ce81655bf477a32fff78df9d8fee12f42fb3a4e9b7eec50359f801f8ae7554527b742876ab8d186;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a16d8299083beea9adf1c0f0a234d9003f64832b697ce2035682aea0dd241dac30cd17ea28f73d5ac322b25fda56775407af0214dd55ef54e19ce37f311d36a6b15b9df064171b400d79564cf167;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdaf61eec035a94ee2888dd2d7589fecbfd604934cd85f88dc22f4bb26b399a104f6b1186234bc9f5a2a2875032e1d92dd1c4fd00cefe38e07edba0100545ab7f41281202a6cb9b58ad731d616f23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197f7d71d692cf023ff5a8e543a5d31ed2f9987bdbac723b376bdb6e8c3f6b3b680633724c591dfd3cb64bc48ba139ef28fa00a0b2c5fa35ebc12fa72e644bbc8e0be3442f605856948f7bacb3093;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132fe675becb9d5c0cdd8a558ed5c388ba6216a812127135f8220137518f0bc7796c4815036915ee5d074202a0a31b76a7dabb277e30e440ae462e5df64d53abe6f069a7a16fba6353de6ba9a5c06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h715003a9ccced2eb653ef669ae72d8385ddcf8bff5e9f75e3e620416fda097007404704bc355f91e12ff7500f1643121989575c78848e9ed983c52425ef20b5f1d24c4613707d30914e4c27786eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196b148c98c8bf0c0cef18e77325eacdbf70084c51040b4083feae8c7af9783f71d4f9b55f5014603c3f7fff7080bb1fe43c84276d9435c1d62ee5d1c23cecc64b816637d80968d21bced1363b10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ed001468f71415c9f4493d3baecc29adb1aa0d9fc9e8cd560c982f2772107dc917d2beab8ce5b536c917364d59b5ba595a5f4aa02afa1381f0b6f91dd6b6bda60bf4235698cb6db7bbac4cde877;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3336ffcb9990781cac13edea976c5638683177d1d8f0369c1107adefb0d126347abb2ea2cba3201e5c063935bd553659da73400364a297936e1261f2e26e9301555354d0369d32a2f72623d8946f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1130356ebb63a659f9d962c9952f71594c98dcce7e5ad34e8d01b7ebec714e564807613b68518ab0631edcdcec2a25c69e4efc0c9cd72a55c3be0a41ecf556766e12b512cb060f8d95af908dccabe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1063ac59eb03ec3f8bb54a1b00f9e216b06fe845243235dcdf22d50cee776cb06562c24c20c35dc0ce678c2cab3cdb51b05beed49aec54cc3974d2e42a7712b1cb806314ac37a6edd99c167301c75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131b515b2d2285a6e1ff4d62faff5a0765fe9fcc34638c3b2ea1417e5c17375d027fee8043ad40c73e1bfb3f67117033ba137d0a6ab0aebdfe5f078a8e938548b0f4e44c0f4d270306db4c64372e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5d16d4cd176b41eb095e74192c2368cdeb8c35e715385b40fd6fe2fe90f00dd6da294a7c4f1d54c30efb3bd6d0cda15a048a2578a8874c00995caa63d1a2af22fcbed5b187851e1b6cba9f316c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c72ebdb272df32a2b6bd0cd6bf31fd557c2bad76fde1a43777dd2049cf38f06a98f32df4632ffe49f7489b42ac8a866031e88eea07c48c9192fbfbd50a5ab9b9f144d6eada3ea718841a7f4db76;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1658968a4dd43b9cfe9e1bc575d3c47dc17ea56277b9a8228a43eb6b8b470626002777b38e87bc6f855fda1de34e31661fb3d7bb0209d7416ab29da124758c9953d5cd2152c6dffb230081eebc972;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57883573d2d7a63bbb6e0fa066dc751bbf53315cefd7f01c037d2657e5df116abbe73713951ccea593b207b3c6cf2ffdfe58a6701a8d2154f74120a10dfc44ce3e1897298266a69dbd0c8fba8e4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h503a98dc251cce52721bb49aed78fc5444fcc417b724b46ce2d3f92bd976d152601a635ed74373208b6009907ed1e15882c7712734739220106a8ec8ef1efa14927d39a0ddf4e0d954b7ef2beb6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1953a677ca1a35f37e9f10ea62c5acd44ce514bf93c4d8054d91d66e805f9bb1345ad2c3d9c7f8609c2bae3766f961ce95d6f4a57583593a0d16fe6e6245d2fdc188b30a8a98898d736b862da6229;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95f89afc4147693533cccf9219e19e4be87e62919fc9bb7b5cab9683d5b67982cb20801f926554e271ae4a2c29018d756dfe2badf12e3830539f88f248662558caf906ac779ce7bf5468d740af24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a502b1a51406da479bfa06dd58b95d19bbbcd5f415910e97161532f98bb4536cacac800e217de4289a41c35e80a3818fd7f5b4d4543fe2262f2acf80885384f7aeaddf3b0cc121f8666882cd97b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19eb34a0654a0069c92a4b93cb9e673b80ba47812aef4739242f6989674416c66577db88ce382dfc8961e7d71bdb998803ecdeaa360a2f05938d013563576bccf3432d730493d0355ecc5da5bffec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he06341e505c8efd958ddcb6c3daac3e12e9e6b601daa3e15ff7275b4a9ea8d20d2b0b4341ab5d3d415a3030468568c11850a392aa8aaa6144a52dd70fb34c397cae5bd7980fdd25f3dcc043c5e42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48e6e8a6c8314218a9d93a54bf6d022a0c238917eccfc9018ff62d38e0a5ba7e7fbfe5b6f26eabdebef342ffa445162caca3777d2096a1a026dd85314de3b1326e5c9bbb4a39c30099b92ffc7a1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1d02cee81e7182c9bff2ed8f8109f8e75eb7d4c0d0a6e331d6c29f5a2248916471b62589657577bd3d8af0bbdb58eef395486fa4745e6bba6079836aeb1a3f760e2a2ad04bfd585adb8034f9311;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16002856618682714cad3bd3913d7df752bc614f40988c59213bc7252eda5421c9d0580ae588cea6b96c8ae5a55527f407669f2614afac0593acbb7b675fe9877755692c9cc45735b303511caf669;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d02a6a8b4d718f32aaff11dd30f47873c23f61d2672b0626aa2985457b7b6768d1a0e5efbd2d55a95b7fd8ce6880a0cc6fa054c2427d6dba657e6a65261f604dd30f7f0d8dc45b8a01911e7363b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f83d26da8190160c3d09b86aec07edffe4b4e492ffea8bc31350b5ba611f4953671912d7155d3c1c20c2e8b2f5b5e70bb30186535375c8fa2df84ae045e5003baca41fe90420cf3f336e55ad70aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd881c201096dd99352a7b654cacb19d58d4ebd270a03c22ed6452c3fbf82e10bc7dec08d5d48f0f479252676c63ad5fc5eee49f6370ebd0a20d1a8ec02a165a53c74ed8a421237a96b716ccdf0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaab7ae5f053412c143a868281cc961f915e79d8439d5cca1867f7640b866aeab663c1647dda9caef1fe69c8cda9a20ea481477fd897487af0f7e55202bb6633283755d907eeb1a32eea1e2600d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e443ed98e322df8e2fbb68d1b362f5d3499ea3eec68425bcd8ec562833da9001f90e43cbfe418dc9edf792595b4851531a4136fddbb2303e6bedd48391ea794ce1b866ec96f948869555c9152c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64d8a7dbce90e5821b5c459e43c8ba7404cda47f9fbd809828dfbceeda197d3659e7b6fbb394de835cd3b6529056d88110dd5e00e12738a4da257e223f8ea145df1755d8c19d432e3229bba1c7e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e3b0c8b2dfff6176a6216d160daefabf7ff728b3bb58430d23e8af7460a9a476b89caa7315eff7f17ac0fe23fb1e024836ac73687da2bade15f72fa56f61d52284af833dca7ef31c7ddebdf71d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3292044ce6f8cffb2324d5e764301ca87208851b2154946db7b43be71a3dbd1221c1488a3b0e52c05b27bf886b4af4629a1b0b6d9c5e35d4ab8d29f085674653b5e1e363ded1be2aba8058b34f5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3052863fb92062f070863f7f3bb2f52efd791a80a4619ce9d04de3113c918d8e3cfa45691e518c0460ae8233d1bd9acd1b077f32b4dece84dcf22641314f15eb2ffb29c51ca7b8d363cd158b041;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e038d18b2766a6c34e329733ab542f352b250c881b794223c2b9b49e93818f96e4991c4cfa1ceb4676bb6f6385dbbdd20b45ad47ec2b82bba10d7d0bea2922442191dba5f54a327dff605c33116;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aba31c93ee9639347ab167dfed10f0e7caba8165bbad5730061bf295401dcb43c1ba82bb5db802bf01d97ad31b58d6e144eaec0d11c56c5ab7cf34a17168e548356c59a9f94857edd5a795286f36;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9c8298f48bf6c9025b759cdc95615afd7e5acc92ee004d5e7b0467ad43cb195aab1579ff56f6b7261da5a9d6688e448e2f55610846588feeb9a579c66e1191b4a6c6805876eea5907a08655d874;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189fdf6378c2d0d95ade77f91a0a3bedb7166334260356eb675dca36e1dc881a859b4d48b91bf4a6580e9cd330d6cd4c632a8d9abf2fe2fc8e85ce271d9e7d82d9bdbfbac58acba9878071803ffa8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he26ad6257f986610f20f342cded9aed4a5d844122d8145074d6e5a55f250b7f15ca2f24576660b7e01fa9899cff80297df2d7d665f14960cbcdbb8ac3dddce110f2c7972d5f103954d640611afee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9f452c029f640251b2a6fd2bd2195340e4e67122aba7ccd53f4e998e89545868745cc32acfa15ac5eed5cd76b1487622f93077d04a1a4c0154c58d24cc4c9ec553a6bec0149d5321bcf75e7947c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc37ea929dec68e23c3840c47114093c09680ef307a8e8dbc7a250a76bba0a0e0c3453df5682d502cab7ba4adf0a0fdcddbe9a47fbe517b3b7052aa63d0790142f5150c23ebd8b88c5dc388cfae1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0cacf3fa75195ce875bdaf43b11352201595122f4620fc6fc571a3766b4f52bd7682cd7a28349025b1224e289698726b6f1776ad20546a8cf4579933b0ce633e816106228e50f6f7ef525a79325;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h282dda7562bb4f5b82b2c93dd484a1bc4574d88d09cb97802c4a69948ee428c97a5a9f3c6b30722899d136529c8c4f92dd85859f6da7cbe61fa111f1615727814d7226b587cce12c7542f515cf0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd14e72cefc9fb4a0d7dbccc2e4338c631be408179480f2bc5c41d736aa75277e3142358812c6cca20f5c28dcb0226ff225da48b818e871d8fb5feb8af9c728fd83a6dcc4ed58e4628346a93982ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d15d3984d914dc0a9445ecf9a4dc4eb0f5e59dbfb44102c58158323013b8a449277c17e3ea701dcdd268502454483ee377d8bd11af094d2d5751051d901527a15ebc5654a0358c626599a2929289;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0f438dc5e95135926c03cf70a9c8a0e89d28feaf9a6f9dd92e25a50302ba1a2c6a132a637ee6f7e95abc35006946a6673d64438c6cb29e27bd2da9be1b028f3bb80b2411202b28cdacdb401176;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7ebc8600b0e0ba6cf91a8bdc72d10f04a58b587c8e26638c376abf8728742210d83557c2052adab9a97c9f165cf174aaa3418f12be92995f32bb13cffe816a12ce4e7a04bd86fc4e5f835c63ece;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a28be3804027de2813c2c407de0c53f7ab057652e7890fd83acfff9dc14a63e16bfb31d3f88b059a797241b5d5f96570817173af0d4ddc2e4985a20b3d571c81b6c7a612688c175782365115dda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9db397f700ee8f90ca292946116eff218f8c92ba39abd3603b13efbaa0c422128f3fa18295ca0fc4c928948eb2effbaeee4877bf2beb1c20451c563b3510bcc4dcc498fd5f2712b57b067b28ce42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169f9de8b1c642e72f22dc8bdfc77cd63e69abab077d02bc5e631e2a1326bd54eaaf038c8612a747b0b3e6622abc213873866bf09b0d7a1074e1c3a7db736f26f6e97826ddf1aeae2ed1aa70587ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5ac02d04ee0c469c7479e02719c1b661d017834faa3d233e5cac332052cab769a8c0c4934c3fd3c1dd52fbf57a203b73b1b282e02e1c6db92cdab938ceee0410ee3c16e61f5c8f3f24c9d70a411;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30a7bc9dbbeae0f751320ae5057bf272e79f0502e66a7bf197d7e3a362b5a710ff8d29e65fb61cff8c0efb0924cb154a193f3e63619622f100b17e77c80fb3be349af4aa77e01e8dfafa73f473;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he68af96b96da88d891e8dea50bb353cb74bbbfdd3f09eb0033e13e0bbbd2ac8c341e8346da7a222e0ee43b26d5020a021aaa0f69776edf06e5c4a297847407fa133cbbe52e4952ec89abc3b2d15e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133d3f3089a25e08e8dd8e2041dba067c71f58b1f7aca58d67253cbc20c72adeccf721a8ebfda51e69203350939001870192e5a109e1e9afa1934c75b918d4fd9faae4aff7fcdc9fbb74fc57e9927;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e5af4ed5b990ba978127ff1f3e265d969c54806f630fa03aebf6e9889d4f68b13c520c91a7b109e475978bc98b2f412d57ccc5b9f89d430c23f893247c8be1a038df8c3b4c1baaa50bd4e73f915;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a91446a999373fa306bb8f53eece3200bdffe5cdfed2554e07bc323f507b8c217475787312ba85258844cf8cdb798e00b5019bdf5c56c603ebfb3f27a347b2cc097f7948f446e6c98236fb55fd1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192c916df330dfd4830ddce12bd9f2b19dee7fa730d0f397590118d60f45495ffb4aa6f824b592e7b2241da63b92706e5eb5b453ed1ccd57e37410780b6c4bac2ee1f488f02e1dd1200925b4df8ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149515b1d841a4865b605cc7e867c3dc150ea51400662e6c6c71b0df89976b5e7eb7e89f653315de8176279ca25911fcbb48acb4a7643af3d740dea4a22cbd879a06566ed7de8b02454d8b2e17ada;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149520c1a72457ae7dec80b12555e5daec3abf41c5c46b68063ea097e54c0855a557a47a62755a767e3f549408ef2ebd0647cdb0566e9c4a87fccbbae7f2b6a12c1ecb7c7171ee73c07cf21b7e5f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff92ae4a0f26d00c361205d07bb9cab7fd42855ba457f1deaeb271d94568028be07e3054e7cc080244a3d57c6956b4425f85e59fe69ed5e73be8300ab2fbebcf248db7cdf0d1e964507402fc0b63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h542840baacb60c421d30f50e136d05be9241af00da69d61410469bc83129e17cbb2c797fff622f0245f05683b007429a6e66600e421dbba77d06e9b88df996d6eef2f226efd00fd3aed4da6e4e6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f180010360d6f42dab42e4548b2a52ad5d31c94a7d564b39dd16b1ea12d4a1fdd4b754de5cac6201b50c34fb8a39f7a41793972a19657c7b28655c8f9a05eae33ee7e50f8b32ee1acf0067b291b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c332cc27178f6ceb855893a5fc1283eb12b078ce19ee9c916c34c54317b4c50e9d9c2eab00063b9c5cd21f04a453133a99163035bcccb9d0f749de1721237f24754b94a1742cc916ce1204d17018;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc644de84fba9f1f039b7acd1d75eae602d74fdd4472e01b578eb90811e71e869a353ef038fcbafb9085ce9e41082f5260af2b5766658bf1b2c643f178a4740831f6d4a476c2eefcda2656848ba47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c63e54afea38c8eadba59ca67d5d2d946831e4f90a7ef84b6762cea238aadc97bfbc3a739a0e08a72b4c4e94896cdd4987dd78d5ce5e9766beed11bd052f67ae68f827fc5d8831747f152c92690e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d50a0c0ee587b7c31291166bccbb7a626fcb1b46cb0a3b85994c829a82bdfcc5caabb7fd5994dfd50eb642fe267c72945e6ca0a82660335d3fa424ea1925f392c7859f7f85adcaa9574c3f5bf559;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he80ef19885339d8bd8c25d17481c8d984075c47a3dbd929ff7501f99eb3e50fe6949377ec4fcb01e9972129d2333eeaad4402c9dad2da8d032d7c56612458c5bc518d0d1af997ff3a17fd97e2d28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8e2b6f4ec0555302523f0b00913d4069436b7f286599253354e5f9787d7bd971aa63c71519599734cbb407b2e6c5ba6aea3bd27874ad525423e0586c9f4b6d97f91c22ce33e1dda13c6ec9b49d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc93c369b786c60771871a6f15cc5f26cf3efe752092fe442aabbaf8296b6ca61c548fe6affbc7051c9d5b70623baca9042173e0fb3ff9024ecf69751ba3c94eadb44a76617173589ad604b59dd8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b193b9aeadc2fef0aaf47c1c7755403f5c7faed8794dc4554da32a1c784e99e3fab76f8d388f0b44477a2f77c72575cd59164e2e2e5781b12124182f0c0fb35426b1b76635ad47fd861a762f12ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2962a98e01a4b80aa05bcd45db2a56a566df80b45aa421da1c9a5442b3229a81ab04760f1f518da2039c6226d35879b781bd42605e2c49503f36b322f84dd03446374cef6d22c5c5db79e45fa17c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1975d4d1859ed3c743bf03e86d383e174edbb479d7775b46c2d7716fb4b07c9be9a0747f6479a53c1735a8382b5e5a52d7c5a1e6782a94f07c01a2559c025702fccd57eee75f8ab088711d09d7bf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158d1c10d873ee65512f54b29765cb7f6908950d11847ea372dea86c50fee594193cb798bce7a8b3171a1a2765073fd1b7ef100bbf208dc580ead8a8bc2fc6167e9adbc7334f882c0c25903ddec3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hefe7323cf7bf19785114a36fc897c253a2a7814b91a51574e9a311eaf7ec287ef07ac8a1e79943128b6502bb16c042e76662a18b657a536cecf8eabb51c03c7859920ca61ca9b1952589a0681c82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f068b5a575bd6957f25c8c66c4e058556fff49ff678edb38feedec11cce4ab0940db51e1ec9a57090b16b7e48d73889c78ee00777b8e141889784ca84c5d0a855207f8a9ca56f5f32fd76f6840e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9304a51c5ee8616066ed06a897370cf8920caf161a35c645a584f861e548631f9419806a5c7842edb42bd18336ba5c54ce4c667f873f7755bfe3cafd7c937a48b5e259fe0e5a6838f67978f1197;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18450db0c4bb2a8d3a6aaa7bd81014cfcab486dd397b5edc2e95744e414d7f721994a7c0f608bc8fbdccb2095941526a0becf47a0a1900fe53e0fc0d70b091c29abb7ce5f7a4bc43409a131d277c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faf68e7eb56edde3e785dcb9bd02946e968239336c3bf981262c7d6f1711610d99a6d077f101d022ecf463a305692031524db323bdf705b62b5cec67b621efa77abcd64b689282b974a5244545d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130622b2c7700ee1e7af99b97f78c38b7f86c8717ed5a892d5e3e51ef67693361cccb1c8959454010e50229142c904991b34e20a0371133466c25139804c5ae0c66f5aa754b53109a775726707a1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b3540b4d9dfcffed1ca26fad8455058cc7c7f3dc0351d0d7790fb773e4e90831a96d415f5d59cfafe366a3a1d1e027dc1989936203e7feb4e4d8aad9e7f5d343be37f1d794dbc584b4ad8189128;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22fbf8c571f20e317b430b539d28686cb39d117e8a1155060547bde609608b962db9aa9e7dc897b4824d9378307407e99ec2ab96789731db8aa9f87f62002e2e11cbce0677f8c6a5b1b4bc9409bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h871d3df9a091273d47e1ce7b5c6fac8e952fbffe17e2fa573a3d69969fd2c4a154e6704fe8bbe80e90d566762fed38ca99b56544863a532994094d279ea341bff5a252713ae76b48dfd977eaae62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he369ebb397437f049d73fefbdfda39ddf03ce758d23122b24d17a91b59f81103e2942b29879445dd1c7a89bcf12606e5592fbbfdb01799c8b0120d139c5b30e9adba63c279d200431f3cfd9a19f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9502b1ce27e0b2fee8645e311a2e9cd1b5bfb4f69fdfe80b2d758ed7cf7cf6a2f20511186c06674a61616928759a70c168ec9c4c04adce3f1d9ccf3c9833612def8d27aac70800a960309d4715b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16196789b8b825650a20789ea26a25c8835e5675af6e7abfc2a510f295ff4b7f5291ab94c1aad6cbba76e6c29133c8f5aacc61dee66e2edb6a6d4b7f2c75ec925b6367fc9f249246393813beb69d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbc3adfd4d0b3be695e14a5b9f7a48dc53e14db1d7afca3541ea9527a0357760408c1dcf0fa548ddccdf6d028e56a3527ee3821e238f3a6a804344e113d62eb1ab150d7318e5e9e7b197a5aae35b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb3cbd314ea85525b1465be5ede3c4dbc035c3556c661301c2541d826417d3abb840b26df99e81c4a7af745be6dd09dae462f64d00de53b62d037c8c5f32f0b15b72727b61e861d35d5ccdd2f38f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8cd8cdf7d05d96959d162185214cc0b42e79edc752259b97225fc4e28bd8f01ec5a4f58020fb66f327ea74a7b73569e8f3441fadcb50368ae7d2c49ad730c429757b82888bc0390c3ee3f8126c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7489e63d392c5404c2df2a87a40e8233913ad5f215a6d2f6a78c9f72490a4ea48d78ba150deed48ad051323bfb377b3a5c16b7da4e78ef1791ab01682b77c697d104aa0c94fc19d489eef9f661c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a710a55d6d25e08873e25e65f4a8d22c852c839f1843964eaae1406c567a809617eb7d9bebc67a85b7e1f36e69ba81abb8ede3a150d8870bfc57b2653642e3adca4a03e5faa25d8e822b05cb456;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcef497caa096cd7ca3aacacdfcf0e6c6c15d75408eab3f39d43068cb1b5b165f1e0be61dca99d0b8f7c915dfd213dd6db435cf2fba95d5b8857c21d9d9a98f7faf929a0b283bb311d7e1dbd46208;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1044515362cac4b1f896c05277308a9c2eea670e4f8d51d87054894a587743fdfbf984cee32c1f2abcda398789da276eb3ce1c36f90f0c2e200a2bd8d448367c2bfde8a830f0cbe789782769951f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152ec5d71e4c6f7e07aa54a767b7cba7082eb37c4b1eb81b693a66a5c16e18f01c983afbe66e5d5c9fe7a8a8b98e1048dc96d46e86d31f43fe0c4b424afad52c77e3294dbae8305a5ddd3226727a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163a85bd42495b16a05ce819569cb8e8dc916891f80988c07972c85d42c849d0734cbc7e02b7a759ffe75e0a896f696daf7fda78302dfc1c8be5d7c8c54aa53ae61396e52d9312cff49db919e0fbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de67b30c905cf4b19e493a6ae13f3d5398a2e2a0c4961b46ff38a03cadc4a3c0379332b52f8496bf73488f6953d922e25c391b94ef3bd62010eb5941d4441a535f664e40e3d8827bfb381e79ce41;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0ed20537e945531fdbd5e368ff7d0a1b31c3a876d7e4ba9b9d9992c8c866d273c8a607ff6260b5ef4b9c034bcb8214f5a98d5aee2810f9d2872e362e7e43d11ec347b584934c96ca569a19d3f1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha79debf3156c980c617d9b2530afe72d5c26824d3de7d0eb7fcfcd357373668d9d177f98083df63fae802827cae53eee781c39513b0e2424a56ddddd22e6582bfda4e501f84011ead560f00b48a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9a4e651f5a39844afa0d9fe26ca2664d0011abe9578340c2b18cd24823e62d365a53777ede55e26cdd2946d97504cad9eb7c0e20202ce46f1cf3372516840e255dc85df0df45ec4b205a6453534;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8db7cbee9a0701d30fcb38ec4d958724a7ba3d01b65a7e1a41ada64dbcb219ec92b7f82fa0d3088fbc8ea6455ea32e60b7aaa5111b6cb2144d8161f2aa1f4b21a16c742b96dc1699ee849c6a8c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e0cd960823b9c302a64fcbb35dfd216e87e5422f3f52c5ce8750c19eda8f4110e671ecdb97c8ccb22151b31add5c0d0a75f7e4a2fe39b1c704e25d9f6c186d5212ae36b1b52a09b172c1fe8d5e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc4bba4a55a0aca52c96e9cecd1da25215cca79a77bfe647163f363b3b0e3d662fe50e811b6f453ebd042ced8b9a2198daa460cb7ae920bfe3425e01552ed23bcbb53e55d299cefdd3bf57229575;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1926a6f27f7927cca8550180f9dfe6f38d86143a942c7c5db5d58c5f8bd9dea8aa5822e3659c8af22292f0df23a0663bcb4e37ae2d5bb13e285ee59fb85c792e7ac984697566146448510da846e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d86d67f9bbc1bb70e97af890848f4b4b90dcc76232effc72b87e333dc97ce229da94345ab47494a9e914bf15a7ba83d99b8edecddbf9e26fd447c069585fb1b4b226809675a8d2dcba687d2cd43f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ba1ab1b73cb0c564461059ae58f2efffdfe8be9cbec564ea573a59e6918d8e0b43bc27db4e6b3e89ee85941dd9598134dbcdaf34eb5042648f1e7ff0beb47a42709e8b3da82012bb85b57511141;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7103c1dc043aac5e2762cfba2f8f6657b33c97ed5160be4f26e04b8e4bfb526e860842736a9ca125700478c8c57d49a6d6e3009c777618dbebc29dd3e0e1024d29213928a39e1fe17557b9db58b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h427c4a1c68d390297cd05e03d4fba9e4b9a5ea0b3c688eee56c8d6a30853d045ddb57888619385e9e8a94a5418966e7f4a8bd47861e66bfc4fe6035f78cad8151b809e817333169b40c2be9a3bc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c103b96ca1db3426013b2463a28391ff755351cf27238d82081add91118e66f5e1ecd3931f84ba0de6522c3f21cb79d178578113d6065ff4d099854201ea0134b40d6d2c0cde6ff909acb6baa99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3325ac4a9ccc514e3dae282f2d9ceee879770f854efed909cf0572f3077fdc48c6718a3a7f492a0711ffdd002c55b6fd0ff4170c2f9131e48e7f591464061fad425c383d5148117f70b33ef2f1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1905b41526306d59f8411b6236cb8add2a4e502b7fadd7dd4f89d65230d24a6218530697a338c791f91f5162995986b9f80c8d2b065c3b59cc9070037166336f9587879a906385e5c0511db2aa1f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d095a56a6024198f0289f3e46c829f3b25f14a5bd0eaa3a6f62931a110675cb797b7e0d0ecfe895fe3e9a13d5d212a485de1378bdae7bd982c3c1882af5d0314a76107b1b82b12845c56d1a966a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb96c4dfcf327fcea70dfce869e36daa3faaec73032b373a09c0c7746d7d624d2081767622a939cc842a1680656813f58d1fd87f641d1cdc3e7e94f6babbfc6d2aff007e51e4c28d4737db1dc13ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bbc8ee061a8e12401ea924011e3124f6780c075d9479e063d519010ab45d1986becb5cbc9cdba3a2af01d2e4f66a1b987226abbd3ffca87b7a3a7676cb1ac9d72b1f9852e481ce12d43e06c82a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52f15d23fa865e81418d612acc4123a8a986e8d7927e6c4a0149cafd03d3d6a8cbdd0a6425cbae48b63f7c992cfc07d3a8a46ff583101267454058005cd166948dfc86997ff271ed7fe7e99aa472;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h156b4ada4833713d765e5b6b7aeb529a9ad1c9c3ff9346f883f938a832ac30db3fe2799b7762df309efed2b10bd170ddcf2b3b04e87e9b3a2afef5de51fbb575b38f93a3b66ada70d5f5536984286;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36387aa47448fd8a640d18d7a9854e93b58983722d96deaa32d2566ec27dee4a5f53fc03b457007a319be55a31355656823a3a2ab8f3b8b98099e0ee83b858065ddd7892291437d227514b23392;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e93dba6325d486f66651f4de4efd1c6e49de8b588cc1189599ed83202dfbe3999f44efe95d49121038ae57ea2c78f09119009354c83c04c14f89070cd91014dc760918fd3dcf07eac3a672aedc3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f1c85756ad2aa2102af7e87512c153427c4295ee922244221d2a8ae9857e6829c9c64c10bdc1ce368690928f7f423226acedab1e832a64f36821741c0d7612a34531e9183ffb9b83c3b5f20c419;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9343d924b37837e0cf0c529841e400225c6a846fe0655c11f31461047027cfd14866f7b814e7a88f94ee7b0a441dcd9b371caa613ad5846fbee65f85d1fc07b3df9c8cb69237f3c34e96559f5b9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54f4a43458ed02f731cea06764394163ddb65fc81d381986ec9cecb6180e179f73f35747ea07fc9f7093cb768fcc0b40ec73be2545d8f84d0b14ffdbfa8fd4f7927b49dd9caad2227803e2370b3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h832e8cce9201c437f141ea430f335cbd3ecb86360c38fa41cd2d3763ddabec0e97568d1e210c9d06b55ddf099870ad4329b145f6dbbf167446e7c480f6d7045c713f101bc7cd6b160aedce7ee2a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b02c442f66b9ed6203271ff70483c264da8defe124f49c1a7fb12a5d83044122ceb0cf0b107d4d89a1b58432ebc2a71c95111982d1bfe761eea40fdf9eb257bbbf4d464fcbbd54879da66cd5aab3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62c2721c70e293baff3d3f49705eab9ea899da09cb5d742c74bc60c59693f41b89ae4e5d46fab8a48fb1e9a1237d83ba8baaf387ba1d3593027f5b99909c6de9d66b5c358c21028e68e3e4112767;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdedb57ab02e72d4e280a9130d43f711b277307e44d07c6fc22ca8bfaead9af368f7ca7900175daf3665b3808e1ac6e24e5890d2ed8c6e2468c1c9461f6d145b3df96f25699517a0d6a16d87b8f9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h174ef0eff342764fba9f0d03fc945b51eb8d1d9bd178d33042e406fdf13477c181dd89e6488e45ca9039450d9451a69e78a4fea8ed903e7ab1ff435af9a74fa8ef3a694fc9270bd2b35cd61bc28aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbb83d9a764cb958f989ff4544b0b83a4339bee96e1d54baed542ce08057a90bc4dd0ad2bef752f7de485c5e720024c3a8dceac4b08b700d6487ad368bb79b615d644fd43aa7158db81c1417b9f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf69d48278232a24af049c92f018670994dca0add9c3713d30ab6cbb1176cad76b9610bb327e511177d04545ba532ec371e30d8379190295021b3ecd03cb854da1294f01e2a027e2ae047f73c61d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173ab5140c545114c9388a99e3999cf18300adcb8da9bec21981d273fe12cf9c241014b53dbb51c654ac7fb635bacdf0102b10a6f838c758a2a441d0352e1da70f4e29cd11c003efcb187cbe5ba56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc0f013a77c63550024da5a4ece3d8b062852328a22570bd3e2bbde7f9d12cc5de4658ebcf073c26f723b825d72574980fc32138c228b05c382b0ca55ac413b3c40eb3d4b571094c8f118f94f858;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7d34e571ef2dc8fe316a2cb144f04109ce904d2acd83f0af13c4f5e703ce4d37428b660c89941f58049fe35104c1767aa23ed85d63dbd1b789778d0f470970036125be71c17f632b2c5f87d5034;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he56aafdd1c5abde3125c421145a8db56857a3f3f5469cfad7d96b5a72094721dd038da36ef847e7f6d5222b694d2d7e555ee53aa3230d958922f31ca1c8857937a3fecb4088f1fbc5ec1006a0ec0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b1a4fc52e29d56246818ba09b932ea5cd6ed28e1f580531c7d9a059e7bb59bb4d94f765b6fdd8641041ce2bae956f351e9f5d55981f4de249416a8715f0812d69bab1dc52c9ea913043f0e11e8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b6fcd2d4687f64ddda7d5293ed6ff2461b7845a39aaf36f77b7cc81abe0255300c492a9b82c6cea7d628079d9be448fbab6572474390a7c4ee1546931d4b9abc5b3896c601d59b535cb1be40d42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha77d1e2af133ec81cbbd80c996bc0429cd4f3d8f8bac946d51afc4954a149e7eb6a86536d4c8058b27ba5b55494bb9d4c68131c7036b763434d92ec004fe578dc59e84d94b44fb607f93bf8817c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49393ff91e5dc7acaa8c2f0337a6b29a39ff886daafc60a2268261caae26e91f39c9cfe9f1c3c02611d0ca255e8d9edd96211a4e80ca74943b72981ad8761afe74c4ba78b72a7525ce98fb5bc400;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123755abff6c6425509bc37bfcc21d6bc6667e0719a7e68d588c0b803b55b8c8976b05b4ef84d2fc562dd02585a0f0d11603fab7898ab079190459bad298beb0c71cdf501b1baaddf89e9e3962a7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4732230734a4fe3c2830641c1f30183702e859fa287125dbeaedd647f512458d1fce8024e59b712fd6269a81f1c18bd540c28af0c40868f023b7c994d689f4efe1eddf6771ef6de4dff49fb0f0be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6011d3c516d42f78c2ef177400a7b9eb4fd1bf4e49ec6d556b0cd862ba7108e91add60ee6f53e2a71a03271c05b7a84ff0b663b4bf32025d4d75d60be0f6536a6e113bb0ad7e599b2dcc92d9726;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1480a0656cc6c0a8c246eacaadd0f85a67dbade0696d1b939b2542ab3de49da6533aa181c9325193a443fa70382730c806acbefdd8170b8cb68cf315844308f82f86f12563aee0701738b247446cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fda9a47ffc932f852ddf6bdd8309471876c3a5ed43913307d8db7dc63ff5385957b47650c82e28b09837204df8ee1e08b3a51e0b788821faa319fb3b6ec5f66ce4c244de4922243414d61bc5619;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h624893554f6144e7ae52d3cb98628d5c36981a6aefe338f85915fe219f628dc63b2a498acd7f82c8782e809d0fcffbdd06525d079d3453540c5d18b096727a948756ce883ceb47f9bab9149c0dcf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7642d26edacc15b2393506ce3f1dc29be3e5884f27aa74730cb2dc574440c2a9e8de6a01a6c6548ed24c961058ca2aa0db32d410293048df43277be41fcabca7d283f2cbddb2521f778dd1797ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67a2d57af12b9da9268dd6212227db0cf60e87e71387ae11f077e87b6892b371fb9f45d758e0921c304f278dbf0009c01c06a592a7cb71adc7ac42b63d330ca7b09810453ac8101fea889327ca64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55111bdcc879036cdd84799248a25f0d9fd8973d7cc8f646cf4a5f3626cf2933cb001ae8f662a7723ae57fe2ff299492e39245885e0019cbbd606e330545d864b32c4c4d60c97709688681630d30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h505305b2da072a05bcb98ff8c8e4fc8fea867175e5bb8d1f399bdb5115f4017f9d1d7511ce94f074a1af8a8bb27f63f0eacbefe3db37d95e49813e4de361df2a46bb90c2a6551879c50b4563f41d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c8ef2a40c8829da37d35898098f9fabd2d5db7441c6d6af2e6fefefe103badbbd12923da892e37193ae359dd4cee31c7f3a595abbef68ae04df2dbd5070d812d56e8095a2497ad2e5d12db53736;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8af8330d2be4a3542409aa6df8e8e97852b9318ff2f31998e87685b5c64c2aee22026fe7d04465268ec8f5bd9d73758a724c900e785f985288bdf83bb4bc2f3d824f584ae57e9371cb75dea89acb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ca5687e3456c3d42ef8165c9ab0a65d4fbb6547d72f252e1ee8c290e9b5cd7653b4c631b395fd0373ef37d9d0a9a56984ac6de26c60a82096d41ec168cf99f9e2554dcdeef06aaa011f418b372d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8c1b233f189f0f627733a19cc649d760642fb1338b743be965e42457576061ce2265e231bb08c3edee2fc69fa21818d1c76605685736ff266bcf4e2d30544e112030d079a9c2476338ec6089cb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31685dd5103468f3186a9dd50b7ba77d5d01c369b0cf9a4ffe0390c0c93762edbbe43f71809f55549eaa0b013af4350f62e67f0d4a395c56141aec6f05c4bcf091cb31545abee0cfe3cdc2dd9148;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0ea39e7415417c9d585b84d71916853ed9219d7fd9a93f5b908de8853deb996d12e87f71ab75406b1517f6394760b667a5d47c33236348720b7b8d37f95012f269aa1057331c97cdf9012aaedc0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80dd0d1451536e4aec498e60bb73eeb23b708ec43b1767309bf29bf18bccb377395123ccdd64b72f6b81fe98be83e2ed313b473df6fb8d1467e0958399a31822f5f1c581c3fb4166553b554433ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h156715ff69498cdaee5b3bff851c35fcf9b7df99685bfbfb1eb8a8c76c3f69ab955cc8372212efca75d338e24fff60c3c9fe12b0d0cd7b1b9ffdaf4da8c42fe90f0757542aa918bc30c9dfa9d413a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153319ddea4cd7a69d78361d4b807743d9bf88430bbd563f71c8a5d3bb37729029adba9bf1c7119b2fcb1e1ef4f2152670ee598b9a3254f1760d09d00265a4ee7559a723497bdea039b81cccdf39d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81a7ccefed9c7704d9904262b0cf79c2995238fb17bc4680edaab524fead41728ccedda3ff70d5763cbf5ab3573a4a8252ae52382937eac882baa51966dca4b34c1fb75cd8f67a042c8f792d7537;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc8bdba0ef2798a0e7971d47e14df62c06e9209f2c903a088fa351602035cf104edc9634e6a55e1df6141bab2530dd16e03aa4ee77a7ad24e102d5d1f523ce9da291b3f989b2aacba391afe5936d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb24d32de85802f2738a57cdcdaacc3db2bf7817f2e8731f5a36da59d129ccc385a9b840b28376f5acc96d078edf461393947fba8a85297eaefd0015ab722264e3da88c4a656170a3ef5c2857816;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1390de9415714aed92ee7fffd6cec1fec589783a86909e9e0b921fd8c9b40835e993847289cd93c669c421d22b11a2abb408305e6691c88c86912de50be27ab3dad8ed7aa685f40acdbf2cdca412f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a9dfe77253d501b5bbd2e295a7e1b189a70d381c31cf7fe518f9a0af39d95001a8c867cc755ff021cc206c72c26c3fd8111fb9d13488f44fdbcbe97df2c793d5ccc5fa824cf3284bae812a7b2f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155af9366cc298f4748c8f65a2384327ce87cb646e30770d522548f73b21bc16471c44f9d0c231515a2815ead469029666c84e208e0fda4f7889783b12a41bb2415b4029791d82ed4d7711186f914;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd7462edf50fb202b56e93bf497d3b27c719395ad539466ccda84561467da197a44eff14484dc9c95c8d54164e61278111d3a91bceed54d21da2472afb1dd94bbd7f21a27c82b7d1333d277696ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1082c690c8169ea097d591d9010512a6ad19d1cca9d3efdde02822c65a43bf2e642c01ee547a4a5c3437011a1604b294eab3d7c9648778cca47859af4054f3722b7b0faa72297ae31391b2a898e3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a731fee95eebf455dabb62e918be6c0b76acf9cb79f81a366e232a86221820a918bb24f298ef269694c8f2bdb444b81a75ce476bd10a8cfaa896cf94d73484bd3cb0e1c2e0743657ce625715b513;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdef875c836bd869711d6e52539eaf308d5d8d1b62fcfe790c252c0a59aae8642376eff3a963e4d1c3e89ec68eb875657ed3f1967aa6c68d23b97700400d94d008f033b9d71d35a9aad68a58e5135;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a84933f77b96c02185e01cf1cf7237a2a8239c72b0e0298c60542f6c688d164aff1b81fd9efc1da9b5ae4b46e21e58e2c66e65d9284ec7c6c7a1fe59592a92fbd48a2a7b4c9f2d21687e88b1f83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acbd9996a97f602efd28e98d3819e5b523521247a420e18810a109f5b5a2e777f10baa97413df80e97644cd881af7375b75e979e567a5c17439001e64a08c321faa3b5ced763091e013162866937;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b74e02c79c5210e4f562bb60e667f603908c322c67c6e0e1776a6939e2ab3f5fe728982c8e27cdde877648227eacffd4c1b4b71274c04538aba818a6ece6881e831a4da1ff09b0f97576f9caa33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f8bb20a0e9da9e792c7e73f5f11d8c10327031eba3e6e2ea7226875243813e9b3d499f84c167149425c74198f62a34a58f7eccaef958bba672d47e42d1d357635af211f274901163dced352e8ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4e827a04ec1e49b4a8ab5cf01f7c2f173711bc4d667ff248b00097f784d5994ae95896edf36834dcaa227b5fee6d71b2136970dad195663e28665b94c945702dcb4daff2ddfcd08c520bb8b1e46;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1dff6a7367973b5749e8679772bd91d423d048fbbe31f7f85582e26e8e5d953941bc3de64c299e8651df92a419c4c0ee349d780d53ff894d2d4a5dc3548a8da3ddee3dfe4b2907c2d823b40bc2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12adb95d30117c10225c755b9ba2702f3ccf364b69806db27d799eff50fbf491a568ab94ef80442f83b2ed61667712058a41aba8fab45be7e99a0f36d49688fafef9320d9b97a41c5b8a5f4d0a764;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8851718a1ff9fbb64147711df6829ab9b382d9171b74d9b04bfe69c8f648bff23faed5745125a3df872fe71e398e1fa81b3eb1613f82d6b3293d7f93438c8ed3c2f12cb596ecee7eda5dd032a0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4be837d7cfb31feb05b7d89f0f8dd8456f6ca73356a9d41e5c0155f73ba39dadfd76c2e615d26e1b7e39ebc0e20e5386590193d088ec47e9500a95bc90240c0c7116c946397c969934b00176fa40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d615b429dad5452cce6a33cae136ab57609ba0aca55e9d8436d4fe4d1c601a49435b2bed8a5542763cbf943818a9aef872fd13075ab2d58056551d7e848363f9c870ddd0599b464bdc03ffb45f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f56e512b323ebdcd3cca2d15be336ee4f4aedf8494ed34d2526395895d498459a9594d2adf05fa7da08bd43bc86620fc9729bbb6736cc0ea396b551c1dc9893189bd265ad0eb14b86a5b5847544;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4165e79e2cd0473012b8ab4067dead100495bfbb709d5309bbcb8e86f1a6452f4701a0b28e9fba445ecd70781413f3d51bf33f847c2e3507ec34e74a8f0024d61b253d7777150e408559b4ba2d98;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104a41171c03647692484edf41a62b26a2a59f58d6e3c496436479ebf63dc0937ac194585a852b0ad68a970399c003083c1244fc4f612d7fe10234c8c494af910982febe5b2260238252f33f832f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd87dd3f4af66f243298284001747606c87ba2228288efaad722d8086a1e8adee57347b008f5c1be863de19b55624940ed97b23821c53cc52fa1126177ea4c36ede1f231173276e2698406064664d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd036e2c007e95ecf5789729c6943ed4ee2671b5a7dc99fdba316521c3210ce0a3e8e847a5297a3d50dcbf687a1efe44af96397db21d04c5690ff06256e14cd960d2bd00ce28dc96e0fd04b8457ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3c5ec7061e4e9712a38c05e7604b4474c4d61197fc9e0008cc2bed11c4f0b9c515121b64bd30c1829c734bcc3e3c777b6dd364690badb801211177758d4a3de712a5fddfa867fbc24ad2e1e1331;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6fe6e2545b38e469821abba0dedb9de36b953004205ba3018d9048a811b112aa4ab15aac62a7a2d47fe874c2182606a051cca82dea3824860dce7206feabd176b87852641bb58a913a597b3416;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53e1531d5a344bd1815107b6a3756f787a24884761ea9300f573d1bc5f04e717142b84b36d5d2c4658be5dec35eef8b000510f8746fe037d2b868b455fb5054bc119273864a45dba9165ca81777a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1705d60286b7f735cdce57037c32a612187ca2e9eb8f2fe4da115b7aeb64faefb66a06f0c0b60470d96cea90ba50475cb8b8401e61a17181aaa00f2e6c59889b64f569022257c07c3f8218479cd48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125afb9d3ad70d196318c0de2e5018b0b1190d80c8d252f6c325cf0ad5ba9d632929f184af9843d32c275c503c0a8393a822122c86ab040cc1f3be588397be5c8097f646b64d4fbb84bf59b03c702;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd12a55db9fc98b0fe183fc979c32fc3648a252cbdba235bfff2434d66270d4196ec1f86a0f0e0660fe5d6622909c5b108a1ef0892c71f77a2b737b4d25f854afd7efdafbcb5147127dd27ff0f7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaac895b19e8b71d3b42076cb67457848ff6fc25e481330c448783f9b0ce68ec480a93b049a494136cc37a33d53185bb1de7755ba8256713d0cf425eb31015fb55a4af09677dff56c6c70373b181;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e17c4bdd65eeb9a78f052f2dcf4ad4b340338d6ff06a125d225af7018bfa8483d9199ce435eca42da3608c372de60902b769ef5301989b0aedfb3c07c53ad56f05f83bee8ce9e8aec241d9f8e814;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67de38cf0716031095453bc2a3c57ceafbb549e7eea8a9871adb01807bc9075f01131e00392c153cac9ca46036c00cd9fa418f64fa2004025748c5b8015444762fb37ccdb9cfd4d5e5b1b637b211;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd2059f659cd0138edf15d2a34ef732ecc65647049c5d6a4712c6ac71236ecd7032787b91bd30e236cc640099f0c3a2cc18db5da2d2a001427809ef8106dbf4ea110f2c14a993afcd321ecfe1a21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c62ef8898463a5037f0937149af9290a2eae0c37c11f16b342d583ce61834b0898362a9765777ad32292668a079cf322d22db44151014b0d13e2cda3abd0bbe9dd3a3f8821a081ba80d5351177f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aeb4a200f9a86ddb6c9b1327c0ff07904f7af847b694e5d622292f47842683023845b8e3f8d3963591090a8c207ff459f9875ba2a0ad2a8e1fb51a195aabfdc28a06c210e3ec4e63405f2ab6de37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcb9fb249343effce13e39b0549e602aae1374d035fe7ce5c263caa3c7428bf301bab5b1d3f025deaa27917be9c6881aba353dbf1ea147a928407aa9102f15b736bca570254c557962e571b9096;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9c9a6a053f5d8083fdb08fefd8eaa8c3c92097287fa8102465bc52dc637ab06660c98b1df3d61da7f35060a91c6eda948f3e5b3c2161fee18585db05dbb86548b3a8836b7aeaccc72e7a1d677b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf31126a0ac9d3b5ced2cb4d0f886d2038be8742391299a5ea99b0780dfa4a2ed13def337ff89064bf5acc4e8a24405eb2516d13f660a789afbc220a71b118547f2b6feada9fdcae2a00570e6386d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7ec3f37f3977bcfc729d70afd988244e7e2f8d7d818d55ef7ab53f084495c0bb910169f353b16bebc8d7b6ef015d9b90784ea4ff2e115b32c2a8a796aa10b09dc805894bbd5b3f84fc018885a62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe37aaef50f07b6cb3b02b16090391699e109d21f39fd3293008d90f700241757cd3e73a8650dc9aa2a04c5c373e5928473884f42e059e1ca3efce68771408b288737135d542a25e144f7b6eb7ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70cf11fcb3a82692f1484a393f3dee48308f8398e5615d170b5f9b5201a542c5b39b7265f69dc374b328ffcbbccfa9e7e061246096bfafd703f8cd1ddd23ee5ea81a7b67f5d8f926d619341fa5e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1418115dad52e34ad885783c0b315746b081e245e8aa58fdf9333ee14b89f8a303bbcef2bf0c2a2128b10c92eff8a4d7a3453b6642fb81e351cf66c8f4693d8b16add5afd94efe08f91f4260e53a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1026137becb364f87aeb9afb472a41021fb97ecc30f822d1a70d988de2b1bad601eb0ebe1aff756c51e38b093cb5f2cf99234084fc74adb6394edc9f23337024748bf36777f1880e6d1de4263c9e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a5b0339ee713e9936a43b4d94f9a948991d205d78d6e0cd58649fb214d13a47c80493974b278692456669319655dfc665856a3b5924c9bb5ef462fd70993584b28ed18618fc2a1ac9bd5ff15f02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bfb01d5f710bf71a8b731664f0a1d0534423ab4dd2dacaa91c28faef7b7c0eca50bc7282fe829abb9e7a4076a96bd3784dc8263aecc7b01b1dd1d9263f2e0bcf840f74c11eb10353d0ad17f8cc9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cc660e423bf469c8f8ea3d3e8ff8ee013886d9b4de1d9bb478fa576f1305f85217cee56a120b2508b176b07d07ae104711a115d58f876a5ae48bb28406c527123eeb377f86d34d834f67189f1ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124cc82ecd136448471751a81e9e7f62f3634e4feb8b06d9cfbb7e273f7f03f6bed8f953480370d727cb427028f19710539e3f162023c0497c255f59b65c85b490948bee84cacecdeca55ddc0ad25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b80cdf6915f6b59531a83e57d9b450a1d41e3d89184526a95cfd382d6f82ccfa9f347f84380f6f41558a03f3ec8abd23c28b242d4177efaaa05a59d004512c9dc4c6d896061efe2e93504bdc1eed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f2215687bfdca5d434213b4d4c0aa19f32242ea04410bc275bb3f29d44f169b4c3f86a27bbb4709aef3a9e165a377f8f94880d72154fb1d5339c6ac50f8687d55870f94b574e92249e54b33fb4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ee5702455ffc3a9d5f42e9e200a3baaee2e84f0b5ed0045cdabd71dbc92f345f13d633bdefda2980e5e53798f80656bcb75f369b4f6d2c308b301a6eb91e8648d57df45cddfc182a56460282482;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbf5fba5fa688db28e4443e2dfd6bd57f4c1fd31f6e8af85d35c7777ba64b75875f3187ab626e465156c054de705886ae4001a3ccbb6ba70a261e66a54d863ed4ea7f2498682c5a9743356d6b2b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5e3c6e8d1b3b3ef8877c6969ce0aabaafe8839da6ce24a698f03ecdc681cf371b42335165c0c07425fd92334abb8c7afd3a0358eeee513f2dd85042069a0d83bdc961526ffb258775ee5ebe1e11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1295f0c57b3bde897710f77f66493456e3ce9e8ff2e2675409396f4d8dc909015bddd72a25d4d31612265ce851c782f1f540e6aec167d5861e90fa457b2e60bbdf0d650b4a83a080fb0996ac80609;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ec4fc6d37bf2aa663eb4adb5487c008312268f2c1d408ed2188a7260351b558775f43bb79ec8dc05bf10a5589a251ec3699c350039d7f8081ce771d2c34bd4ae0f466e8e4e16932860f781c5497;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e448848606dbe132ae5de00caf9e4dc7a37644c8df98873409675a8e5e48ccd0b9b20970ca559b714354c79135b9c7d28f7a7f232e0ad894a7e20711995c386b0d8d0dd7cdd963e7927bd0efd11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95684a85193c24b3ba61e8a5e90f951cfaa58056d0b10a0ff766b75c5762a60a4ee9c2f42d26a0f4fd8f83e8afdffff8be7feb863525cfe1a597c552848db255de05a5be196a2c1d19c17c4fa2d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e98a03eaf1c83514c68f31ffb981fe32d2c3396c6fdd554495e496a0cce50cd6c299699a559dc96a262e84379f73829d0692081bab7cc25d3610df0f392c2539804160b54fbb5500c1d33d7f770;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd8d9117ecffaf18cb6d03b7d7cd8d478f2a229b0aa2bf7dc437091962648698e08c0bd0647159115509d7079b2894d52b212ab67a03b0662d4f2b39505a89fe337ecb417eec973198b001331134;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a46f8e8e6233593783bce74a967c1dcf87ef86936ba8f13866414472903910a1fbccf3977671e28639b73d0e5d2c8cc1f75a285349fea2d65d1ce6aa5458762830398c5326aef736915ca402bc7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h250d1cb89b9d638a8d131a9bf752b662ec98741e58c8199d1e8e0492d9ca638e5d822aa98e83a4120f61c3ab0844c6e34113754304dab8b312afad0193965936b075e8cbd2e18ee0408c43ffa458;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186a4ab26c330d2a39aab93d2c61cadf6ab076b928b02165e5e91627ebfcbaeb306f18c4af3468b08cdbf5864cb012df1c7fdea5230b23252c268ef67eb329211e0593be4e259b168232a6bdead6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c752abd8ec0b2f625a00595f40c1aa1845a6eb54a8dbfc01aa22d1baf85657c8eab678079571d183532ceb5aa22c56c9d81a55be309ecf82ae66018b9e0b3f611b6fb6c220f752dd225c4c81ff5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ade3c21b4ef18c50f25ee434f8d45124a0e0d965b266fdb50122684d42b59783fd686d6d7d62e6830dab0be49b4d7c85cc45b18f8c047c697f2ee1eaa609b2b5e31d2871156021d17b28b5110d4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195f23e087f5c55d148f22d42c07a35cc9abe8fc93f68c554ba26aee09b771623e6816d4f6d4a01dce60b20575c5bfb31ef71947f5729ec8548b00f6ae9dd76e0fc617d6325e6e8a6c7015d7e9a3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1971fe55d24f8451b8f6cd698b1e45b00af6dd75fb8f6c84be719a9c60006c88e5dfd470301da00f5aede198ae36f1fb8d8bfb23b28fa89f73c3d20d3e3b728baa9a14f03813908860d2a73e6ad90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d71974789a8212347acb3b6c3b9834b94c8e053e44aef986a47228446ae2115500bf3a607eb42398564cc529016b6079d00d805b03ac233869acb5cc1e37e8c915aeeda4537ccf0f4b15b017e639;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77b36f05bd73a4a88cd016e6ea3810d3715163d5553d6b6eecf15ee599be75d1f56d0392e8e14979cd38e97555ba8534c5c67e95fa6b799068e838d1d45d2d2b04995648b5762dc46faaea4ab25f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1016591ed4e9570833e3dcdbb2da45d25fce46cb2fcee4276d088cb771a00f6dd47327bae8653792057e8b97498aab74a4290fc5769d4af307cb13bf9a83a5edf88bfde3d9dfccbd0bdfa2aeaf6f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h147a0438b1389cee30ae686b539de5c2c8e0c8f43de5af20cd5048d9201fc8bddba823850e9822639d5ce4f8d876e80a4f470cb08abad0309cd990ef600d28928283658fcf97683ec1bb345f71dce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5ad786a725bd11b208a3b52ab1ab97bea2dc94e882a0ee3d4d69a36d39559cf3962ef2edec68f0774338a00a452789e23e07c1eeae3da1abf89b4126c8dc748217b91b329eb531529b0bcca8e19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128f6150c643d36f56660b928c81b8b98d247542a7d01642c14643e7e985ac4e90bb9da128d7eae80c1359289908082e3250ccd5055f89edbde7eb5371c9b692877f1886fa43312049c41b2bb3d58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e61d52db0fa10153a2ee9f1431e4ddb5d56d933a25f4680b679ce3ee35ab5a976ec07e7658f2af63fa15f7a3212099619d3296839b8ca946d60b62b9c8f1886c76796d3f32c0485af668526870cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148cdba573468b7e189a75f82728f04171b0b3c8068fca632f047b2dadcdc909ce2deafc45f8f83066eb378acf914a45fd989299da395e9aa0a72e3958b93f6c11c61554a3739f8e2a0e20882b211;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2b2b447f316dbcd76e705c9824b0598ca80b843d4d6eca30a883aca522a4f11cf6011dedb44b2fa2f5316362dae60a883e7d4a089a204eab78b1233cc5179854e9fd6d97e3c1c2b782beb5ba1ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136ebb0c731e1936cbff9e402a71be7ff03efb3ec47c9d46eefc8579f9c5087ff4e41ed355142308c95cb90e80b29699d7b4115f11485d1c35345c3c6e764abcd196aa65142d89942f230ea99360d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b1af1c226b6bc2b1fdeb11a1b4daf0afb614a09f2b84fad424097321472b01fd2549f89fb704f498ef056ae4bf172b4f24fb84de2a0d121d4022e53ace12b338d248dfd4be903dc477bee481b3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h890828fbaee162c2477303754bc89ba8a59f24e60d4a7da8f2afc8d2a793856ff8b925942b0baeef0728608546152e45bd2d56debece46491d680de4a417fa9a773b690949e67603fb1998fe672f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcafc248afd36d79c0a4427c9917f1273ee1e7b0bb3f5af15aad4ce6b8111bcb5bfbe24faee64360c43af41631395d19953404685c3dcf749c90c4a9bdd877a857d6dcc332bcf43df195862476334;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e2ea4344a08dc2fa633f8369f04c796ad9b9f376a9f51fb74ffe098aa8bc9b8011e2a0ebf507cd7d49789cb0817e5e06be9d132341ba5edae44c4b6126e6b7f8dcb90dca1be0faaacbd6a966612;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab09b67db47c3255d64ccbd5cfeb5b1c87d9f7d986aa8a6efbd582e11e6b475d6d408647d7d7549bbf2867c0e2faa420a47d3c6c094350806928e041a59ca6960f0b998a01bab05fa180a5071739;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4252e789787815b2f930056bca7e4eba5b5f11124c1f6c7076cf7da3deee9ba2a4850b99628a7300ecdd3cd7e62adad7653c0629b5fdcc51420dc368719e9b6e4187c656858cebae3c646d0d5cce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd65361ee3dd3fb11507ed2721b9e393c6e644b6db9ff31fb9b19db7a1725130b51073d58ce966d1c474d8afbbc3a304572ac8b48334f7c7718b8cf9a99a368f01796fe65a9433caca7c993555cdf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2b5725e0e74606e159f2a27bcbab619cdfe1613df33a07915b14c420e287887f3db0ee2318d770a822168d1ed4120d8199e75334914bb78f8bed95f7229c67eab2b623f938602293f18ecb5949;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a67043d50ec629f2f4a3911d0fafea29f0ea42ae6609b35f3acb5154b8037371f4994d9e0f569f239736324031aad734310dc4ae45e6c8025fe2a1c3e04ac3d7152f9de7073aa2575743a15efb33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h276bffc511363e6e7898b3d908dabd41a3979f554776c747a232cc08fe5c39c50e1485f1b5884da3c5fb548eb7cf9b356a344d906c47e39949a917b2772e1fa39eb4f93a82f12db56a038645883f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h848480db1bceb7b1e81a3ef0636c224cad3a333e156dd2e1e739df9792f1c7b4d461ad2ef141d1378a912d41d6f5d414e39e08efbad108588da40a5e80fbcefc400c3b13224ac13dcd1762ab8d16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142dee15aed657470894fe120cbd5086ae213ad25a91a7d769fd0d97aa18ae9bf24b78e8d8c73e505977e278096f94edb013f6247be27e663028cdbf20c5a7e875c3d1edfbc616932aae2e797dec1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha71551a5bb2102f89c8bb576b07240c78e92e86acee016a725e4caa3d2c413f288d893a6f680faf42e604eb800fa2046037d1ee621080d15fb1519cb651b7fbabfff55aa4828aedae8b38202df14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198cdaef9ec69474667eb6399fcb135124a61d482bf2c0c8a9aa06ce3b2aae62053cf51f820c62d68de1fe0466d3264229830a3d8f8d90f6d6a77f15b06c55188685b9de494bb4dc28238b4663603;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90506ed3ec35139befc23d3214571774406937b6c323c6347547b091c55a8bd76559280ad6c023d1a106d08c946e95d08f772ff5d1be9a27c11a871cb81352e2525b4c33e7512f2321c2c5d3abbf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0cf363fd34d07f1e7266b2d248d0fc5d699056ba679e2a667a1ec1f6a7ca05aa0f5b2eb63ac25a0b743736b2b246541866c6d6825b5bdca5b2f1cb89d499aecf17285321814b9bfa67a17cf2560;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f6c0e5810629fe42110154fe98a185a3942bf3537f604510d2350ab75a646c02ad3f2fdf2487ce931538aa91b7d6480387d134d6dd0c9b5c56995b8a3df14d861b55d4e36b2c3838314fca8bee3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf629f63812023d223aa125a5d4f23bdc7adb7e1fd234e7ade181a92461fd60aae870cecc0a027980c749f7afc2b26ebf892a1d449a7b9bcb4cb789a917af7703f5320ecd4842d0e84be2b1d58784;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcbcfc684a2ebb14da0c14c180f105987a9cc425fda1a7c4bb70876ddb3d4740347bec36a766c41eb2682e03fd2ea04447f54644ad0ce8e1145b432422332984d770177802cb98b8011f822cf4c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1874d643f8f134c4a6c0c4446888f18a02057a152b8b024867efcdaeef5dea5e9ca51b0a1f22a156a72b0cd424faddc3a03fc25f16f0fb47431e790903819e5f37169d897778ae9d7bacbd4e92b26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haeefbc3edaec619384e8053d658d6612b3f0970899259e4205dc9c94f467509b784fc4f58e3f2670a64fe6b4edba462617db59dfcd03a363a5cfd0ffcf20317b5e9e4663bccb5e3ed16af6ed786e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54bc452876e3b993a270771539a0206e70f8bef35e5e8fc501895ad971834a141d4d9e68dbd795ed9173c1b19808680f219b49e3414a52a88b814222a9c13e0e777a369d200d757d628a7f18d496;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5d349be1971e2a145261baa862070b14f724f2cdbc4513cf423d5b3ee21aba450689d3a60c0537522d6941254789728d6ed1480cec015478d024d2b76a705567e880408eee5c6e98cf307a5e55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h822bebb9bf02bb28e972c964b1557375a08adc901393d72d34ce23fb7d6d8522862ae1c3d443f99fc55a917a0786bf6375c4d731e665ad3d6e6baf7b43f192a069c6531a524927cbd2c0861cb4eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19742fd8dcd1563aa2fa103ec2df3939f0c55af9c25c9be9e23e859b8ccbd0e8666b28b28983a05e1c913c5098628fbed0e75925451a443d2a41151c0104f2fff9a71334ebd9d1228d83dc35c56da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a10b8686cd99b16d023d0a7cab65f0a59aadab130e1346be9e1932fe3ec52243a71e08d92796f9d04fee9cd15551480879e9189fa1f4488c4d0b0f5c4ba2b56c2bc1537c775f0e63c0be253d7af5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf6c621babf366da7d9d4fbbf79537dde84f22c3b017a4d7b029ba442524f0eb2001ec9591973d4b6d83764182a424847429b447e7704449da7b813b495f728d00d82018ac576da8894702e0949e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139f080369d1d9fb749eb08a2405178c795f0b7ebdc6b7193720238740d203bcecacf860a2cc26a68c715f85d644e46d83cdd638c1a7de0bf0ca66c08a86b294ed3bbdbf6fc020a1b7223a5d4b32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183e4027c270d72aa9c00d6b223760eccf1e87baa7d71ad5f65b5fe291fc0736409808ef383e0ff2d32493b1c1d6e319fcdd11f3607352e5661f2bea9d545b354f4c7f2c82dada9d19864c13584e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcaafec875a1693099d582a517fdab78f6bd559fb432a85d6e78276bf37dfa7d5638a7609d367352b81bde988dee301654c7006495a15f579e106bb9784a759ecae622c233a1d864041b7e6a815f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he465327c35b8129b9c88e6577b7bb27f85018bb3bffc72edc2825fb143a43e06f0663eb739e514f7822a22490703ecb8d31a88c99a1d279b8134876f28f2a8ec3b82e743b2c20bc82f9d805b5b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha33496f9ae00c225170c1af039a96fd1db653d8ae905aa923c8604a9b1b73e807ae9b21b6f8689686442bdc99f16bb721f8a097766c51024f39208129ddea09844c330fcee89e9889e462fe900f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb373aa70427169c6eaab035ae6345814aa7f8390fbfa3d822a1ff383ea0e6d5898e5fe11c0a3c721ffe3941b2d128bed91091abec7fafb2ce0e116671b96aa56b5f79045bcf014bb124f121a8419;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e033c881fb9ea458cd80facc122a5a56af3132ef22ba988c8ec34a87361478b65c8cda0cc53b5dfb7d504b291c0df1325bf14adcf11d762a9b1be84f4a75fe4a507e8a3c5751326237c57016b4a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb0e0b434e7b56ee5410e188950baf5cdf58ad335f6399b0ebd4ddafb5012fadd7497046f9678ce3c281fe64c47d92a6ebf36015f8ff3a23c0877a4eeaedab5fa973ee59aa353a04907e668e55b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eed4f42fc699d1811c3bb27fc10388ec3788cbf91b9a344c049afd66516837d92b39f820627e5d4ca2ea51b965d94de29de217dc3a5c7aaac67ea5f533820ba27dc79aa40443b03fd24331518a34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120437093e2ee4f6edbf60bb54ad9b1e70ef4476f0d8f315b97e106be32dbfaf8095d364beb6b02658ead9b6412c1b1ca7cadf2b65bfb86d737a2f187ffc95685420c966c404aed49a0080d24bfb1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10373b22eefa28291565bddc0bfe73e896406d780241578cb0eccb4b24688f26cba5f9d199129dd7efa8f8b35f58508856781208611342aaa6eb6f55b36bad9eb396187bfcfcff57274d23e5a5789;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa952dda409d803e7c947b706c4fac57b0319f0b1da58aef49b351447314a113d2727fbedb04fe747cbfce0f7c350e0040134a050bf5795beb43f73a0555234a4f4af0234ed6622c5b626d0f9954;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46624e88ff489debb2c765e93dc4d65611e312986477e5645b0e6afab71b3b6db53cbbe8cc0d995d172923dcef7df0ead6a93d6ae70c8f5cd36457eaef76471474c292b4594f4fd89b2e6a9dd610;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd0b83be823545dc4844e8e06b1d680826feae44f04231740ad797773796ba37f1419be37a975457677deb69222e2f2145a907202408ee7b4ad3f77935b8cbd9c956868b06ef2da9c0778f6ac57d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1cd2f87f199f21e14e14d6f4e92d63c97a8f32ad877de5eb545c42fbe262da3f83bcfcde5d8ec1a1800ed9d96414da394109ffa4b9ebda99be91f1a41cea8fdde9b61fc9e1697b24deecfdb026e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2b4f2f6e8b873948c7307e1d71369e38f4325081e4a9d5fc5f26c7b9411f8b09fbb6d9300cf704298dd179e64aa4b4c0eb738a77b862c063b4a52085a53e36476ec597a07709954ecefb6163b49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c2923bc343e2749f6f1bd1d9d8c2eebe27232b600c0f3a3a098eabdc20dd20230a75351d2ab4adf7382d67dd84acb5e5a53a0ff9fd1a7c414b476f0711bc4a941439554080d55deb1b88d5958cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d186e2f69eb79a728a37846112d18e38a4923385c1899e2430b88e9dfad1abaf0fafec5a4c6bbef554635490797b19c23fb2c7330fce01435aa9c3ec1938235980467679c20ed1644c46067c601;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h288cc67cd6da116622bf8b0db028b28d53ad78de367d7b1f20f6ee09bdd1d1f10bfeab12fa450720c56c467f62a2b5cc1e8b198cc25149d21ce2086ba2ef982d42d34f456c8e7b71ea075217b0a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17857a24711b526644ed9fa03b47f6694eb7b8931b4ca42487b7c9519fc6f14d6b430bc8e849b2baebb754d530e587b179efca98cd3ab41594817c2890dd6eae50842895ba992b8b9fa3b28084d3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19276b4a222241164351151eb3b45d4d8080aab767b0f342f53df17c33b49ecd407e49e4b32ba6b2de7e629de3ae155a0134cfd2ce07fab94f81ebb7f1f6a84eaab17310c2d85147d02004f97d874;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h662afe0f8eab55df0d226b12a4720e716db7ed5512c5733169f45674517fe64452c0f8fe50e2b629189ecdb28ae05988489b46469e3376a29a6282030e56d481f405511aba137cbfb7a39af51c99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc28a2ebbb85a3ae85e8dc955d89f89e190317171325638054532fbe4137044bdf9934429ddcd50daae33a61e65503e71cebaca6e69dad1405fe45427c88a73e177cf64b28e651f01aaaa824e33b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd9384028976203225cb46a36f3acce847b95bb3fd44dbef649a3c20ce4bbd76dbeb7887df804120afb4ab0a6cc5b068f3b355456598a5cea22be2cf57288a2125c208ce929b26549f02970016b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heca599a5c991b0b767b79392ae7c557297a2831c70a9717c77662521f34eb356e0936ffa5bf89dfb3831bac68f1377bf041dff3a80e7db904b8742578bd417521fe5858a553f7bdd1b8b9b385412;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cda4f5b3183ec795d1412aaf1b081f9f3635d05c0963054132f7d6484cd4628d9e5345d8968addff7a64a639fe7f19debe5a77f0f865339dd38490501822ca7259e79690b92b4df613d6a941319;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc39662cb42abfc1c0b38ffe855de37c2a7dfb20615411fa9b0eb8fe1b11b44a2b6ab06425a2a43d90171c3f8a1e237c00906151cc9c204de41c9e68fc4810fd8b2b13eb4f9bac850397aa54b29f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8906fae7a371dfa3866fb005466796a112e6f155a179ebc5b53c7541cb5e665e882182f83864fed4996fd41e0ad47254011301b12f66cc4c833c8aefe240af280e25bba5e5af02f670727d8ce87;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc88d1fd402728245dd5caa1e0ed290285ea2697473607e1d23a289093b8e5ceb7e0a1a699242245333b76214ac7504d81653403b8e63c4e74b553c4c3ff28b76f9aa5cf3ed579fe7a64722faf48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f3d4a89afe5599101d153ec031ea178e32d4bc75c3cd136857db162678ff7c90c39ddcd5d64b38a1592bff840c801fd5eb25cd1b81382fcc6be64b18e917c9682d996f0c34cfbee7ad0d5af0e03;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ec88093915cfe423e3e1f83dbc34129c26c01dbfb63d6796cc6f2da2dce00843b36d399b3348f9d95074d49e14d3c0c5ba2869d522a726dc1eee79f65fc8f9a59e1cd979df36aade9d772e93b2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdb48ef4302e9ae8ea92d26045eb720a5179081c4cb5f585f0d617f8ad0cab31678db73c234f19a55c465c0ef9f4e9112e55788c36cb6b128685464a7d7fd22191240f042d2dbb227957340921eb;
        #1
        $finish();
    end
endmodule
