module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    compressor_CLA512_32 compressor_CLA512_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA512_32(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [110:0] stage1_0;
   wire [198:0] stage1_1;
   wire [187:0] stage1_2;
   wire [276:0] stage1_3;
   wire [244:0] stage1_4;
   wire [205:0] stage1_5;
   wire [242:0] stage1_6;
   wire [185:0] stage1_7;
   wire [348:0] stage1_8;
   wire [211:0] stage1_9;
   wire [181:0] stage1_10;
   wire [205:0] stage1_11;
   wire [221:0] stage1_12;
   wire [231:0] stage1_13;
   wire [231:0] stage1_14;
   wire [236:0] stage1_15;
   wire [213:0] stage1_16;
   wire [223:0] stage1_17;
   wire [202:0] stage1_18;
   wire [262:0] stage1_19;
   wire [213:0] stage1_20;
   wire [269:0] stage1_21;
   wire [273:0] stage1_22;
   wire [165:0] stage1_23;
   wire [220:0] stage1_24;
   wire [273:0] stage1_25;
   wire [190:0] stage1_26;
   wire [199:0] stage1_27;
   wire [247:0] stage1_28;
   wire [242:0] stage1_29;
   wire [206:0] stage1_30;
   wire [242:0] stage1_31;
   wire [149:0] stage1_32;
   wire [70:0] stage1_33;
   wire [62:0] stage2_0;
   wire [55:0] stage2_1;
   wire [94:0] stage2_2;
   wire [76:0] stage2_3;
   wire [118:0] stage2_4;
   wire [93:0] stage2_5;
   wire [95:0] stage2_6;
   wire [108:0] stage2_7;
   wire [97:0] stage2_8;
   wire [107:0] stage2_9;
   wire [94:0] stage2_10;
   wire [115:0] stage2_11;
   wire [101:0] stage2_12;
   wire [123:0] stage2_13;
   wire [69:0] stage2_14;
   wire [97:0] stage2_15;
   wire [124:0] stage2_16;
   wire [127:0] stage2_17;
   wire [72:0] stage2_18;
   wire [97:0] stage2_19;
   wire [109:0] stage2_20;
   wire [124:0] stage2_21;
   wire [94:0] stage2_22;
   wire [122:0] stage2_23;
   wire [89:0] stage2_24;
   wire [102:0] stage2_25;
   wire [99:0] stage2_26;
   wire [84:0] stage2_27;
   wire [170:0] stage2_28;
   wire [142:0] stage2_29;
   wire [91:0] stage2_30;
   wire [101:0] stage2_31;
   wire [73:0] stage2_32;
   wire [59:0] stage2_33;
   wire [34:0] stage2_34;
   wire [11:0] stage2_35;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [35:0] stage3_2;
   wire [27:0] stage3_3;
   wire [46:0] stage3_4;
   wire [58:0] stage3_5;
   wire [37:0] stage3_6;
   wire [46:0] stage3_7;
   wire [92:0] stage3_8;
   wire [49:0] stage3_9;
   wire [37:0] stage3_10;
   wire [54:0] stage3_11;
   wire [46:0] stage3_12;
   wire [36:0] stage3_13;
   wire [55:0] stage3_14;
   wire [70:0] stage3_15;
   wire [66:0] stage3_16;
   wire [76:0] stage3_17;
   wire [34:0] stage3_18;
   wire [69:0] stage3_19;
   wire [29:0] stage3_20;
   wire [62:0] stage3_21;
   wire [50:0] stage3_22;
   wire [45:0] stage3_23;
   wire [60:0] stage3_24;
   wire [48:0] stage3_25;
   wire [50:0] stage3_26;
   wire [54:0] stage3_27;
   wire [73:0] stage3_28;
   wire [57:0] stage3_29;
   wire [70:0] stage3_30;
   wire [57:0] stage3_31;
   wire [57:0] stage3_32;
   wire [26:0] stage3_33;
   wire [26:0] stage3_34;
   wire [12:0] stage3_35;
   wire [5:0] stage3_36;
   wire [1:0] stage3_37;
   wire [10:0] stage4_0;
   wire [15:0] stage4_1;
   wire [12:0] stage4_2;
   wire [22:0] stage4_3;
   wire [23:0] stage4_4;
   wire [45:0] stage4_5;
   wire [22:0] stage4_6;
   wire [14:0] stage4_7;
   wire [28:0] stage4_8;
   wire [41:0] stage4_9;
   wire [17:0] stage4_10;
   wire [42:0] stage4_11;
   wire [23:0] stage4_12;
   wire [18:0] stage4_13;
   wire [34:0] stage4_14;
   wire [38:0] stage4_15;
   wire [19:0] stage4_16;
   wire [42:0] stage4_17;
   wire [28:0] stage4_18;
   wire [31:0] stage4_19;
   wire [18:0] stage4_20;
   wire [18:0] stage4_21;
   wire [30:0] stage4_22;
   wire [37:0] stage4_23;
   wire [29:0] stage4_24;
   wire [18:0] stage4_25;
   wire [22:0] stage4_26;
   wire [26:0] stage4_27;
   wire [24:0] stage4_28;
   wire [25:0] stage4_29;
   wire [26:0] stage4_30;
   wire [30:0] stage4_31;
   wire [42:0] stage4_32;
   wire [18:0] stage4_33;
   wire [12:0] stage4_34;
   wire [14:0] stage4_35;
   wire [10:0] stage4_36;
   wire [2:0] stage4_37;
   wire [10:0] stage5_0;
   wire [10:0] stage5_1;
   wire [9:0] stage5_2;
   wire [5:0] stage5_3;
   wire [9:0] stage5_4;
   wire [10:0] stage5_5;
   wire [12:0] stage5_6;
   wire [19:0] stage5_7;
   wire [9:0] stage5_8;
   wire [10:0] stage5_9;
   wire [12:0] stage5_10;
   wire [15:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [9:0] stage5_14;
   wire [12:0] stage5_15;
   wire [14:0] stage5_16;
   wire [14:0] stage5_17;
   wire [16:0] stage5_18;
   wire [23:0] stage5_19;
   wire [13:0] stage5_20;
   wire [8:0] stage5_21;
   wire [16:0] stage5_22;
   wire [9:0] stage5_23;
   wire [13:0] stage5_24;
   wire [11:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [16:0] stage5_30;
   wire [12:0] stage5_31;
   wire [25:0] stage5_32;
   wire [10:0] stage5_33;
   wire [9:0] stage5_34;
   wire [7:0] stage5_35;
   wire [3:0] stage5_36;
   wire [6:0] stage5_37;
   wire [1:0] stage5_38;
   wire [6:0] stage6_0;
   wire [4:0] stage6_1;
   wire [5:0] stage6_2;
   wire [5:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [3:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [5:0] stage6_9;
   wire [3:0] stage6_10;
   wire [7:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [14:0] stage6_19;
   wire [5:0] stage6_20;
   wire [12:0] stage6_21;
   wire [7:0] stage6_22;
   wire [3:0] stage6_23;
   wire [5:0] stage6_24;
   wire [5:0] stage6_25;
   wire [4:0] stage6_26;
   wire [7:0] stage6_27;
   wire [4:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [7:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [9:0] stage6_34;
   wire [5:0] stage6_35;
   wire [2:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;
   wire [1:0] stage6_39;
   wire [0:0] stage6_40;
   wire [6:0] stage7_0;
   wire [0:0] stage7_1;
   wire [6:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [1:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [2:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [4:0] stage7_19;
   wire [5:0] stage7_20;
   wire [2:0] stage7_21;
   wire [5:0] stage7_22;
   wire [6:0] stage7_23;
   wire [0:0] stage7_24;
   wire [1:0] stage7_25;
   wire [2:0] stage7_26;
   wire [2:0] stage7_27;
   wire [6:0] stage7_28;
   wire [4:0] stage7_29;
   wire [0:0] stage7_30;
   wire [8:0] stage7_31;
   wire [0:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [2:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[11]},
      {stage0_3[22]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[12]},
      {stage0_3[23]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[13]},
      {stage0_3[24]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[14]},
      {stage0_3[25]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[15]},
      {stage0_3[26]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[16]},
      {stage0_3[27]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[17]},
      {stage0_3[28]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[18]},
      {stage0_3[29]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_2[19]},
      {stage0_3[30]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_2[20]},
      {stage0_3[31]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_2[21]},
      {stage0_3[32]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_2[22]},
      {stage0_3[33]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_2[23]},
      {stage0_3[34]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_2[24]},
      {stage0_3[35]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_2[25]},
      {stage0_3[36]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_2[26]},
      {stage0_3[37]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_2[27]},
      {stage0_3[38]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_2[28]},
      {stage0_3[39]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_2[29]},
      {stage0_3[40]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_2[30]},
      {stage0_3[41]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_2[31]},
      {stage0_3[42]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_2[32]},
      {stage0_3[43]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_2[33]},
      {stage0_3[44]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_2[34]},
      {stage0_3[45]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_2[35]},
      {stage0_3[46]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_2[36]},
      {stage0_3[47]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_2[37]},
      {stage0_3[48]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_2[38]},
      {stage0_3[49]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_2[39]},
      {stage0_3[50]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_2[40]},
      {stage0_3[51]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_2[41]},
      {stage0_3[52]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453]},
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459]},
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[460], stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465]},
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[466], stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471]},
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[472], stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483]},
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489]},
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc606_5 gpc99 (
      {stage0_0[490], stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495]},
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc606_5 gpc100 (
      {stage0_0[496], stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501]},
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[0],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[1],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[2],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[3],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[4],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[5],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[6],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[7],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[8],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[9],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[10],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[11],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[12],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[13],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[14],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[15],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[16],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[17],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[18],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[19],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[20],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[21],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[22],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[23],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[24],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[25],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[26],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[27],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[28],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[29],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[30],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[31],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[32],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[33],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[34],stage1_4[135],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[35],stage1_4[136],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[36],stage1_4[137],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[37],stage1_4[138],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452]},
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage1_5[38],stage1_4[139],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400]},
      {stage0_3[287]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[39],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405]},
      {stage0_3[288]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[40],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage0_3[289]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[41],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415]},
      {stage0_3[290]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[42],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage0_3[291]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[43],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_3[292]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[44],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430]},
      {stage0_3[293]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[45],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[431], stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435]},
      {stage0_3[294]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[46],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[436], stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440]},
      {stage0_3[295]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[47],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[441], stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445]},
      {stage0_3[296]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[48],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449], stage0_2[450]},
      {stage0_3[297]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[49],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_3[298]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[50],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460]},
      {stage0_3[299]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[51],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[461], stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465]},
      {stage0_3[300]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[52],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[466], stage0_2[467], stage0_2[468], stage0_2[469], stage0_2[470]},
      {stage0_3[301]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[53],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[471], stage0_2[472], stage0_2[473], stage0_2[474], stage0_2[475]},
      {stage0_3[302]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[54],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479], stage0_2[480]},
      {stage0_3[303]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[55],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage0_4[102]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[17],stage1_5[56],stage1_4[157],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313]},
      {stage0_4[103]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[18],stage1_5[57],stage1_4[158],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage0_4[104]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[19],stage1_5[58],stage1_4[159],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323]},
      {stage0_4[105]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[20],stage1_5[59],stage1_4[160],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328]},
      {stage0_4[106]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[21],stage1_5[60],stage1_4[161],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage0_4[107]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[22],stage1_5[61],stage1_4[162],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage0_4[108]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[23],stage1_5[62],stage1_4[163],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[109]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[24],stage1_5[63],stage1_4[164],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[110]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[25],stage1_5[64],stage1_4[165],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[111]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[26],stage1_5[65],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[112]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[27],stage1_5[66],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[113]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[28],stage1_5[67],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[114]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[29],stage1_5[68],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[115]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[30],stage1_5[69],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[116]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[31],stage1_5[70],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[117]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[32],stage1_5[71],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[118]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[33],stage1_5[72],stage1_4[173],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[119]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[34],stage1_5[73],stage1_4[174],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[120]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[35],stage1_5[74],stage1_4[175],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[121]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[36],stage1_5[75],stage1_4[176],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[122]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[37],stage1_5[76],stage1_4[177],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[123]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[38],stage1_5[77],stage1_4[178],stage1_3[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[22],stage1_6[39],stage1_5[78],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[23],stage1_6[40],stage1_5[79],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[24],stage1_6[41],stage1_5[80],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[25],stage1_6[42],stage1_5[81],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[26],stage1_6[43],stage1_5[82],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[27],stage1_6[44],stage1_5[83],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[28],stage1_6[45],stage1_5[84],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[29],stage1_6[46],stage1_5[85],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[30],stage1_6[47],stage1_5[86],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[31],stage1_6[48],stage1_5[87],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[32],stage1_6[49],stage1_5[88],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[33],stage1_6[50],stage1_5[89],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[34],stage1_6[51],stage1_5[90],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[35],stage1_6[52],stage1_5[91],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[36],stage1_6[53],stage1_5[92],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[37],stage1_6[54],stage1_5[93],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[38],stage1_6[55],stage1_5[94],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[39],stage1_6[56],stage1_5[95],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[40],stage1_6[57],stage1_5[96],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[41],stage1_6[58],stage1_5[97],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[42],stage1_6[59],stage1_5[98],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[43],stage1_6[60],stage1_5[99],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[44],stage1_6[61],stage1_5[100],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[45],stage1_6[62],stage1_5[101],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[46],stage1_6[63],stage1_5[102],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[47],stage1_6[64],stage1_5[103],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[48],stage1_6[65],stage1_5[104],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[49],stage1_6[66],stage1_5[105],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[50],stage1_6[67],stage1_5[106],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[51],stage1_6[68],stage1_5[107],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[52],stage1_6[69],stage1_5[108],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[53],stage1_6[70],stage1_5[109],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[54],stage1_6[71],stage1_5[110],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[55],stage1_6[72],stage1_5[111],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[56],stage1_6[73],stage1_5[112],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[57],stage1_6[74],stage1_5[113],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[58],stage1_6[75],stage1_5[114],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[59],stage1_6[76],stage1_5[115],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[60],stage1_6[77],stage1_5[116],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[61],stage1_6[78],stage1_5[117],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[62],stage1_6[79],stage1_5[118],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[63],stage1_6[80],stage1_5[119],stage1_4[220]}
   );
   gpc606_5 gpc221 (
      {stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[64],stage1_6[81],stage1_5[120],stage1_4[221]}
   );
   gpc606_5 gpc222 (
      {stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[65],stage1_6[82],stage1_5[121],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[66],stage1_6[83],stage1_5[122],stage1_4[223]}
   );
   gpc606_5 gpc224 (
      {stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[67],stage1_6[84],stage1_5[123],stage1_4[224]}
   );
   gpc606_5 gpc225 (
      {stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[68],stage1_6[85],stage1_5[124],stage1_4[225]}
   );
   gpc606_5 gpc226 (
      {stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[69],stage1_6[86],stage1_5[125],stage1_4[226]}
   );
   gpc606_5 gpc227 (
      {stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[70],stage1_6[87],stage1_5[126],stage1_4[227]}
   );
   gpc606_5 gpc228 (
      {stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[71],stage1_6[88],stage1_5[127],stage1_4[228]}
   );
   gpc606_5 gpc229 (
      {stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[72],stage1_6[89],stage1_5[128],stage1_4[229]}
   );
   gpc606_5 gpc230 (
      {stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[73],stage1_6[90],stage1_5[129],stage1_4[230]}
   );
   gpc606_5 gpc231 (
      {stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[74],stage1_6[91],stage1_5[130],stage1_4[231]}
   );
   gpc606_5 gpc232 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[75],stage1_6[92],stage1_5[131],stage1_4[232]}
   );
   gpc606_5 gpc233 (
      {stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[76],stage1_6[93],stage1_5[132],stage1_4[233]}
   );
   gpc606_5 gpc234 (
      {stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[77],stage1_6[94],stage1_5[133],stage1_4[234]}
   );
   gpc606_5 gpc235 (
      {stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[78],stage1_6[95],stage1_5[134],stage1_4[235]}
   );
   gpc606_5 gpc236 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[79],stage1_6[96],stage1_5[135],stage1_4[236]}
   );
   gpc615_5 gpc237 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[132]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[80],stage1_6[97],stage1_5[136],stage1_4[237]}
   );
   gpc615_5 gpc238 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[133]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[81],stage1_6[98],stage1_5[137],stage1_4[238]}
   );
   gpc615_5 gpc239 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[134]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[82],stage1_6[99],stage1_5[138],stage1_4[239]}
   );
   gpc615_5 gpc240 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[135]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[83],stage1_6[100],stage1_5[139],stage1_4[240]}
   );
   gpc615_5 gpc241 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[136]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[84],stage1_6[101],stage1_5[140],stage1_4[241]}
   );
   gpc615_5 gpc242 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[137]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[85],stage1_6[102],stage1_5[141],stage1_4[242]}
   );
   gpc615_5 gpc243 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[138]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[86],stage1_6[103],stage1_5[142],stage1_4[243]}
   );
   gpc615_5 gpc244 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[139]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[87],stage1_6[104],stage1_5[143],stage1_4[244]}
   );
   gpc606_5 gpc245 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[66],stage1_7[88],stage1_6[105],stage1_5[144]}
   );
   gpc606_5 gpc246 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[67],stage1_7[89],stage1_6[106],stage1_5[145]}
   );
   gpc606_5 gpc247 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[68],stage1_7[90],stage1_6[107],stage1_5[146]}
   );
   gpc606_5 gpc248 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[69],stage1_7[91],stage1_6[108],stage1_5[147]}
   );
   gpc606_5 gpc249 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[70],stage1_7[92],stage1_6[109],stage1_5[148]}
   );
   gpc606_5 gpc250 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[71],stage1_7[93],stage1_6[110],stage1_5[149]}
   );
   gpc606_5 gpc251 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[72],stage1_7[94],stage1_6[111],stage1_5[150]}
   );
   gpc606_5 gpc252 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[73],stage1_7[95],stage1_6[112],stage1_5[151]}
   );
   gpc606_5 gpc253 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[74],stage1_7[96],stage1_6[113],stage1_5[152]}
   );
   gpc606_5 gpc254 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[75],stage1_7[97],stage1_6[114],stage1_5[153]}
   );
   gpc606_5 gpc255 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[76],stage1_7[98],stage1_6[115],stage1_5[154]}
   );
   gpc606_5 gpc256 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[77],stage1_7[99],stage1_6[116],stage1_5[155]}
   );
   gpc606_5 gpc257 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[78],stage1_7[100],stage1_6[117],stage1_5[156]}
   );
   gpc606_5 gpc258 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[79],stage1_7[101],stage1_6[118],stage1_5[157]}
   );
   gpc606_5 gpc259 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[80],stage1_7[102],stage1_6[119],stage1_5[158]}
   );
   gpc606_5 gpc260 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[81],stage1_7[103],stage1_6[120],stage1_5[159]}
   );
   gpc606_5 gpc261 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[82],stage1_7[104],stage1_6[121],stage1_5[160]}
   );
   gpc606_5 gpc262 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[83],stage1_7[105],stage1_6[122],stage1_5[161]}
   );
   gpc606_5 gpc263 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[84],stage1_7[106],stage1_6[123],stage1_5[162]}
   );
   gpc606_5 gpc264 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[85],stage1_7[107],stage1_6[124],stage1_5[163]}
   );
   gpc606_5 gpc265 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[86],stage1_7[108],stage1_6[125],stage1_5[164]}
   );
   gpc606_5 gpc266 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[87],stage1_7[109],stage1_6[126],stage1_5[165]}
   );
   gpc606_5 gpc267 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276], stage0_5[277]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[88],stage1_7[110],stage1_6[127],stage1_5[166]}
   );
   gpc606_5 gpc268 (
      {stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282], stage0_5[283]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[89],stage1_7[111],stage1_6[128],stage1_5[167]}
   );
   gpc606_5 gpc269 (
      {stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288], stage0_5[289]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[90],stage1_7[112],stage1_6[129],stage1_5[168]}
   );
   gpc606_5 gpc270 (
      {stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[91],stage1_7[113],stage1_6[130],stage1_5[169]}
   );
   gpc606_5 gpc271 (
      {stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[92],stage1_7[114],stage1_6[131],stage1_5[170]}
   );
   gpc606_5 gpc272 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306], stage0_5[307]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[93],stage1_7[115],stage1_6[132],stage1_5[171]}
   );
   gpc606_5 gpc273 (
      {stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312], stage0_5[313]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[94],stage1_7[116],stage1_6[133],stage1_5[172]}
   );
   gpc606_5 gpc274 (
      {stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318], stage0_5[319]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[95],stage1_7[117],stage1_6[134],stage1_5[173]}
   );
   gpc606_5 gpc275 (
      {stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[96],stage1_7[118],stage1_6[135],stage1_5[174]}
   );
   gpc606_5 gpc276 (
      {stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[97],stage1_7[119],stage1_6[136],stage1_5[175]}
   );
   gpc606_5 gpc277 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336], stage0_5[337]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[98],stage1_7[120],stage1_6[137],stage1_5[176]}
   );
   gpc606_5 gpc278 (
      {stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342], stage0_5[343]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[99],stage1_7[121],stage1_6[138],stage1_5[177]}
   );
   gpc606_5 gpc279 (
      {stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348], stage0_5[349]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[100],stage1_7[122],stage1_6[139],stage1_5[178]}
   );
   gpc606_5 gpc280 (
      {stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354], stage0_5[355]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[101],stage1_7[123],stage1_6[140],stage1_5[179]}
   );
   gpc606_5 gpc281 (
      {stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360], stage0_5[361]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[102],stage1_7[124],stage1_6[141],stage1_5[180]}
   );
   gpc606_5 gpc282 (
      {stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366], stage0_5[367]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[103],stage1_7[125],stage1_6[142],stage1_5[181]}
   );
   gpc606_5 gpc283 (
      {stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372], stage0_5[373]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[104],stage1_7[126],stage1_6[143],stage1_5[182]}
   );
   gpc606_5 gpc284 (
      {stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378], stage0_5[379]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[105],stage1_7[127],stage1_6[144],stage1_5[183]}
   );
   gpc606_5 gpc285 (
      {stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384], stage0_5[385]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[106],stage1_7[128],stage1_6[145],stage1_5[184]}
   );
   gpc606_5 gpc286 (
      {stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390], stage0_5[391]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[107],stage1_7[129],stage1_6[146],stage1_5[185]}
   );
   gpc606_5 gpc287 (
      {stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396], stage0_5[397]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[108],stage1_7[130],stage1_6[147],stage1_5[186]}
   );
   gpc606_5 gpc288 (
      {stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402], stage0_5[403]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[109],stage1_7[131],stage1_6[148],stage1_5[187]}
   );
   gpc606_5 gpc289 (
      {stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408], stage0_5[409]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[110],stage1_7[132],stage1_6[149],stage1_5[188]}
   );
   gpc606_5 gpc290 (
      {stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414], stage0_5[415]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[111],stage1_7[133],stage1_6[150],stage1_5[189]}
   );
   gpc606_5 gpc291 (
      {stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420], stage0_5[421]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[112],stage1_7[134],stage1_6[151],stage1_5[190]}
   );
   gpc606_5 gpc292 (
      {stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426], stage0_5[427]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[113],stage1_7[135],stage1_6[152],stage1_5[191]}
   );
   gpc606_5 gpc293 (
      {stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432], stage0_5[433]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[114],stage1_7[136],stage1_6[153],stage1_5[192]}
   );
   gpc606_5 gpc294 (
      {stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438], stage0_5[439]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[115],stage1_7[137],stage1_6[154],stage1_5[193]}
   );
   gpc606_5 gpc295 (
      {stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444], stage0_5[445]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[116],stage1_7[138],stage1_6[155],stage1_5[194]}
   );
   gpc606_5 gpc296 (
      {stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450], stage0_5[451]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[117],stage1_7[139],stage1_6[156],stage1_5[195]}
   );
   gpc606_5 gpc297 (
      {stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456], stage0_5[457]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[118],stage1_7[140],stage1_6[157],stage1_5[196]}
   );
   gpc606_5 gpc298 (
      {stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462], stage0_5[463]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[119],stage1_7[141],stage1_6[158],stage1_5[197]}
   );
   gpc606_5 gpc299 (
      {stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468], stage0_5[469]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[120],stage1_7[142],stage1_6[159],stage1_5[198]}
   );
   gpc606_5 gpc300 (
      {stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474], stage0_5[475]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[121],stage1_7[143],stage1_6[160],stage1_5[199]}
   );
   gpc606_5 gpc301 (
      {stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480], stage0_5[481]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[122],stage1_7[144],stage1_6[161],stage1_5[200]}
   );
   gpc606_5 gpc302 (
      {stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486], stage0_5[487]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[123],stage1_7[145],stage1_6[162],stage1_5[201]}
   );
   gpc606_5 gpc303 (
      {stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492], stage0_5[493]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[124],stage1_7[146],stage1_6[163],stage1_5[202]}
   );
   gpc606_5 gpc304 (
      {stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498], stage0_5[499]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[125],stage1_7[147],stage1_6[164],stage1_5[203]}
   );
   gpc606_5 gpc305 (
      {stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504], stage0_5[505]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[126],stage1_7[148],stage1_6[165],stage1_5[204]}
   );
   gpc606_5 gpc306 (
      {stage0_5[506], stage0_5[507], stage0_5[508], stage0_5[509], stage0_5[510], stage0_5[511]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[127],stage1_7[149],stage1_6[166],stage1_5[205]}
   );
   gpc615_5 gpc307 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[372]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[62],stage1_8[128],stage1_7[150],stage1_6[167]}
   );
   gpc615_5 gpc308 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[373]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[63],stage1_8[129],stage1_7[151],stage1_6[168]}
   );
   gpc615_5 gpc309 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[374]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[64],stage1_8[130],stage1_7[152],stage1_6[169]}
   );
   gpc615_5 gpc310 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[375]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[65],stage1_8[131],stage1_7[153],stage1_6[170]}
   );
   gpc615_5 gpc311 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[376]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[66],stage1_8[132],stage1_7[154],stage1_6[171]}
   );
   gpc615_5 gpc312 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[377]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[67],stage1_8[133],stage1_7[155],stage1_6[172]}
   );
   gpc615_5 gpc313 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[378]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[68],stage1_8[134],stage1_7[156],stage1_6[173]}
   );
   gpc615_5 gpc314 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[379]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[69],stage1_8[135],stage1_7[157],stage1_6[174]}
   );
   gpc615_5 gpc315 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[380]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[70],stage1_8[136],stage1_7[158],stage1_6[175]}
   );
   gpc615_5 gpc316 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[381]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[71],stage1_8[137],stage1_7[159],stage1_6[176]}
   );
   gpc615_5 gpc317 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[60]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[10],stage1_9[72],stage1_8[138],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[61]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[11],stage1_9[73],stage1_8[139],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[62]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[12],stage1_9[74],stage1_8[140],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[63]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[13],stage1_9[75],stage1_8[141],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[64]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[14],stage1_9[76],stage1_8[142],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[65]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[15],stage1_9[77],stage1_8[143],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[66]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[16],stage1_9[78],stage1_8[144],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[67]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[17],stage1_9[79],stage1_8[145],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[68]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[18],stage1_9[80],stage1_8[146],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[69]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[19],stage1_9[81],stage1_8[147],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[70]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[20],stage1_9[82],stage1_8[148],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[71]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[21],stage1_9[83],stage1_8[149],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[72]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[22],stage1_9[84],stage1_8[150],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[73]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[23],stage1_9[85],stage1_8[151],stage1_7[173]}
   );
   gpc615_5 gpc331 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[74]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[24],stage1_9[86],stage1_8[152],stage1_7[174]}
   );
   gpc615_5 gpc332 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[75]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[25],stage1_9[87],stage1_8[153],stage1_7[175]}
   );
   gpc615_5 gpc333 (
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466]},
      {stage0_8[76]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[26],stage1_9[88],stage1_8[154],stage1_7[176]}
   );
   gpc615_5 gpc334 (
      {stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471]},
      {stage0_8[77]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[27],stage1_9[89],stage1_8[155],stage1_7[177]}
   );
   gpc615_5 gpc335 (
      {stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475], stage0_7[476]},
      {stage0_8[78]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[28],stage1_9[90],stage1_8[156],stage1_7[178]}
   );
   gpc615_5 gpc336 (
      {stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480], stage0_7[481]},
      {stage0_8[79]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[29],stage1_9[91],stage1_8[157],stage1_7[179]}
   );
   gpc615_5 gpc337 (
      {stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485], stage0_7[486]},
      {stage0_8[80]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[30],stage1_9[92],stage1_8[158],stage1_7[180]}
   );
   gpc615_5 gpc338 (
      {stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490], stage0_7[491]},
      {stage0_8[81]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[31],stage1_9[93],stage1_8[159],stage1_7[181]}
   );
   gpc615_5 gpc339 (
      {stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495], stage0_7[496]},
      {stage0_8[82]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[32],stage1_9[94],stage1_8[160],stage1_7[182]}
   );
   gpc615_5 gpc340 (
      {stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500], stage0_7[501]},
      {stage0_8[83]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[33],stage1_9[95],stage1_8[161],stage1_7[183]}
   );
   gpc615_5 gpc341 (
      {stage0_7[502], stage0_7[503], stage0_7[504], stage0_7[505], stage0_7[506]},
      {stage0_8[84]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[34],stage1_9[96],stage1_8[162],stage1_7[184]}
   );
   gpc615_5 gpc342 (
      {stage0_7[507], stage0_7[508], stage0_7[509], stage0_7[510], stage0_7[511]},
      {stage0_8[85]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[35],stage1_9[97],stage1_8[163],stage1_7[185]}
   );
   gpc606_5 gpc343 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[26],stage1_10[36],stage1_9[98],stage1_8[164]}
   );
   gpc606_5 gpc344 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[27],stage1_10[37],stage1_9[99],stage1_8[165]}
   );
   gpc606_5 gpc345 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[28],stage1_10[38],stage1_9[100],stage1_8[166]}
   );
   gpc606_5 gpc346 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[29],stage1_10[39],stage1_9[101],stage1_8[167]}
   );
   gpc606_5 gpc347 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[30],stage1_10[40],stage1_9[102],stage1_8[168]}
   );
   gpc606_5 gpc348 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[31],stage1_10[41],stage1_9[103],stage1_8[169]}
   );
   gpc606_5 gpc349 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[32],stage1_10[42],stage1_9[104],stage1_8[170]}
   );
   gpc606_5 gpc350 (
      {stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[33],stage1_10[43],stage1_9[105],stage1_8[171]}
   );
   gpc606_5 gpc351 (
      {stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[34],stage1_10[44],stage1_9[106],stage1_8[172]}
   );
   gpc606_5 gpc352 (
      {stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[35],stage1_10[45],stage1_9[107],stage1_8[173]}
   );
   gpc606_5 gpc353 (
      {stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[36],stage1_10[46],stage1_9[108],stage1_8[174]}
   );
   gpc606_5 gpc354 (
      {stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[37],stage1_10[47],stage1_9[109],stage1_8[175]}
   );
   gpc606_5 gpc355 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[38],stage1_10[48],stage1_9[110],stage1_8[176]}
   );
   gpc606_5 gpc356 (
      {stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[39],stage1_10[49],stage1_9[111],stage1_8[177]}
   );
   gpc606_5 gpc357 (
      {stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[40],stage1_10[50],stage1_9[112],stage1_8[178]}
   );
   gpc606_5 gpc358 (
      {stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[41],stage1_10[51],stage1_9[113],stage1_8[179]}
   );
   gpc606_5 gpc359 (
      {stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[42],stage1_10[52],stage1_9[114],stage1_8[180]}
   );
   gpc606_5 gpc360 (
      {stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[43],stage1_10[53],stage1_9[115],stage1_8[181]}
   );
   gpc606_5 gpc361 (
      {stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[44],stage1_10[54],stage1_9[116],stage1_8[182]}
   );
   gpc606_5 gpc362 (
      {stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[45],stage1_10[55],stage1_9[117],stage1_8[183]}
   );
   gpc606_5 gpc363 (
      {stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[46],stage1_10[56],stage1_9[118],stage1_8[184]}
   );
   gpc606_5 gpc364 (
      {stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[47],stage1_10[57],stage1_9[119],stage1_8[185]}
   );
   gpc606_5 gpc365 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[48],stage1_10[58],stage1_9[120],stage1_8[186]}
   );
   gpc606_5 gpc366 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[49],stage1_10[59],stage1_9[121],stage1_8[187]}
   );
   gpc606_5 gpc367 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[50],stage1_10[60],stage1_9[122],stage1_8[188]}
   );
   gpc606_5 gpc368 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[51],stage1_10[61],stage1_9[123],stage1_8[189]}
   );
   gpc606_5 gpc369 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[52],stage1_10[62],stage1_9[124],stage1_8[190]}
   );
   gpc606_5 gpc370 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[53],stage1_10[63],stage1_9[125],stage1_8[191]}
   );
   gpc606_5 gpc371 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[54],stage1_10[64],stage1_9[126],stage1_8[192]}
   );
   gpc606_5 gpc372 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[55],stage1_10[65],stage1_9[127],stage1_8[193]}
   );
   gpc606_5 gpc373 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[56],stage1_10[66],stage1_9[128],stage1_8[194]}
   );
   gpc606_5 gpc374 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[57],stage1_10[67],stage1_9[129],stage1_8[195]}
   );
   gpc606_5 gpc375 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[58],stage1_10[68],stage1_9[130],stage1_8[196]}
   );
   gpc606_5 gpc376 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[59],stage1_10[69],stage1_9[131],stage1_8[197]}
   );
   gpc606_5 gpc377 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[60],stage1_10[70],stage1_9[132],stage1_8[198]}
   );
   gpc606_5 gpc378 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[61],stage1_10[71],stage1_9[133],stage1_8[199]}
   );
   gpc606_5 gpc379 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[62],stage1_10[72],stage1_9[134],stage1_8[200]}
   );
   gpc606_5 gpc380 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[63],stage1_10[73],stage1_9[135],stage1_8[201]}
   );
   gpc606_5 gpc381 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[64],stage1_10[74],stage1_9[136],stage1_8[202]}
   );
   gpc606_5 gpc382 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[65],stage1_10[75],stage1_9[137],stage1_8[203]}
   );
   gpc606_5 gpc383 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[66],stage1_10[76],stage1_9[138],stage1_8[204]}
   );
   gpc615_5 gpc384 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_9[156]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[67],stage1_10[77],stage1_9[139],stage1_8[205]}
   );
   gpc615_5 gpc385 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_9[157]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[68],stage1_10[78],stage1_9[140],stage1_8[206]}
   );
   gpc615_5 gpc386 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346]},
      {stage0_9[158]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[69],stage1_10[79],stage1_9[141],stage1_8[207]}
   );
   gpc615_5 gpc387 (
      {stage0_8[347], stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351]},
      {stage0_9[159]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[70],stage1_10[80],stage1_9[142],stage1_8[208]}
   );
   gpc615_5 gpc388 (
      {stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355], stage0_8[356]},
      {stage0_9[160]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[71],stage1_10[81],stage1_9[143],stage1_8[209]}
   );
   gpc615_5 gpc389 (
      {stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_9[161]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[72],stage1_10[82],stage1_9[144],stage1_8[210]}
   );
   gpc615_5 gpc390 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_9[162]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[73],stage1_10[83],stage1_9[145],stage1_8[211]}
   );
   gpc615_5 gpc391 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_9[163]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[74],stage1_10[84],stage1_9[146],stage1_8[212]}
   );
   gpc615_5 gpc392 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376]},
      {stage0_9[164]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[75],stage1_10[85],stage1_9[147],stage1_8[213]}
   );
   gpc606_5 gpc393 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[50],stage1_11[76],stage1_10[86],stage1_9[148]}
   );
   gpc606_5 gpc394 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[51],stage1_11[77],stage1_10[87],stage1_9[149]}
   );
   gpc606_5 gpc395 (
      {stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[52],stage1_11[78],stage1_10[88],stage1_9[150]}
   );
   gpc606_5 gpc396 (
      {stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[53],stage1_11[79],stage1_10[89],stage1_9[151]}
   );
   gpc606_5 gpc397 (
      {stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[54],stage1_11[80],stage1_10[90],stage1_9[152]}
   );
   gpc606_5 gpc398 (
      {stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[55],stage1_11[81],stage1_10[91],stage1_9[153]}
   );
   gpc606_5 gpc399 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[56],stage1_11[82],stage1_10[92],stage1_9[154]}
   );
   gpc606_5 gpc400 (
      {stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[57],stage1_11[83],stage1_10[93],stage1_9[155]}
   );
   gpc606_5 gpc401 (
      {stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[58],stage1_11[84],stage1_10[94],stage1_9[156]}
   );
   gpc606_5 gpc402 (
      {stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[59],stage1_11[85],stage1_10[95],stage1_9[157]}
   );
   gpc606_5 gpc403 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[60],stage1_11[86],stage1_10[96],stage1_9[158]}
   );
   gpc606_5 gpc404 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[61],stage1_11[87],stage1_10[97],stage1_9[159]}
   );
   gpc606_5 gpc405 (
      {stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[62],stage1_11[88],stage1_10[98],stage1_9[160]}
   );
   gpc606_5 gpc406 (
      {stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[63],stage1_11[89],stage1_10[99],stage1_9[161]}
   );
   gpc606_5 gpc407 (
      {stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[64],stage1_11[90],stage1_10[100],stage1_9[162]}
   );
   gpc606_5 gpc408 (
      {stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[65],stage1_11[91],stage1_10[101],stage1_9[163]}
   );
   gpc606_5 gpc409 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[66],stage1_11[92],stage1_10[102],stage1_9[164]}
   );
   gpc606_5 gpc410 (
      {stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[67],stage1_11[93],stage1_10[103],stage1_9[165]}
   );
   gpc606_5 gpc411 (
      {stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[68],stage1_11[94],stage1_10[104],stage1_9[166]}
   );
   gpc606_5 gpc412 (
      {stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[69],stage1_11[95],stage1_10[105],stage1_9[167]}
   );
   gpc606_5 gpc413 (
      {stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[70],stage1_11[96],stage1_10[106],stage1_9[168]}
   );
   gpc606_5 gpc414 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[71],stage1_11[97],stage1_10[107],stage1_9[169]}
   );
   gpc606_5 gpc415 (
      {stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[72],stage1_11[98],stage1_10[108],stage1_9[170]}
   );
   gpc606_5 gpc416 (
      {stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[73],stage1_11[99],stage1_10[109],stage1_9[171]}
   );
   gpc606_5 gpc417 (
      {stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[74],stage1_11[100],stage1_10[110],stage1_9[172]}
   );
   gpc606_5 gpc418 (
      {stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[75],stage1_11[101],stage1_10[111],stage1_9[173]}
   );
   gpc606_5 gpc419 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[76],stage1_11[102],stage1_10[112],stage1_9[174]}
   );
   gpc606_5 gpc420 (
      {stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[77],stage1_11[103],stage1_10[113],stage1_9[175]}
   );
   gpc606_5 gpc421 (
      {stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[78],stage1_11[104],stage1_10[114],stage1_9[176]}
   );
   gpc606_5 gpc422 (
      {stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[79],stage1_11[105],stage1_10[115],stage1_9[177]}
   );
   gpc606_5 gpc423 (
      {stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[80],stage1_11[106],stage1_10[116],stage1_9[178]}
   );
   gpc606_5 gpc424 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[81],stage1_11[107],stage1_10[117],stage1_9[179]}
   );
   gpc606_5 gpc425 (
      {stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[82],stage1_11[108],stage1_10[118],stage1_9[180]}
   );
   gpc606_5 gpc426 (
      {stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[83],stage1_11[109],stage1_10[119],stage1_9[181]}
   );
   gpc606_5 gpc427 (
      {stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[84],stage1_11[110],stage1_10[120],stage1_9[182]}
   );
   gpc606_5 gpc428 (
      {stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[85],stage1_11[111],stage1_10[121],stage1_9[183]}
   );
   gpc606_5 gpc429 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[86],stage1_11[112],stage1_10[122],stage1_9[184]}
   );
   gpc606_5 gpc430 (
      {stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[87],stage1_11[113],stage1_10[123],stage1_9[185]}
   );
   gpc606_5 gpc431 (
      {stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[88],stage1_11[114],stage1_10[124],stage1_9[186]}
   );
   gpc615_5 gpc432 (
      {stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403]},
      {stage0_10[300]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[89],stage1_11[115],stage1_10[125],stage1_9[187]}
   );
   gpc615_5 gpc433 (
      {stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_10[301]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[90],stage1_11[116],stage1_10[126],stage1_9[188]}
   );
   gpc615_5 gpc434 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_10[302]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[91],stage1_11[117],stage1_10[127],stage1_9[189]}
   );
   gpc615_5 gpc435 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418]},
      {stage0_10[303]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[92],stage1_11[118],stage1_10[128],stage1_9[190]}
   );
   gpc615_5 gpc436 (
      {stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_10[304]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[93],stage1_11[119],stage1_10[129],stage1_9[191]}
   );
   gpc615_5 gpc437 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428]},
      {stage0_10[305]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[94],stage1_11[120],stage1_10[130],stage1_9[192]}
   );
   gpc615_5 gpc438 (
      {stage0_9[429], stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433]},
      {stage0_10[306]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[95],stage1_11[121],stage1_10[131],stage1_9[193]}
   );
   gpc615_5 gpc439 (
      {stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437], stage0_9[438]},
      {stage0_10[307]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[96],stage1_11[122],stage1_10[132],stage1_9[194]}
   );
   gpc615_5 gpc440 (
      {stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_10[308]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[97],stage1_11[123],stage1_10[133],stage1_9[195]}
   );
   gpc615_5 gpc441 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448]},
      {stage0_10[309]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[98],stage1_11[124],stage1_10[134],stage1_9[196]}
   );
   gpc615_5 gpc442 (
      {stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_10[310]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[99],stage1_11[125],stage1_10[135],stage1_9[197]}
   );
   gpc615_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458]},
      {stage0_10[311]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[100],stage1_11[126],stage1_10[136],stage1_9[198]}
   );
   gpc615_5 gpc444 (
      {stage0_9[459], stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463]},
      {stage0_10[312]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[101],stage1_11[127],stage1_10[137],stage1_9[199]}
   );
   gpc615_5 gpc445 (
      {stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467], stage0_9[468]},
      {stage0_10[313]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[102],stage1_11[128],stage1_10[138],stage1_9[200]}
   );
   gpc615_5 gpc446 (
      {stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_10[314]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[103],stage1_11[129],stage1_10[139],stage1_9[201]}
   );
   gpc615_5 gpc447 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478]},
      {stage0_10[315]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[104],stage1_11[130],stage1_10[140],stage1_9[202]}
   );
   gpc615_5 gpc448 (
      {stage0_9[479], stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483]},
      {stage0_10[316]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[105],stage1_11[131],stage1_10[141],stage1_9[203]}
   );
   gpc615_5 gpc449 (
      {stage0_9[484], stage0_9[485], stage0_9[486], stage0_9[487], stage0_9[488]},
      {stage0_10[317]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[106],stage1_11[132],stage1_10[142],stage1_9[204]}
   );
   gpc615_5 gpc450 (
      {stage0_9[489], stage0_9[490], stage0_9[491], stage0_9[492], stage0_9[493]},
      {stage0_10[318]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[107],stage1_11[133],stage1_10[143],stage1_9[205]}
   );
   gpc615_5 gpc451 (
      {stage0_9[494], stage0_9[495], stage0_9[496], stage0_9[497], stage0_9[498]},
      {stage0_10[319]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[108],stage1_11[134],stage1_10[144],stage1_9[206]}
   );
   gpc615_5 gpc452 (
      {stage0_9[499], stage0_9[500], stage0_9[501], stage0_9[502], stage0_9[503]},
      {stage0_10[320]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[109],stage1_11[135],stage1_10[145],stage1_9[207]}
   );
   gpc615_5 gpc453 (
      {stage0_9[504], stage0_9[505], stage0_9[506], stage0_9[507], stage0_9[508]},
      {stage0_10[321]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[110],stage1_11[136],stage1_10[146],stage1_9[208]}
   );
   gpc606_5 gpc454 (
      {stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[61],stage1_12[111],stage1_11[137],stage1_10[147]}
   );
   gpc606_5 gpc455 (
      {stage0_10[328], stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[62],stage1_12[112],stage1_11[138],stage1_10[148]}
   );
   gpc606_5 gpc456 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[63],stage1_12[113],stage1_11[139],stage1_10[149]}
   );
   gpc606_5 gpc457 (
      {stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[64],stage1_12[114],stage1_11[140],stage1_10[150]}
   );
   gpc606_5 gpc458 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[65],stage1_12[115],stage1_11[141],stage1_10[151]}
   );
   gpc606_5 gpc459 (
      {stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[66],stage1_12[116],stage1_11[142],stage1_10[152]}
   );
   gpc606_5 gpc460 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[67],stage1_12[117],stage1_11[143],stage1_10[153]}
   );
   gpc606_5 gpc461 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[68],stage1_12[118],stage1_11[144],stage1_10[154]}
   );
   gpc606_5 gpc462 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[69],stage1_12[119],stage1_11[145],stage1_10[155]}
   );
   gpc606_5 gpc463 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[70],stage1_12[120],stage1_11[146],stage1_10[156]}
   );
   gpc606_5 gpc464 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[71],stage1_12[121],stage1_11[147],stage1_10[157]}
   );
   gpc606_5 gpc465 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[72],stage1_12[122],stage1_11[148],stage1_10[158]}
   );
   gpc606_5 gpc466 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[73],stage1_12[123],stage1_11[149],stage1_10[159]}
   );
   gpc606_5 gpc467 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[74],stage1_12[124],stage1_11[150],stage1_10[160]}
   );
   gpc606_5 gpc468 (
      {stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[75],stage1_12[125],stage1_11[151],stage1_10[161]}
   );
   gpc615_5 gpc469 (
      {stage0_10[412], stage0_10[413], stage0_10[414], stage0_10[415], stage0_10[416]},
      {stage0_11[366]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[76],stage1_12[126],stage1_11[152],stage1_10[162]}
   );
   gpc615_5 gpc470 (
      {stage0_10[417], stage0_10[418], stage0_10[419], stage0_10[420], stage0_10[421]},
      {stage0_11[367]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[77],stage1_12[127],stage1_11[153],stage1_10[163]}
   );
   gpc615_5 gpc471 (
      {stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425], stage0_10[426]},
      {stage0_11[368]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[78],stage1_12[128],stage1_11[154],stage1_10[164]}
   );
   gpc615_5 gpc472 (
      {stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage0_11[369]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[79],stage1_12[129],stage1_11[155],stage1_10[165]}
   );
   gpc615_5 gpc473 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[370]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[80],stage1_12[130],stage1_11[156],stage1_10[166]}
   );
   gpc615_5 gpc474 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[371]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[81],stage1_12[131],stage1_11[157],stage1_10[167]}
   );
   gpc615_5 gpc475 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[372]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[82],stage1_12[132],stage1_11[158],stage1_10[168]}
   );
   gpc615_5 gpc476 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[373]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[83],stage1_12[133],stage1_11[159],stage1_10[169]}
   );
   gpc615_5 gpc477 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[374]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[84],stage1_12[134],stage1_11[160],stage1_10[170]}
   );
   gpc615_5 gpc478 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[375]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[85],stage1_12[135],stage1_11[161],stage1_10[171]}
   );
   gpc615_5 gpc479 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[376]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[86],stage1_12[136],stage1_11[162],stage1_10[172]}
   );
   gpc615_5 gpc480 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[377]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[87],stage1_12[137],stage1_11[163],stage1_10[173]}
   );
   gpc615_5 gpc481 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[378]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[88],stage1_12[138],stage1_11[164],stage1_10[174]}
   );
   gpc615_5 gpc482 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[379]},
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage1_14[28],stage1_13[89],stage1_12[139],stage1_11[165],stage1_10[175]}
   );
   gpc615_5 gpc483 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[380]},
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage1_14[29],stage1_13[90],stage1_12[140],stage1_11[166],stage1_10[176]}
   );
   gpc615_5 gpc484 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[381]},
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage1_14[30],stage1_13[91],stage1_12[141],stage1_11[167],stage1_10[177]}
   );
   gpc615_5 gpc485 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[382]},
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage1_14[31],stage1_13[92],stage1_12[142],stage1_11[168],stage1_10[178]}
   );
   gpc615_5 gpc486 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[383]},
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage1_14[32],stage1_13[93],stage1_12[143],stage1_11[169],stage1_10[179]}
   );
   gpc615_5 gpc487 (
      {stage0_10[502], stage0_10[503], stage0_10[504], stage0_10[505], stage0_10[506]},
      {stage0_11[384]},
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage1_14[33],stage1_13[94],stage1_12[144],stage1_11[170],stage1_10[180]}
   );
   gpc615_5 gpc488 (
      {stage0_10[507], stage0_10[508], stage0_10[509], stage0_10[510], stage0_10[511]},
      {stage0_11[385]},
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage1_14[34],stage1_13[95],stage1_12[145],stage1_11[171],stage1_10[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[210]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[35],stage1_13[96],stage1_12[146],stage1_11[172]}
   );
   gpc615_5 gpc490 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[211]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[36],stage1_13[97],stage1_12[147],stage1_11[173]}
   );
   gpc615_5 gpc491 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[212]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[37],stage1_13[98],stage1_12[148],stage1_11[174]}
   );
   gpc615_5 gpc492 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[213]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[38],stage1_13[99],stage1_12[149],stage1_11[175]}
   );
   gpc615_5 gpc493 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[214]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[39],stage1_13[100],stage1_12[150],stage1_11[176]}
   );
   gpc615_5 gpc494 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[215]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[40],stage1_13[101],stage1_12[151],stage1_11[177]}
   );
   gpc615_5 gpc495 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[216]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[41],stage1_13[102],stage1_12[152],stage1_11[178]}
   );
   gpc615_5 gpc496 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[217]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[42],stage1_13[103],stage1_12[153],stage1_11[179]}
   );
   gpc615_5 gpc497 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[218]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[43],stage1_13[104],stage1_12[154],stage1_11[180]}
   );
   gpc615_5 gpc498 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[219]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[44],stage1_13[105],stage1_12[155],stage1_11[181]}
   );
   gpc615_5 gpc499 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[220]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[45],stage1_13[106],stage1_12[156],stage1_11[182]}
   );
   gpc615_5 gpc500 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[221]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[46],stage1_13[107],stage1_12[157],stage1_11[183]}
   );
   gpc615_5 gpc501 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[222]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[47],stage1_13[108],stage1_12[158],stage1_11[184]}
   );
   gpc615_5 gpc502 (
      {stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage0_12[223]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[48],stage1_13[109],stage1_12[159],stage1_11[185]}
   );
   gpc615_5 gpc503 (
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460]},
      {stage0_12[224]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[49],stage1_13[110],stage1_12[160],stage1_11[186]}
   );
   gpc615_5 gpc504 (
      {stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_12[225]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[50],stage1_13[111],stage1_12[161],stage1_11[187]}
   );
   gpc615_5 gpc505 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[226]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[51],stage1_13[112],stage1_12[162],stage1_11[188]}
   );
   gpc615_5 gpc506 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[227]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[52],stage1_13[113],stage1_12[163],stage1_11[189]}
   );
   gpc615_5 gpc507 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[228]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[53],stage1_13[114],stage1_12[164],stage1_11[190]}
   );
   gpc615_5 gpc508 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[229]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[54],stage1_13[115],stage1_12[165],stage1_11[191]}
   );
   gpc615_5 gpc509 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[230]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[55],stage1_13[116],stage1_12[166],stage1_11[192]}
   );
   gpc615_5 gpc510 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[231]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[56],stage1_13[117],stage1_12[167],stage1_11[193]}
   );
   gpc615_5 gpc511 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[232]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[57],stage1_13[118],stage1_12[168],stage1_11[194]}
   );
   gpc606_5 gpc512 (
      {stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[23],stage1_14[58],stage1_13[119],stage1_12[169]}
   );
   gpc606_5 gpc513 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[24],stage1_14[59],stage1_13[120],stage1_12[170]}
   );
   gpc606_5 gpc514 (
      {stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[25],stage1_14[60],stage1_13[121],stage1_12[171]}
   );
   gpc606_5 gpc515 (
      {stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[26],stage1_14[61],stage1_13[122],stage1_12[172]}
   );
   gpc606_5 gpc516 (
      {stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[27],stage1_14[62],stage1_13[123],stage1_12[173]}
   );
   gpc606_5 gpc517 (
      {stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[28],stage1_14[63],stage1_13[124],stage1_12[174]}
   );
   gpc606_5 gpc518 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[29],stage1_14[64],stage1_13[125],stage1_12[175]}
   );
   gpc606_5 gpc519 (
      {stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[30],stage1_14[65],stage1_13[126],stage1_12[176]}
   );
   gpc606_5 gpc520 (
      {stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[31],stage1_14[66],stage1_13[127],stage1_12[177]}
   );
   gpc606_5 gpc521 (
      {stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[32],stage1_14[67],stage1_13[128],stage1_12[178]}
   );
   gpc606_5 gpc522 (
      {stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[33],stage1_14[68],stage1_13[129],stage1_12[179]}
   );
   gpc606_5 gpc523 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[34],stage1_14[69],stage1_13[130],stage1_12[180]}
   );
   gpc606_5 gpc524 (
      {stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[35],stage1_14[70],stage1_13[131],stage1_12[181]}
   );
   gpc606_5 gpc525 (
      {stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[36],stage1_14[71],stage1_13[132],stage1_12[182]}
   );
   gpc615_5 gpc526 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[138]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[37],stage1_14[72],stage1_13[133],stage1_12[183]}
   );
   gpc615_5 gpc527 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[139]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[38],stage1_14[73],stage1_13[134],stage1_12[184]}
   );
   gpc615_5 gpc528 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[140]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[39],stage1_14[74],stage1_13[135],stage1_12[185]}
   );
   gpc615_5 gpc529 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[141]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[40],stage1_14[75],stage1_13[136],stage1_12[186]}
   );
   gpc615_5 gpc530 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[142]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[41],stage1_14[76],stage1_13[137],stage1_12[187]}
   );
   gpc615_5 gpc531 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[143]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[42],stage1_14[77],stage1_13[138],stage1_12[188]}
   );
   gpc615_5 gpc532 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[144]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[43],stage1_14[78],stage1_13[139],stage1_12[189]}
   );
   gpc615_5 gpc533 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[145]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[44],stage1_14[79],stage1_13[140],stage1_12[190]}
   );
   gpc615_5 gpc534 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[146]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[45],stage1_14[80],stage1_13[141],stage1_12[191]}
   );
   gpc615_5 gpc535 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[147]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[46],stage1_14[81],stage1_13[142],stage1_12[192]}
   );
   gpc615_5 gpc536 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[148]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[47],stage1_14[82],stage1_13[143],stage1_12[193]}
   );
   gpc615_5 gpc537 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[149]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[48],stage1_14[83],stage1_13[144],stage1_12[194]}
   );
   gpc615_5 gpc538 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[150]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[49],stage1_14[84],stage1_13[145],stage1_12[195]}
   );
   gpc615_5 gpc539 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[151]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[50],stage1_14[85],stage1_13[146],stage1_12[196]}
   );
   gpc615_5 gpc540 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[152]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[51],stage1_14[86],stage1_13[147],stage1_12[197]}
   );
   gpc615_5 gpc541 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[153]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[52],stage1_14[87],stage1_13[148],stage1_12[198]}
   );
   gpc615_5 gpc542 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[154]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[53],stage1_14[88],stage1_13[149],stage1_12[199]}
   );
   gpc615_5 gpc543 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[155]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[54],stage1_14[89],stage1_13[150],stage1_12[200]}
   );
   gpc615_5 gpc544 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[156]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[55],stage1_14[90],stage1_13[151],stage1_12[201]}
   );
   gpc615_5 gpc545 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[157]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[56],stage1_14[91],stage1_13[152],stage1_12[202]}
   );
   gpc615_5 gpc546 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[158]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[57],stage1_14[92],stage1_13[153],stage1_12[203]}
   );
   gpc615_5 gpc547 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[159]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[58],stage1_14[93],stage1_13[154],stage1_12[204]}
   );
   gpc615_5 gpc548 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[160]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[59],stage1_14[94],stage1_13[155],stage1_12[205]}
   );
   gpc615_5 gpc549 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[161]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[60],stage1_14[95],stage1_13[156],stage1_12[206]}
   );
   gpc615_5 gpc550 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[162]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[61],stage1_14[96],stage1_13[157],stage1_12[207]}
   );
   gpc615_5 gpc551 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[163]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[62],stage1_14[97],stage1_13[158],stage1_12[208]}
   );
   gpc615_5 gpc552 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[164]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[63],stage1_14[98],stage1_13[159],stage1_12[209]}
   );
   gpc615_5 gpc553 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[165]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[64],stage1_14[99],stage1_13[160],stage1_12[210]}
   );
   gpc615_5 gpc554 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[166]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[65],stage1_14[100],stage1_13[161],stage1_12[211]}
   );
   gpc615_5 gpc555 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[167]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[66],stage1_14[101],stage1_13[162],stage1_12[212]}
   );
   gpc615_5 gpc556 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[168]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[67],stage1_14[102],stage1_13[163],stage1_12[213]}
   );
   gpc615_5 gpc557 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[169]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[68],stage1_14[103],stage1_13[164],stage1_12[214]}
   );
   gpc615_5 gpc558 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[170]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[69],stage1_14[104],stage1_13[165],stage1_12[215]}
   );
   gpc615_5 gpc559 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[171]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[70],stage1_14[105],stage1_13[166],stage1_12[216]}
   );
   gpc615_5 gpc560 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[172]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[71],stage1_14[106],stage1_13[167],stage1_12[217]}
   );
   gpc615_5 gpc561 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[173]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[72],stage1_14[107],stage1_13[168],stage1_12[218]}
   );
   gpc615_5 gpc562 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[174]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[73],stage1_14[108],stage1_13[169],stage1_12[219]}
   );
   gpc615_5 gpc563 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[175]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[74],stage1_14[109],stage1_13[170],stage1_12[220]}
   );
   gpc615_5 gpc564 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[176]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[75],stage1_14[110],stage1_13[171],stage1_12[221]}
   );
   gpc606_5 gpc565 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[53],stage1_15[76],stage1_14[111],stage1_13[172]}
   );
   gpc606_5 gpc566 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[54],stage1_15[77],stage1_14[112],stage1_13[173]}
   );
   gpc606_5 gpc567 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[55],stage1_15[78],stage1_14[113],stage1_13[174]}
   );
   gpc606_5 gpc568 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[56],stage1_15[79],stage1_14[114],stage1_13[175]}
   );
   gpc606_5 gpc569 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[57],stage1_15[80],stage1_14[115],stage1_13[176]}
   );
   gpc606_5 gpc570 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[58],stage1_15[81],stage1_14[116],stage1_13[177]}
   );
   gpc606_5 gpc571 (
      {stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[59],stage1_15[82],stage1_14[117],stage1_13[178]}
   );
   gpc606_5 gpc572 (
      {stage0_13[219], stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[60],stage1_15[83],stage1_14[118],stage1_13[179]}
   );
   gpc606_5 gpc573 (
      {stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[61],stage1_15[84],stage1_14[119],stage1_13[180]}
   );
   gpc606_5 gpc574 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[62],stage1_15[85],stage1_14[120],stage1_13[181]}
   );
   gpc606_5 gpc575 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241], stage0_13[242]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[63],stage1_15[86],stage1_14[121],stage1_13[182]}
   );
   gpc606_5 gpc576 (
      {stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246], stage0_13[247], stage0_13[248]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[64],stage1_15[87],stage1_14[122],stage1_13[183]}
   );
   gpc606_5 gpc577 (
      {stage0_13[249], stage0_13[250], stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[65],stage1_15[88],stage1_14[123],stage1_13[184]}
   );
   gpc606_5 gpc578 (
      {stage0_13[255], stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[66],stage1_15[89],stage1_14[124],stage1_13[185]}
   );
   gpc606_5 gpc579 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[67],stage1_15[90],stage1_14[125],stage1_13[186]}
   );
   gpc606_5 gpc580 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271], stage0_13[272]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[68],stage1_15[91],stage1_14[126],stage1_13[187]}
   );
   gpc606_5 gpc581 (
      {stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276], stage0_13[277], stage0_13[278]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[69],stage1_15[92],stage1_14[127],stage1_13[188]}
   );
   gpc606_5 gpc582 (
      {stage0_13[279], stage0_13[280], stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[70],stage1_15[93],stage1_14[128],stage1_13[189]}
   );
   gpc606_5 gpc583 (
      {stage0_13[285], stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[71],stage1_15[94],stage1_14[129],stage1_13[190]}
   );
   gpc606_5 gpc584 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[72],stage1_15[95],stage1_14[130],stage1_13[191]}
   );
   gpc606_5 gpc585 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301], stage0_13[302]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[73],stage1_15[96],stage1_14[131],stage1_13[192]}
   );
   gpc606_5 gpc586 (
      {stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306], stage0_13[307], stage0_13[308]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[74],stage1_15[97],stage1_14[132],stage1_13[193]}
   );
   gpc606_5 gpc587 (
      {stage0_13[309], stage0_13[310], stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[75],stage1_15[98],stage1_14[133],stage1_13[194]}
   );
   gpc606_5 gpc588 (
      {stage0_13[315], stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[76],stage1_15[99],stage1_14[134],stage1_13[195]}
   );
   gpc606_5 gpc589 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[77],stage1_15[100],stage1_14[135],stage1_13[196]}
   );
   gpc606_5 gpc590 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331], stage0_13[332]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[78],stage1_15[101],stage1_14[136],stage1_13[197]}
   );
   gpc606_5 gpc591 (
      {stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336], stage0_13[337], stage0_13[338]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[79],stage1_15[102],stage1_14[137],stage1_13[198]}
   );
   gpc606_5 gpc592 (
      {stage0_13[339], stage0_13[340], stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[80],stage1_15[103],stage1_14[138],stage1_13[199]}
   );
   gpc606_5 gpc593 (
      {stage0_13[345], stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[81],stage1_15[104],stage1_14[139],stage1_13[200]}
   );
   gpc606_5 gpc594 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[82],stage1_15[105],stage1_14[140],stage1_13[201]}
   );
   gpc606_5 gpc595 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361], stage0_13[362]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[83],stage1_15[106],stage1_14[141],stage1_13[202]}
   );
   gpc606_5 gpc596 (
      {stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366], stage0_13[367], stage0_13[368]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[84],stage1_15[107],stage1_14[142],stage1_13[203]}
   );
   gpc606_5 gpc597 (
      {stage0_13[369], stage0_13[370], stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[85],stage1_15[108],stage1_14[143],stage1_13[204]}
   );
   gpc606_5 gpc598 (
      {stage0_13[375], stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[86],stage1_15[109],stage1_14[144],stage1_13[205]}
   );
   gpc606_5 gpc599 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[87],stage1_15[110],stage1_14[145],stage1_13[206]}
   );
   gpc606_5 gpc600 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391], stage0_13[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[88],stage1_15[111],stage1_14[146],stage1_13[207]}
   );
   gpc606_5 gpc601 (
      {stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396], stage0_13[397], stage0_13[398]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[89],stage1_15[112],stage1_14[147],stage1_13[208]}
   );
   gpc606_5 gpc602 (
      {stage0_13[399], stage0_13[400], stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[90],stage1_15[113],stage1_14[148],stage1_13[209]}
   );
   gpc606_5 gpc603 (
      {stage0_13[405], stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[91],stage1_15[114],stage1_14[149],stage1_13[210]}
   );
   gpc606_5 gpc604 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[92],stage1_15[115],stage1_14[150],stage1_13[211]}
   );
   gpc606_5 gpc605 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421], stage0_13[422]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[93],stage1_15[116],stage1_14[151],stage1_13[212]}
   );
   gpc606_5 gpc606 (
      {stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426], stage0_13[427], stage0_13[428]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[94],stage1_15[117],stage1_14[152],stage1_13[213]}
   );
   gpc606_5 gpc607 (
      {stage0_13[429], stage0_13[430], stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[95],stage1_15[118],stage1_14[153],stage1_13[214]}
   );
   gpc606_5 gpc608 (
      {stage0_13[435], stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[96],stage1_15[119],stage1_14[154],stage1_13[215]}
   );
   gpc606_5 gpc609 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[97],stage1_15[120],stage1_14[155],stage1_13[216]}
   );
   gpc606_5 gpc610 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451], stage0_13[452]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[98],stage1_15[121],stage1_14[156],stage1_13[217]}
   );
   gpc606_5 gpc611 (
      {stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456], stage0_13[457], stage0_13[458]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[99],stage1_15[122],stage1_14[157],stage1_13[218]}
   );
   gpc606_5 gpc612 (
      {stage0_13[459], stage0_13[460], stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[100],stage1_15[123],stage1_14[158],stage1_13[219]}
   );
   gpc606_5 gpc613 (
      {stage0_13[465], stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[101],stage1_15[124],stage1_14[159],stage1_13[220]}
   );
   gpc606_5 gpc614 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475], stage0_13[476]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[102],stage1_15[125],stage1_14[160],stage1_13[221]}
   );
   gpc606_5 gpc615 (
      {stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480], stage0_13[481], stage0_13[482]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[103],stage1_15[126],stage1_14[161],stage1_13[222]}
   );
   gpc606_5 gpc616 (
      {stage0_13[483], stage0_13[484], stage0_13[485], stage0_13[486], stage0_13[487], stage0_13[488]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[104],stage1_15[127],stage1_14[162],stage1_13[223]}
   );
   gpc606_5 gpc617 (
      {stage0_13[489], stage0_13[490], stage0_13[491], stage0_13[492], stage0_13[493], stage0_13[494]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[105],stage1_15[128],stage1_14[163],stage1_13[224]}
   );
   gpc606_5 gpc618 (
      {stage0_13[495], stage0_13[496], stage0_13[497], stage0_13[498], stage0_13[499], stage0_13[500]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[106],stage1_15[129],stage1_14[164],stage1_13[225]}
   );
   gpc606_5 gpc619 (
      {stage0_13[501], stage0_13[502], stage0_13[503], stage0_13[504], stage0_13[505], stage0_13[506]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[107],stage1_15[130],stage1_14[165],stage1_13[226]}
   );
   gpc606_5 gpc620 (
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[55],stage1_16[108],stage1_15[131],stage1_14[166]}
   );
   gpc606_5 gpc621 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[56],stage1_16[109],stage1_15[132],stage1_14[167]}
   );
   gpc606_5 gpc622 (
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[57],stage1_16[110],stage1_15[133],stage1_14[168]}
   );
   gpc606_5 gpc623 (
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[58],stage1_16[111],stage1_15[134],stage1_14[169]}
   );
   gpc606_5 gpc624 (
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[59],stage1_16[112],stage1_15[135],stage1_14[170]}
   );
   gpc606_5 gpc625 (
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[60],stage1_16[113],stage1_15[136],stage1_14[171]}
   );
   gpc606_5 gpc626 (
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[61],stage1_16[114],stage1_15[137],stage1_14[172]}
   );
   gpc606_5 gpc627 (
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[62],stage1_16[115],stage1_15[138],stage1_14[173]}
   );
   gpc606_5 gpc628 (
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[63],stage1_16[116],stage1_15[139],stage1_14[174]}
   );
   gpc606_5 gpc629 (
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[64],stage1_16[117],stage1_15[140],stage1_14[175]}
   );
   gpc606_5 gpc630 (
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[65],stage1_16[118],stage1_15[141],stage1_14[176]}
   );
   gpc606_5 gpc631 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[66],stage1_16[119],stage1_15[142],stage1_14[177]}
   );
   gpc606_5 gpc632 (
      {stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[67],stage1_16[120],stage1_15[143],stage1_14[178]}
   );
   gpc606_5 gpc633 (
      {stage0_14[396], stage0_14[397], stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[68],stage1_16[121],stage1_15[144],stage1_14[179]}
   );
   gpc606_5 gpc634 (
      {stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[69],stage1_16[122],stage1_15[145],stage1_14[180]}
   );
   gpc606_5 gpc635 (
      {stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[70],stage1_16[123],stage1_15[146],stage1_14[181]}
   );
   gpc606_5 gpc636 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[71],stage1_16[124],stage1_15[147],stage1_14[182]}
   );
   gpc606_5 gpc637 (
      {stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423], stage0_14[424], stage0_14[425]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[72],stage1_16[125],stage1_15[148],stage1_14[183]}
   );
   gpc606_5 gpc638 (
      {stage0_14[426], stage0_14[427], stage0_14[428], stage0_14[429], stage0_14[430], stage0_14[431]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[73],stage1_16[126],stage1_15[149],stage1_14[184]}
   );
   gpc606_5 gpc639 (
      {stage0_14[432], stage0_14[433], stage0_14[434], stage0_14[435], stage0_14[436], stage0_14[437]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[74],stage1_16[127],stage1_15[150],stage1_14[185]}
   );
   gpc606_5 gpc640 (
      {stage0_14[438], stage0_14[439], stage0_14[440], stage0_14[441], stage0_14[442], stage0_14[443]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[75],stage1_16[128],stage1_15[151],stage1_14[186]}
   );
   gpc606_5 gpc641 (
      {stage0_14[444], stage0_14[445], stage0_14[446], stage0_14[447], stage0_14[448], stage0_14[449]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[76],stage1_16[129],stage1_15[152],stage1_14[187]}
   );
   gpc606_5 gpc642 (
      {stage0_14[450], stage0_14[451], stage0_14[452], stage0_14[453], stage0_14[454], stage0_14[455]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[77],stage1_16[130],stage1_15[153],stage1_14[188]}
   );
   gpc606_5 gpc643 (
      {stage0_14[456], stage0_14[457], stage0_14[458], stage0_14[459], stage0_14[460], stage0_14[461]},
      {stage0_16[138], stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143]},
      {stage1_18[23],stage1_17[78],stage1_16[131],stage1_15[154],stage1_14[189]}
   );
   gpc615_5 gpc644 (
      {stage0_14[462], stage0_14[463], stage0_14[464], stage0_14[465], stage0_14[466]},
      {stage0_15[330]},
      {stage0_16[144], stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149]},
      {stage1_18[24],stage1_17[79],stage1_16[132],stage1_15[155],stage1_14[190]}
   );
   gpc615_5 gpc645 (
      {stage0_14[467], stage0_14[468], stage0_14[469], stage0_14[470], stage0_14[471]},
      {stage0_15[331]},
      {stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155]},
      {stage1_18[25],stage1_17[80],stage1_16[133],stage1_15[156],stage1_14[191]}
   );
   gpc606_5 gpc646 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[26],stage1_17[81],stage1_16[134],stage1_15[157]}
   );
   gpc606_5 gpc647 (
      {stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[27],stage1_17[82],stage1_16[135],stage1_15[158]}
   );
   gpc606_5 gpc648 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[28],stage1_17[83],stage1_16[136],stage1_15[159]}
   );
   gpc606_5 gpc649 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[29],stage1_17[84],stage1_16[137],stage1_15[160]}
   );
   gpc615_5 gpc650 (
      {stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360]},
      {stage0_16[156]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[30],stage1_17[85],stage1_16[138],stage1_15[161]}
   );
   gpc615_5 gpc651 (
      {stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage0_16[157]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[31],stage1_17[86],stage1_16[139],stage1_15[162]}
   );
   gpc615_5 gpc652 (
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370]},
      {stage0_16[158]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[32],stage1_17[87],stage1_16[140],stage1_15[163]}
   );
   gpc615_5 gpc653 (
      {stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375]},
      {stage0_16[159]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[33],stage1_17[88],stage1_16[141],stage1_15[164]}
   );
   gpc615_5 gpc654 (
      {stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380]},
      {stage0_16[160]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[34],stage1_17[89],stage1_16[142],stage1_15[165]}
   );
   gpc615_5 gpc655 (
      {stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385]},
      {stage0_16[161]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[35],stage1_17[90],stage1_16[143],stage1_15[166]}
   );
   gpc615_5 gpc656 (
      {stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390]},
      {stage0_16[162]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[36],stage1_17[91],stage1_16[144],stage1_15[167]}
   );
   gpc615_5 gpc657 (
      {stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage0_16[163]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[37],stage1_17[92],stage1_16[145],stage1_15[168]}
   );
   gpc615_5 gpc658 (
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400]},
      {stage0_16[164]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[38],stage1_17[93],stage1_16[146],stage1_15[169]}
   );
   gpc615_5 gpc659 (
      {stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405]},
      {stage0_16[165]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[39],stage1_17[94],stage1_16[147],stage1_15[170]}
   );
   gpc615_5 gpc660 (
      {stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410]},
      {stage0_16[166]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[40],stage1_17[95],stage1_16[148],stage1_15[171]}
   );
   gpc615_5 gpc661 (
      {stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415]},
      {stage0_16[167]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[41],stage1_17[96],stage1_16[149],stage1_15[172]}
   );
   gpc615_5 gpc662 (
      {stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420]},
      {stage0_16[168]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[42],stage1_17[97],stage1_16[150],stage1_15[173]}
   );
   gpc615_5 gpc663 (
      {stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage0_16[169]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[43],stage1_17[98],stage1_16[151],stage1_15[174]}
   );
   gpc615_5 gpc664 (
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430]},
      {stage0_16[170]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[44],stage1_17[99],stage1_16[152],stage1_15[175]}
   );
   gpc615_5 gpc665 (
      {stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435]},
      {stage0_16[171]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[45],stage1_17[100],stage1_16[153],stage1_15[176]}
   );
   gpc615_5 gpc666 (
      {stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440]},
      {stage0_16[172]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[46],stage1_17[101],stage1_16[154],stage1_15[177]}
   );
   gpc615_5 gpc667 (
      {stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445]},
      {stage0_16[173]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[47],stage1_17[102],stage1_16[155],stage1_15[178]}
   );
   gpc615_5 gpc668 (
      {stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450]},
      {stage0_16[174]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[48],stage1_17[103],stage1_16[156],stage1_15[179]}
   );
   gpc615_5 gpc669 (
      {stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage0_16[175]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[49],stage1_17[104],stage1_16[157],stage1_15[180]}
   );
   gpc606_5 gpc670 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[24],stage1_18[50],stage1_17[105],stage1_16[158]}
   );
   gpc606_5 gpc671 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[25],stage1_18[51],stage1_17[106],stage1_16[159]}
   );
   gpc606_5 gpc672 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[26],stage1_18[52],stage1_17[107],stage1_16[160]}
   );
   gpc606_5 gpc673 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[27],stage1_18[53],stage1_17[108],stage1_16[161]}
   );
   gpc606_5 gpc674 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[28],stage1_18[54],stage1_17[109],stage1_16[162]}
   );
   gpc606_5 gpc675 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[29],stage1_18[55],stage1_17[110],stage1_16[163]}
   );
   gpc606_5 gpc676 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[30],stage1_18[56],stage1_17[111],stage1_16[164]}
   );
   gpc606_5 gpc677 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[31],stage1_18[57],stage1_17[112],stage1_16[165]}
   );
   gpc606_5 gpc678 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[32],stage1_18[58],stage1_17[113],stage1_16[166]}
   );
   gpc606_5 gpc679 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[33],stage1_18[59],stage1_17[114],stage1_16[167]}
   );
   gpc606_5 gpc680 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[34],stage1_18[60],stage1_17[115],stage1_16[168]}
   );
   gpc606_5 gpc681 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[35],stage1_18[61],stage1_17[116],stage1_16[169]}
   );
   gpc606_5 gpc682 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[36],stage1_18[62],stage1_17[117],stage1_16[170]}
   );
   gpc606_5 gpc683 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[37],stage1_18[63],stage1_17[118],stage1_16[171]}
   );
   gpc606_5 gpc684 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[38],stage1_18[64],stage1_17[119],stage1_16[172]}
   );
   gpc606_5 gpc685 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[39],stage1_18[65],stage1_17[120],stage1_16[173]}
   );
   gpc606_5 gpc686 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[40],stage1_18[66],stage1_17[121],stage1_16[174]}
   );
   gpc606_5 gpc687 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[41],stage1_18[67],stage1_17[122],stage1_16[175]}
   );
   gpc606_5 gpc688 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[42],stage1_18[68],stage1_17[123],stage1_16[176]}
   );
   gpc606_5 gpc689 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[43],stage1_18[69],stage1_17[124],stage1_16[177]}
   );
   gpc606_5 gpc690 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[44],stage1_18[70],stage1_17[125],stage1_16[178]}
   );
   gpc606_5 gpc691 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[45],stage1_18[71],stage1_17[126],stage1_16[179]}
   );
   gpc606_5 gpc692 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[46],stage1_18[72],stage1_17[127],stage1_16[180]}
   );
   gpc606_5 gpc693 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[47],stage1_18[73],stage1_17[128],stage1_16[181]}
   );
   gpc606_5 gpc694 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[48],stage1_18[74],stage1_17[129],stage1_16[182]}
   );
   gpc606_5 gpc695 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[49],stage1_18[75],stage1_17[130],stage1_16[183]}
   );
   gpc606_5 gpc696 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[50],stage1_18[76],stage1_17[131],stage1_16[184]}
   );
   gpc606_5 gpc697 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[51],stage1_18[77],stage1_17[132],stage1_16[185]}
   );
   gpc606_5 gpc698 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[52],stage1_18[78],stage1_17[133],stage1_16[186]}
   );
   gpc606_5 gpc699 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[53],stage1_18[79],stage1_17[134],stage1_16[187]}
   );
   gpc606_5 gpc700 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[54],stage1_18[80],stage1_17[135],stage1_16[188]}
   );
   gpc606_5 gpc701 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[55],stage1_18[81],stage1_17[136],stage1_16[189]}
   );
   gpc606_5 gpc702 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[56],stage1_18[82],stage1_17[137],stage1_16[190]}
   );
   gpc606_5 gpc703 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[57],stage1_18[83],stage1_17[138],stage1_16[191]}
   );
   gpc606_5 gpc704 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[58],stage1_18[84],stage1_17[139],stage1_16[192]}
   );
   gpc606_5 gpc705 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[59],stage1_18[85],stage1_17[140],stage1_16[193]}
   );
   gpc606_5 gpc706 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[60],stage1_18[86],stage1_17[141],stage1_16[194]}
   );
   gpc606_5 gpc707 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[61],stage1_18[87],stage1_17[142],stage1_16[195]}
   );
   gpc606_5 gpc708 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[62],stage1_18[88],stage1_17[143],stage1_16[196]}
   );
   gpc606_5 gpc709 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[63],stage1_18[89],stage1_17[144],stage1_16[197]}
   );
   gpc606_5 gpc710 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[64],stage1_18[90],stage1_17[145],stage1_16[198]}
   );
   gpc606_5 gpc711 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[65],stage1_18[91],stage1_17[146],stage1_16[199]}
   );
   gpc606_5 gpc712 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[66],stage1_18[92],stage1_17[147],stage1_16[200]}
   );
   gpc606_5 gpc713 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[67],stage1_18[93],stage1_17[148],stage1_16[201]}
   );
   gpc606_5 gpc714 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[68],stage1_18[94],stage1_17[149],stage1_16[202]}
   );
   gpc606_5 gpc715 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[69],stage1_18[95],stage1_17[150],stage1_16[203]}
   );
   gpc606_5 gpc716 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[70],stage1_18[96],stage1_17[151],stage1_16[204]}
   );
   gpc606_5 gpc717 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[71],stage1_18[97],stage1_17[152],stage1_16[205]}
   );
   gpc606_5 gpc718 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[72],stage1_18[98],stage1_17[153],stage1_16[206]}
   );
   gpc606_5 gpc719 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[73],stage1_18[99],stage1_17[154],stage1_16[207]}
   );
   gpc606_5 gpc720 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[74],stage1_18[100],stage1_17[155],stage1_16[208]}
   );
   gpc606_5 gpc721 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[75],stage1_18[101],stage1_17[156],stage1_16[209]}
   );
   gpc606_5 gpc722 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[76],stage1_18[102],stage1_17[157],stage1_16[210]}
   );
   gpc606_5 gpc723 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[77],stage1_18[103],stage1_17[158],stage1_16[211]}
   );
   gpc606_5 gpc724 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[78],stage1_18[104],stage1_17[159],stage1_16[212]}
   );
   gpc606_5 gpc725 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[79],stage1_18[105],stage1_17[160],stage1_16[213]}
   );
   gpc606_5 gpc726 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[56],stage1_19[80],stage1_18[106],stage1_17[161]}
   );
   gpc606_5 gpc727 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[57],stage1_19[81],stage1_18[107],stage1_17[162]}
   );
   gpc606_5 gpc728 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[58],stage1_19[82],stage1_18[108],stage1_17[163]}
   );
   gpc606_5 gpc729 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[59],stage1_19[83],stage1_18[109],stage1_17[164]}
   );
   gpc606_5 gpc730 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[60],stage1_19[84],stage1_18[110],stage1_17[165]}
   );
   gpc606_5 gpc731 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[61],stage1_19[85],stage1_18[111],stage1_17[166]}
   );
   gpc606_5 gpc732 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[62],stage1_19[86],stage1_18[112],stage1_17[167]}
   );
   gpc606_5 gpc733 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[63],stage1_19[87],stage1_18[113],stage1_17[168]}
   );
   gpc606_5 gpc734 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[64],stage1_19[88],stage1_18[114],stage1_17[169]}
   );
   gpc606_5 gpc735 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[65],stage1_19[89],stage1_18[115],stage1_17[170]}
   );
   gpc606_5 gpc736 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[66],stage1_19[90],stage1_18[116],stage1_17[171]}
   );
   gpc606_5 gpc737 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[67],stage1_19[91],stage1_18[117],stage1_17[172]}
   );
   gpc606_5 gpc738 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[68],stage1_19[92],stage1_18[118],stage1_17[173]}
   );
   gpc606_5 gpc739 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[69],stage1_19[93],stage1_18[119],stage1_17[174]}
   );
   gpc606_5 gpc740 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[70],stage1_19[94],stage1_18[120],stage1_17[175]}
   );
   gpc606_5 gpc741 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[71],stage1_19[95],stage1_18[121],stage1_17[176]}
   );
   gpc606_5 gpc742 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[72],stage1_19[96],stage1_18[122],stage1_17[177]}
   );
   gpc606_5 gpc743 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[73],stage1_19[97],stage1_18[123],stage1_17[178]}
   );
   gpc606_5 gpc744 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[74],stage1_19[98],stage1_18[124],stage1_17[179]}
   );
   gpc606_5 gpc745 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[75],stage1_19[99],stage1_18[125],stage1_17[180]}
   );
   gpc606_5 gpc746 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[76],stage1_19[100],stage1_18[126],stage1_17[181]}
   );
   gpc606_5 gpc747 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[77],stage1_19[101],stage1_18[127],stage1_17[182]}
   );
   gpc606_5 gpc748 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[78],stage1_19[102],stage1_18[128],stage1_17[183]}
   );
   gpc606_5 gpc749 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[79],stage1_19[103],stage1_18[129],stage1_17[184]}
   );
   gpc606_5 gpc750 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[80],stage1_19[104],stage1_18[130],stage1_17[185]}
   );
   gpc606_5 gpc751 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[81],stage1_19[105],stage1_18[131],stage1_17[186]}
   );
   gpc606_5 gpc752 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[82],stage1_19[106],stage1_18[132],stage1_17[187]}
   );
   gpc606_5 gpc753 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[83],stage1_19[107],stage1_18[133],stage1_17[188]}
   );
   gpc606_5 gpc754 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[84],stage1_19[108],stage1_18[134],stage1_17[189]}
   );
   gpc606_5 gpc755 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[85],stage1_19[109],stage1_18[135],stage1_17[190]}
   );
   gpc606_5 gpc756 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[86],stage1_19[110],stage1_18[136],stage1_17[191]}
   );
   gpc606_5 gpc757 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[87],stage1_19[111],stage1_18[137],stage1_17[192]}
   );
   gpc606_5 gpc758 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[88],stage1_19[112],stage1_18[138],stage1_17[193]}
   );
   gpc606_5 gpc759 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[89],stage1_19[113],stage1_18[139],stage1_17[194]}
   );
   gpc606_5 gpc760 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[90],stage1_19[114],stage1_18[140],stage1_17[195]}
   );
   gpc606_5 gpc761 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[91],stage1_19[115],stage1_18[141],stage1_17[196]}
   );
   gpc606_5 gpc762 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[92],stage1_19[116],stage1_18[142],stage1_17[197]}
   );
   gpc606_5 gpc763 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[93],stage1_19[117],stage1_18[143],stage1_17[198]}
   );
   gpc606_5 gpc764 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[94],stage1_19[118],stage1_18[144],stage1_17[199]}
   );
   gpc606_5 gpc765 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[95],stage1_19[119],stage1_18[145],stage1_17[200]}
   );
   gpc606_5 gpc766 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[240], stage0_19[241], stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245]},
      {stage1_21[40],stage1_20[96],stage1_19[120],stage1_18[146],stage1_17[201]}
   );
   gpc606_5 gpc767 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[246], stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage1_21[41],stage1_20[97],stage1_19[121],stage1_18[147],stage1_17[202]}
   );
   gpc606_5 gpc768 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256], stage0_19[257]},
      {stage1_21[42],stage1_20[98],stage1_19[122],stage1_18[148],stage1_17[203]}
   );
   gpc606_5 gpc769 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261], stage0_19[262], stage0_19[263]},
      {stage1_21[43],stage1_20[99],stage1_19[123],stage1_18[149],stage1_17[204]}
   );
   gpc606_5 gpc770 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[264], stage0_19[265], stage0_19[266], stage0_19[267], stage0_19[268], stage0_19[269]},
      {stage1_21[44],stage1_20[100],stage1_19[124],stage1_18[150],stage1_17[205]}
   );
   gpc606_5 gpc771 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[270], stage0_19[271], stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275]},
      {stage1_21[45],stage1_20[101],stage1_19[125],stage1_18[151],stage1_17[206]}
   );
   gpc606_5 gpc772 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[276], stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage1_21[46],stage1_20[102],stage1_19[126],stage1_18[152],stage1_17[207]}
   );
   gpc606_5 gpc773 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286], stage0_19[287]},
      {stage1_21[47],stage1_20[103],stage1_19[127],stage1_18[153],stage1_17[208]}
   );
   gpc606_5 gpc774 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291], stage0_19[292], stage0_19[293]},
      {stage1_21[48],stage1_20[104],stage1_19[128],stage1_18[154],stage1_17[209]}
   );
   gpc606_5 gpc775 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[294], stage0_19[295], stage0_19[296], stage0_19[297], stage0_19[298], stage0_19[299]},
      {stage1_21[49],stage1_20[105],stage1_19[129],stage1_18[155],stage1_17[210]}
   );
   gpc606_5 gpc776 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[300], stage0_19[301], stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305]},
      {stage1_21[50],stage1_20[106],stage1_19[130],stage1_18[156],stage1_17[211]}
   );
   gpc606_5 gpc777 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[306], stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage1_21[51],stage1_20[107],stage1_19[131],stage1_18[157],stage1_17[212]}
   );
   gpc606_5 gpc778 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316], stage0_19[317]},
      {stage1_21[52],stage1_20[108],stage1_19[132],stage1_18[158],stage1_17[213]}
   );
   gpc606_5 gpc779 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321], stage0_19[322], stage0_19[323]},
      {stage1_21[53],stage1_20[109],stage1_19[133],stage1_18[159],stage1_17[214]}
   );
   gpc606_5 gpc780 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[324], stage0_19[325], stage0_19[326], stage0_19[327], stage0_19[328], stage0_19[329]},
      {stage1_21[54],stage1_20[110],stage1_19[134],stage1_18[160],stage1_17[215]}
   );
   gpc606_5 gpc781 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[330], stage0_19[331], stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335]},
      {stage1_21[55],stage1_20[111],stage1_19[135],stage1_18[161],stage1_17[216]}
   );
   gpc606_5 gpc782 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[336], stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage1_21[56],stage1_20[112],stage1_19[136],stage1_18[162],stage1_17[217]}
   );
   gpc606_5 gpc783 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346], stage0_19[347]},
      {stage1_21[57],stage1_20[113],stage1_19[137],stage1_18[163],stage1_17[218]}
   );
   gpc606_5 gpc784 (
      {stage0_17[492], stage0_17[493], stage0_17[494], stage0_17[495], stage0_17[496], stage0_17[497]},
      {stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351], stage0_19[352], stage0_19[353]},
      {stage1_21[58],stage1_20[114],stage1_19[138],stage1_18[164],stage1_17[219]}
   );
   gpc606_5 gpc785 (
      {stage0_17[498], stage0_17[499], stage0_17[500], stage0_17[501], stage0_17[502], stage0_17[503]},
      {stage0_19[354], stage0_19[355], stage0_19[356], stage0_19[357], stage0_19[358], stage0_19[359]},
      {stage1_21[59],stage1_20[115],stage1_19[139],stage1_18[165],stage1_17[220]}
   );
   gpc606_5 gpc786 (
      {stage0_17[504], stage0_17[505], stage0_17[506], stage0_17[507], stage0_17[508], stage0_17[509]},
      {stage0_19[360], stage0_19[361], stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365]},
      {stage1_21[60],stage1_20[116],stage1_19[140],stage1_18[166],stage1_17[221]}
   );
   gpc615_5 gpc787 (
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340]},
      {stage0_19[366]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[61],stage1_20[117],stage1_19[141],stage1_18[167]}
   );
   gpc615_5 gpc788 (
      {stage0_18[341], stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345]},
      {stage0_19[367]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[62],stage1_20[118],stage1_19[142],stage1_18[168]}
   );
   gpc615_5 gpc789 (
      {stage0_18[346], stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350]},
      {stage0_19[368]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[63],stage1_20[119],stage1_19[143],stage1_18[169]}
   );
   gpc615_5 gpc790 (
      {stage0_18[351], stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355]},
      {stage0_19[369]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[64],stage1_20[120],stage1_19[144],stage1_18[170]}
   );
   gpc615_5 gpc791 (
      {stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360]},
      {stage0_19[370]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[65],stage1_20[121],stage1_19[145],stage1_18[171]}
   );
   gpc615_5 gpc792 (
      {stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage0_19[371]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[66],stage1_20[122],stage1_19[146],stage1_18[172]}
   );
   gpc615_5 gpc793 (
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370]},
      {stage0_19[372]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[67],stage1_20[123],stage1_19[147],stage1_18[173]}
   );
   gpc615_5 gpc794 (
      {stage0_18[371], stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375]},
      {stage0_19[373]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[68],stage1_20[124],stage1_19[148],stage1_18[174]}
   );
   gpc615_5 gpc795 (
      {stage0_18[376], stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380]},
      {stage0_19[374]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[69],stage1_20[125],stage1_19[149],stage1_18[175]}
   );
   gpc615_5 gpc796 (
      {stage0_18[381], stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385]},
      {stage0_19[375]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[70],stage1_20[126],stage1_19[150],stage1_18[176]}
   );
   gpc615_5 gpc797 (
      {stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390]},
      {stage0_19[376]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[71],stage1_20[127],stage1_19[151],stage1_18[177]}
   );
   gpc615_5 gpc798 (
      {stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage0_19[377]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[72],stage1_20[128],stage1_19[152],stage1_18[178]}
   );
   gpc615_5 gpc799 (
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400]},
      {stage0_19[378]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[73],stage1_20[129],stage1_19[153],stage1_18[179]}
   );
   gpc615_5 gpc800 (
      {stage0_18[401], stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405]},
      {stage0_19[379]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[74],stage1_20[130],stage1_19[154],stage1_18[180]}
   );
   gpc615_5 gpc801 (
      {stage0_18[406], stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410]},
      {stage0_19[380]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[75],stage1_20[131],stage1_19[155],stage1_18[181]}
   );
   gpc615_5 gpc802 (
      {stage0_18[411], stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415]},
      {stage0_19[381]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[76],stage1_20[132],stage1_19[156],stage1_18[182]}
   );
   gpc615_5 gpc803 (
      {stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420]},
      {stage0_19[382]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[77],stage1_20[133],stage1_19[157],stage1_18[183]}
   );
   gpc615_5 gpc804 (
      {stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage0_19[383]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[78],stage1_20[134],stage1_19[158],stage1_18[184]}
   );
   gpc615_5 gpc805 (
      {stage0_18[426], stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430]},
      {stage0_19[384]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[79],stage1_20[135],stage1_19[159],stage1_18[185]}
   );
   gpc615_5 gpc806 (
      {stage0_18[431], stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435]},
      {stage0_19[385]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[80],stage1_20[136],stage1_19[160],stage1_18[186]}
   );
   gpc615_5 gpc807 (
      {stage0_18[436], stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440]},
      {stage0_19[386]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[81],stage1_20[137],stage1_19[161],stage1_18[187]}
   );
   gpc615_5 gpc808 (
      {stage0_18[441], stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445]},
      {stage0_19[387]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[82],stage1_20[138],stage1_19[162],stage1_18[188]}
   );
   gpc615_5 gpc809 (
      {stage0_18[446], stage0_18[447], stage0_18[448], stage0_18[449], stage0_18[450]},
      {stage0_19[388]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[83],stage1_20[139],stage1_19[163],stage1_18[189]}
   );
   gpc615_5 gpc810 (
      {stage0_18[451], stage0_18[452], stage0_18[453], stage0_18[454], stage0_18[455]},
      {stage0_19[389]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[84],stage1_20[140],stage1_19[164],stage1_18[190]}
   );
   gpc615_5 gpc811 (
      {stage0_18[456], stage0_18[457], stage0_18[458], stage0_18[459], stage0_18[460]},
      {stage0_19[390]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[85],stage1_20[141],stage1_19[165],stage1_18[191]}
   );
   gpc615_5 gpc812 (
      {stage0_18[461], stage0_18[462], stage0_18[463], stage0_18[464], stage0_18[465]},
      {stage0_19[391]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[86],stage1_20[142],stage1_19[166],stage1_18[192]}
   );
   gpc615_5 gpc813 (
      {stage0_18[466], stage0_18[467], stage0_18[468], stage0_18[469], stage0_18[470]},
      {stage0_19[392]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[87],stage1_20[143],stage1_19[167],stage1_18[193]}
   );
   gpc615_5 gpc814 (
      {stage0_18[471], stage0_18[472], stage0_18[473], stage0_18[474], stage0_18[475]},
      {stage0_19[393]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[88],stage1_20[144],stage1_19[168],stage1_18[194]}
   );
   gpc615_5 gpc815 (
      {stage0_18[476], stage0_18[477], stage0_18[478], stage0_18[479], stage0_18[480]},
      {stage0_19[394]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[89],stage1_20[145],stage1_19[169],stage1_18[195]}
   );
   gpc615_5 gpc816 (
      {stage0_18[481], stage0_18[482], stage0_18[483], stage0_18[484], stage0_18[485]},
      {stage0_19[395]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[90],stage1_20[146],stage1_19[170],stage1_18[196]}
   );
   gpc615_5 gpc817 (
      {stage0_18[486], stage0_18[487], stage0_18[488], stage0_18[489], stage0_18[490]},
      {stage0_19[396]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[91],stage1_20[147],stage1_19[171],stage1_18[197]}
   );
   gpc615_5 gpc818 (
      {stage0_18[491], stage0_18[492], stage0_18[493], stage0_18[494], stage0_18[495]},
      {stage0_19[397]},
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage1_22[31],stage1_21[92],stage1_20[148],stage1_19[172],stage1_18[198]}
   );
   gpc615_5 gpc819 (
      {stage0_18[496], stage0_18[497], stage0_18[498], stage0_18[499], stage0_18[500]},
      {stage0_19[398]},
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage1_22[32],stage1_21[93],stage1_20[149],stage1_19[173],stage1_18[199]}
   );
   gpc615_5 gpc820 (
      {stage0_18[501], stage0_18[502], stage0_18[503], stage0_18[504], stage0_18[505]},
      {stage0_19[399]},
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage1_22[33],stage1_21[94],stage1_20[150],stage1_19[174],stage1_18[200]}
   );
   gpc615_5 gpc821 (
      {stage0_18[506], stage0_18[507], stage0_18[508], stage0_18[509], stage0_18[510]},
      {stage0_19[400]},
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage1_22[34],stage1_21[95],stage1_20[151],stage1_19[175],stage1_18[201]}
   );
   gpc615_5 gpc822 (
      {stage0_19[401], stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405]},
      {stage0_20[210]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[35],stage1_21[96],stage1_20[152],stage1_19[176]}
   );
   gpc615_5 gpc823 (
      {stage0_19[406], stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410]},
      {stage0_20[211]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[36],stage1_21[97],stage1_20[153],stage1_19[177]}
   );
   gpc615_5 gpc824 (
      {stage0_19[411], stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415]},
      {stage0_20[212]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[37],stage1_21[98],stage1_20[154],stage1_19[178]}
   );
   gpc615_5 gpc825 (
      {stage0_19[416], stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420]},
      {stage0_20[213]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[38],stage1_21[99],stage1_20[155],stage1_19[179]}
   );
   gpc615_5 gpc826 (
      {stage0_19[421], stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425]},
      {stage0_20[214]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[39],stage1_21[100],stage1_20[156],stage1_19[180]}
   );
   gpc615_5 gpc827 (
      {stage0_19[426], stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430]},
      {stage0_20[215]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[40],stage1_21[101],stage1_20[157],stage1_19[181]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[6],stage1_22[41],stage1_21[102],stage1_20[158]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[7],stage1_22[42],stage1_21[103],stage1_20[159]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[8],stage1_22[43],stage1_21[104],stage1_20[160]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[9],stage1_22[44],stage1_21[105],stage1_20[161]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[10],stage1_22[45],stage1_21[106],stage1_20[162]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[11],stage1_22[46],stage1_21[107],stage1_20[163]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[12],stage1_22[47],stage1_21[108],stage1_20[164]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[13],stage1_22[48],stage1_21[109],stage1_20[165]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[14],stage1_22[49],stage1_21[110],stage1_20[166]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[15],stage1_22[50],stage1_21[111],stage1_20[167]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[16],stage1_22[51],stage1_21[112],stage1_20[168]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[17],stage1_22[52],stage1_21[113],stage1_20[169]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[18],stage1_22[53],stage1_21[114],stage1_20[170]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[19],stage1_22[54],stage1_21[115],stage1_20[171]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[20],stage1_22[55],stage1_21[116],stage1_20[172]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[21],stage1_22[56],stage1_21[117],stage1_20[173]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[22],stage1_22[57],stage1_21[118],stage1_20[174]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[23],stage1_22[58],stage1_21[119],stage1_20[175]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[24],stage1_22[59],stage1_21[120],stage1_20[176]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[25],stage1_22[60],stage1_21[121],stage1_20[177]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[26],stage1_22[61],stage1_21[122],stage1_20[178]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[27],stage1_22[62],stage1_21[123],stage1_20[179]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[28],stage1_22[63],stage1_21[124],stage1_20[180]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[29],stage1_22[64],stage1_21[125],stage1_20[181]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[30],stage1_22[65],stage1_21[126],stage1_20[182]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[31],stage1_22[66],stage1_21[127],stage1_20[183]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[32],stage1_22[67],stage1_21[128],stage1_20[184]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[33],stage1_22[68],stage1_21[129],stage1_20[185]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[34],stage1_22[69],stage1_21[130],stage1_20[186]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[35],stage1_22[70],stage1_21[131],stage1_20[187]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[36],stage1_22[71],stage1_21[132],stage1_20[188]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[37],stage1_22[72],stage1_21[133],stage1_20[189]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[38],stage1_22[73],stage1_21[134],stage1_20[190]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[39],stage1_22[74],stage1_21[135],stage1_20[191]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[40],stage1_22[75],stage1_21[136],stage1_20[192]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[41],stage1_22[76],stage1_21[137],stage1_20[193]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[42],stage1_22[77],stage1_21[138],stage1_20[194]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[43],stage1_22[78],stage1_21[139],stage1_20[195]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[44],stage1_22[79],stage1_21[140],stage1_20[196]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[45],stage1_22[80],stage1_21[141],stage1_20[197]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[46],stage1_22[81],stage1_21[142],stage1_20[198]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[47],stage1_22[82],stage1_21[143],stage1_20[199]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[48],stage1_22[83],stage1_21[144],stage1_20[200]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[49],stage1_22[84],stage1_21[145],stage1_20[201]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[50],stage1_22[85],stage1_21[146],stage1_20[202]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[51],stage1_22[86],stage1_21[147],stage1_20[203]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[52],stage1_22[87],stage1_21[148],stage1_20[204]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[53],stage1_22[88],stage1_21[149],stage1_20[205]}
   );
   gpc606_5 gpc876 (
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[48],stage1_23[54],stage1_22[89],stage1_21[150]}
   );
   gpc606_5 gpc877 (
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[49],stage1_23[55],stage1_22[90],stage1_21[151]}
   );
   gpc606_5 gpc878 (
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[50],stage1_23[56],stage1_22[91],stage1_21[152]}
   );
   gpc606_5 gpc879 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[51],stage1_23[57],stage1_22[92],stage1_21[153]}
   );
   gpc606_5 gpc880 (
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[52],stage1_23[58],stage1_22[93],stage1_21[154]}
   );
   gpc606_5 gpc881 (
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[53],stage1_23[59],stage1_22[94],stage1_21[155]}
   );
   gpc606_5 gpc882 (
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[54],stage1_23[60],stage1_22[95],stage1_21[156]}
   );
   gpc606_5 gpc883 (
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[55],stage1_23[61],stage1_22[96],stage1_21[157]}
   );
   gpc606_5 gpc884 (
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[56],stage1_23[62],stage1_22[97],stage1_21[158]}
   );
   gpc606_5 gpc885 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[57],stage1_23[63],stage1_22[98],stage1_21[159]}
   );
   gpc606_5 gpc886 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[58],stage1_23[64],stage1_22[99],stage1_21[160]}
   );
   gpc606_5 gpc887 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[59],stage1_23[65],stage1_22[100],stage1_21[161]}
   );
   gpc606_5 gpc888 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[60],stage1_23[66],stage1_22[101],stage1_21[162]}
   );
   gpc606_5 gpc889 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[61],stage1_23[67],stage1_22[102],stage1_21[163]}
   );
   gpc606_5 gpc890 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[62],stage1_23[68],stage1_22[103],stage1_21[164]}
   );
   gpc606_5 gpc891 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[63],stage1_23[69],stage1_22[104],stage1_21[165]}
   );
   gpc606_5 gpc892 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[64],stage1_23[70],stage1_22[105],stage1_21[166]}
   );
   gpc606_5 gpc893 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[65],stage1_23[71],stage1_22[106],stage1_21[167]}
   );
   gpc606_5 gpc894 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[66],stage1_23[72],stage1_22[107],stage1_21[168]}
   );
   gpc606_5 gpc895 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[67],stage1_23[73],stage1_22[108],stage1_21[169]}
   );
   gpc606_5 gpc896 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[68],stage1_23[74],stage1_22[109],stage1_21[170]}
   );
   gpc606_5 gpc897 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[69],stage1_23[75],stage1_22[110],stage1_21[171]}
   );
   gpc606_5 gpc898 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[70],stage1_23[76],stage1_22[111],stage1_21[172]}
   );
   gpc606_5 gpc899 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[71],stage1_23[77],stage1_22[112],stage1_21[173]}
   );
   gpc606_5 gpc900 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[72],stage1_23[78],stage1_22[113],stage1_21[174]}
   );
   gpc606_5 gpc901 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[73],stage1_23[79],stage1_22[114],stage1_21[175]}
   );
   gpc606_5 gpc902 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[74],stage1_23[80],stage1_22[115],stage1_21[176]}
   );
   gpc606_5 gpc903 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[75],stage1_23[81],stage1_22[116],stage1_21[177]}
   );
   gpc606_5 gpc904 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[76],stage1_23[82],stage1_22[117],stage1_21[178]}
   );
   gpc606_5 gpc905 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[77],stage1_23[83],stage1_22[118],stage1_21[179]}
   );
   gpc606_5 gpc906 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[78],stage1_23[84],stage1_22[119],stage1_21[180]}
   );
   gpc606_5 gpc907 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[79],stage1_23[85],stage1_22[120],stage1_21[181]}
   );
   gpc606_5 gpc908 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[80],stage1_23[86],stage1_22[121],stage1_21[182]}
   );
   gpc606_5 gpc909 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[81],stage1_23[87],stage1_22[122],stage1_21[183]}
   );
   gpc606_5 gpc910 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[82],stage1_23[88],stage1_22[123],stage1_21[184]}
   );
   gpc606_5 gpc911 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[83],stage1_23[89],stage1_22[124],stage1_21[185]}
   );
   gpc606_5 gpc912 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[84],stage1_23[90],stage1_22[125],stage1_21[186]}
   );
   gpc606_5 gpc913 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[85],stage1_23[91],stage1_22[126],stage1_21[187]}
   );
   gpc606_5 gpc914 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[86],stage1_23[92],stage1_22[127],stage1_21[188]}
   );
   gpc606_5 gpc915 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[87],stage1_23[93],stage1_22[128],stage1_21[189]}
   );
   gpc615_5 gpc916 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280]},
      {stage0_22[288]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[88],stage1_23[94],stage1_22[129],stage1_21[190]}
   );
   gpc615_5 gpc917 (
      {stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[289]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[89],stage1_23[95],stage1_22[130],stage1_21[191]}
   );
   gpc615_5 gpc918 (
      {stage0_21[286], stage0_21[287], stage0_21[288], stage0_21[289], stage0_21[290]},
      {stage0_22[290]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[90],stage1_23[96],stage1_22[131],stage1_21[192]}
   );
   gpc615_5 gpc919 (
      {stage0_21[291], stage0_21[292], stage0_21[293], stage0_21[294], stage0_21[295]},
      {stage0_22[291]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[91],stage1_23[97],stage1_22[132],stage1_21[193]}
   );
   gpc615_5 gpc920 (
      {stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299], stage0_21[300]},
      {stage0_22[292]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[92],stage1_23[98],stage1_22[133],stage1_21[194]}
   );
   gpc615_5 gpc921 (
      {stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_22[293]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[93],stage1_23[99],stage1_22[134],stage1_21[195]}
   );
   gpc615_5 gpc922 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310]},
      {stage0_22[294]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[94],stage1_23[100],stage1_22[135],stage1_21[196]}
   );
   gpc615_5 gpc923 (
      {stage0_21[311], stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315]},
      {stage0_22[295]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[95],stage1_23[101],stage1_22[136],stage1_21[197]}
   );
   gpc615_5 gpc924 (
      {stage0_21[316], stage0_21[317], stage0_21[318], stage0_21[319], stage0_21[320]},
      {stage0_22[296]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[96],stage1_23[102],stage1_22[137],stage1_21[198]}
   );
   gpc615_5 gpc925 (
      {stage0_21[321], stage0_21[322], stage0_21[323], stage0_21[324], stage0_21[325]},
      {stage0_22[297]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[97],stage1_23[103],stage1_22[138],stage1_21[199]}
   );
   gpc615_5 gpc926 (
      {stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329], stage0_21[330]},
      {stage0_22[298]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[98],stage1_23[104],stage1_22[139],stage1_21[200]}
   );
   gpc615_5 gpc927 (
      {stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_22[299]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[99],stage1_23[105],stage1_22[140],stage1_21[201]}
   );
   gpc615_5 gpc928 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340]},
      {stage0_22[300]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[100],stage1_23[106],stage1_22[141],stage1_21[202]}
   );
   gpc615_5 gpc929 (
      {stage0_21[341], stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345]},
      {stage0_22[301]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[101],stage1_23[107],stage1_22[142],stage1_21[203]}
   );
   gpc615_5 gpc930 (
      {stage0_21[346], stage0_21[347], stage0_21[348], stage0_21[349], stage0_21[350]},
      {stage0_22[302]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[102],stage1_23[108],stage1_22[143],stage1_21[204]}
   );
   gpc615_5 gpc931 (
      {stage0_21[351], stage0_21[352], stage0_21[353], stage0_21[354], stage0_21[355]},
      {stage0_22[303]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[103],stage1_23[109],stage1_22[144],stage1_21[205]}
   );
   gpc615_5 gpc932 (
      {stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359], stage0_21[360]},
      {stage0_22[304]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[104],stage1_23[110],stage1_22[145],stage1_21[206]}
   );
   gpc615_5 gpc933 (
      {stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_22[305]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[105],stage1_23[111],stage1_22[146],stage1_21[207]}
   );
   gpc615_5 gpc934 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370]},
      {stage0_22[306]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[106],stage1_23[112],stage1_22[147],stage1_21[208]}
   );
   gpc615_5 gpc935 (
      {stage0_21[371], stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375]},
      {stage0_22[307]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[107],stage1_23[113],stage1_22[148],stage1_21[209]}
   );
   gpc615_5 gpc936 (
      {stage0_21[376], stage0_21[377], stage0_21[378], stage0_21[379], stage0_21[380]},
      {stage0_22[308]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[108],stage1_23[114],stage1_22[149],stage1_21[210]}
   );
   gpc615_5 gpc937 (
      {stage0_21[381], stage0_21[382], stage0_21[383], stage0_21[384], stage0_21[385]},
      {stage0_22[309]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[109],stage1_23[115],stage1_22[150],stage1_21[211]}
   );
   gpc615_5 gpc938 (
      {stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389], stage0_21[390]},
      {stage0_22[310]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[110],stage1_23[116],stage1_22[151],stage1_21[212]}
   );
   gpc615_5 gpc939 (
      {stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_22[311]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[111],stage1_23[117],stage1_22[152],stage1_21[213]}
   );
   gpc615_5 gpc940 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400]},
      {stage0_22[312]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[112],stage1_23[118],stage1_22[153],stage1_21[214]}
   );
   gpc615_5 gpc941 (
      {stage0_21[401], stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405]},
      {stage0_22[313]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[113],stage1_23[119],stage1_22[154],stage1_21[215]}
   );
   gpc615_5 gpc942 (
      {stage0_21[406], stage0_21[407], stage0_21[408], stage0_21[409], stage0_21[410]},
      {stage0_22[314]},
      {stage0_23[396], stage0_23[397], stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401]},
      {stage1_25[66],stage1_24[114],stage1_23[120],stage1_22[155],stage1_21[216]}
   );
   gpc615_5 gpc943 (
      {stage0_21[411], stage0_21[412], stage0_21[413], stage0_21[414], stage0_21[415]},
      {stage0_22[315]},
      {stage0_23[402], stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage1_25[67],stage1_24[115],stage1_23[121],stage1_22[156],stage1_21[217]}
   );
   gpc615_5 gpc944 (
      {stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419], stage0_21[420]},
      {stage0_22[316]},
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412], stage0_23[413]},
      {stage1_25[68],stage1_24[116],stage1_23[122],stage1_22[157],stage1_21[218]}
   );
   gpc615_5 gpc945 (
      {stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_22[317]},
      {stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417], stage0_23[418], stage0_23[419]},
      {stage1_25[69],stage1_24[117],stage1_23[123],stage1_22[158],stage1_21[219]}
   );
   gpc615_5 gpc946 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430]},
      {stage0_22[318]},
      {stage0_23[420], stage0_23[421], stage0_23[422], stage0_23[423], stage0_23[424], stage0_23[425]},
      {stage1_25[70],stage1_24[118],stage1_23[124],stage1_22[159],stage1_21[220]}
   );
   gpc615_5 gpc947 (
      {stage0_21[431], stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435]},
      {stage0_22[319]},
      {stage0_23[426], stage0_23[427], stage0_23[428], stage0_23[429], stage0_23[430], stage0_23[431]},
      {stage1_25[71],stage1_24[119],stage1_23[125],stage1_22[160],stage1_21[221]}
   );
   gpc615_5 gpc948 (
      {stage0_21[436], stage0_21[437], stage0_21[438], stage0_21[439], stage0_21[440]},
      {stage0_22[320]},
      {stage0_23[432], stage0_23[433], stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437]},
      {stage1_25[72],stage1_24[120],stage1_23[126],stage1_22[161],stage1_21[222]}
   );
   gpc615_5 gpc949 (
      {stage0_21[441], stage0_21[442], stage0_21[443], stage0_21[444], stage0_21[445]},
      {stage0_22[321]},
      {stage0_23[438], stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage1_25[73],stage1_24[121],stage1_23[127],stage1_22[162],stage1_21[223]}
   );
   gpc615_5 gpc950 (
      {stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449], stage0_21[450]},
      {stage0_22[322]},
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448], stage0_23[449]},
      {stage1_25[74],stage1_24[122],stage1_23[128],stage1_22[163],stage1_21[224]}
   );
   gpc615_5 gpc951 (
      {stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_22[323]},
      {stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453], stage0_23[454], stage0_23[455]},
      {stage1_25[75],stage1_24[123],stage1_23[129],stage1_22[164],stage1_21[225]}
   );
   gpc615_5 gpc952 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460]},
      {stage0_22[324]},
      {stage0_23[456], stage0_23[457], stage0_23[458], stage0_23[459], stage0_23[460], stage0_23[461]},
      {stage1_25[76],stage1_24[124],stage1_23[130],stage1_22[165],stage1_21[226]}
   );
   gpc615_5 gpc953 (
      {stage0_21[461], stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465]},
      {stage0_22[325]},
      {stage0_23[462], stage0_23[463], stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467]},
      {stage1_25[77],stage1_24[125],stage1_23[131],stage1_22[166],stage1_21[227]}
   );
   gpc615_5 gpc954 (
      {stage0_21[466], stage0_21[467], stage0_21[468], stage0_21[469], stage0_21[470]},
      {stage0_22[326]},
      {stage0_23[468], stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage1_25[78],stage1_24[126],stage1_23[132],stage1_22[167],stage1_21[228]}
   );
   gpc606_5 gpc955 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[79],stage1_24[127],stage1_23[133],stage1_22[168]}
   );
   gpc606_5 gpc956 (
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[80],stage1_24[128],stage1_23[134],stage1_22[169]}
   );
   gpc606_5 gpc957 (
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[81],stage1_24[129],stage1_23[135],stage1_22[170]}
   );
   gpc606_5 gpc958 (
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[82],stage1_24[130],stage1_23[136],stage1_22[171]}
   );
   gpc606_5 gpc959 (
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[83],stage1_24[131],stage1_23[137],stage1_22[172]}
   );
   gpc606_5 gpc960 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[84],stage1_24[132],stage1_23[138],stage1_22[173]}
   );
   gpc606_5 gpc961 (
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[85],stage1_24[133],stage1_23[139],stage1_22[174]}
   );
   gpc606_5 gpc962 (
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[86],stage1_24[134],stage1_23[140],stage1_22[175]}
   );
   gpc606_5 gpc963 (
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[87],stage1_24[135],stage1_23[141],stage1_22[176]}
   );
   gpc606_5 gpc964 (
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[88],stage1_24[136],stage1_23[142],stage1_22[177]}
   );
   gpc606_5 gpc965 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391], stage0_22[392]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[89],stage1_24[137],stage1_23[143],stage1_22[178]}
   );
   gpc615_5 gpc966 (
      {stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396], stage0_22[397]},
      {stage0_23[474]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[90],stage1_24[138],stage1_23[144],stage1_22[179]}
   );
   gpc615_5 gpc967 (
      {stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401], stage0_22[402]},
      {stage0_23[475]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[91],stage1_24[139],stage1_23[145],stage1_22[180]}
   );
   gpc615_5 gpc968 (
      {stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage0_23[476]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[92],stage1_24[140],stage1_23[146],stage1_22[181]}
   );
   gpc615_5 gpc969 (
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412]},
      {stage0_23[477]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[93],stage1_24[141],stage1_23[147],stage1_22[182]}
   );
   gpc615_5 gpc970 (
      {stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417]},
      {stage0_23[478]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[94],stage1_24[142],stage1_23[148],stage1_22[183]}
   );
   gpc615_5 gpc971 (
      {stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421], stage0_22[422]},
      {stage0_23[479]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[95],stage1_24[143],stage1_23[149],stage1_22[184]}
   );
   gpc615_5 gpc972 (
      {stage0_23[480], stage0_23[481], stage0_23[482], stage0_23[483], stage0_23[484]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[96],stage1_24[144],stage1_23[150]}
   );
   gpc615_5 gpc973 (
      {stage0_23[485], stage0_23[486], stage0_23[487], stage0_23[488], stage0_23[489]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[97],stage1_24[145],stage1_23[151]}
   );
   gpc615_5 gpc974 (
      {stage0_23[490], stage0_23[491], stage0_23[492], stage0_23[493], stage0_23[494]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[98],stage1_24[146],stage1_23[152]}
   );
   gpc615_5 gpc975 (
      {stage0_23[495], stage0_23[496], stage0_23[497], stage0_23[498], stage0_23[499]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[99],stage1_24[147],stage1_23[153]}
   );
   gpc606_5 gpc976 (
      {stage0_24[106], stage0_24[107], stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[4],stage1_26[21],stage1_25[100],stage1_24[148]}
   );
   gpc606_5 gpc977 (
      {stage0_24[112], stage0_24[113], stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[5],stage1_26[22],stage1_25[101],stage1_24[149]}
   );
   gpc606_5 gpc978 (
      {stage0_24[118], stage0_24[119], stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[6],stage1_26[23],stage1_25[102],stage1_24[150]}
   );
   gpc606_5 gpc979 (
      {stage0_24[124], stage0_24[125], stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[7],stage1_26[24],stage1_25[103],stage1_24[151]}
   );
   gpc606_5 gpc980 (
      {stage0_24[130], stage0_24[131], stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[8],stage1_26[25],stage1_25[104],stage1_24[152]}
   );
   gpc606_5 gpc981 (
      {stage0_24[136], stage0_24[137], stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[9],stage1_26[26],stage1_25[105],stage1_24[153]}
   );
   gpc606_5 gpc982 (
      {stage0_24[142], stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[10],stage1_26[27],stage1_25[106],stage1_24[154]}
   );
   gpc606_5 gpc983 (
      {stage0_24[148], stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[11],stage1_26[28],stage1_25[107],stage1_24[155]}
   );
   gpc606_5 gpc984 (
      {stage0_24[154], stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[12],stage1_26[29],stage1_25[108],stage1_24[156]}
   );
   gpc606_5 gpc985 (
      {stage0_24[160], stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[13],stage1_26[30],stage1_25[109],stage1_24[157]}
   );
   gpc606_5 gpc986 (
      {stage0_24[166], stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[14],stage1_26[31],stage1_25[110],stage1_24[158]}
   );
   gpc606_5 gpc987 (
      {stage0_24[172], stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[15],stage1_26[32],stage1_25[111],stage1_24[159]}
   );
   gpc606_5 gpc988 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[16],stage1_26[33],stage1_25[112],stage1_24[160]}
   );
   gpc606_5 gpc989 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[17],stage1_26[34],stage1_25[113],stage1_24[161]}
   );
   gpc606_5 gpc990 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[18],stage1_26[35],stage1_25[114],stage1_24[162]}
   );
   gpc606_5 gpc991 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[19],stage1_26[36],stage1_25[115],stage1_24[163]}
   );
   gpc606_5 gpc992 (
      {stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[20],stage1_26[37],stage1_25[116],stage1_24[164]}
   );
   gpc606_5 gpc993 (
      {stage0_24[208], stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[21],stage1_26[38],stage1_25[117],stage1_24[165]}
   );
   gpc606_5 gpc994 (
      {stage0_24[214], stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[22],stage1_26[39],stage1_25[118],stage1_24[166]}
   );
   gpc606_5 gpc995 (
      {stage0_24[220], stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[23],stage1_26[40],stage1_25[119],stage1_24[167]}
   );
   gpc606_5 gpc996 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[24],stage1_26[41],stage1_25[120],stage1_24[168]}
   );
   gpc606_5 gpc997 (
      {stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[25],stage1_26[42],stage1_25[121],stage1_24[169]}
   );
   gpc606_5 gpc998 (
      {stage0_24[238], stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[26],stage1_26[43],stage1_25[122],stage1_24[170]}
   );
   gpc606_5 gpc999 (
      {stage0_24[244], stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[27],stage1_26[44],stage1_25[123],stage1_24[171]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[250], stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[28],stage1_26[45],stage1_25[124],stage1_24[172]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[29],stage1_26[46],stage1_25[125],stage1_24[173]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[30],stage1_26[47],stage1_25[126],stage1_24[174]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[268], stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[31],stage1_26[48],stage1_25[127],stage1_24[175]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[274], stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[32],stage1_26[49],stage1_25[128],stage1_24[176]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[280], stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[33],stage1_26[50],stage1_25[129],stage1_24[177]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[34],stage1_26[51],stage1_25[130],stage1_24[178]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[35],stage1_26[52],stage1_25[131],stage1_24[179]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[298], stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[36],stage1_26[53],stage1_25[132],stage1_24[180]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[304], stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[37],stage1_26[54],stage1_25[133],stage1_24[181]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[310], stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[38],stage1_26[55],stage1_25[134],stage1_24[182]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[39],stage1_26[56],stage1_25[135],stage1_24[183]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[40],stage1_26[57],stage1_25[136],stage1_24[184]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[328], stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[41],stage1_26[58],stage1_25[137],stage1_24[185]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[334], stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[42],stage1_26[59],stage1_25[138],stage1_24[186]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[340], stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[43],stage1_26[60],stage1_25[139],stage1_24[187]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[44],stage1_26[61],stage1_25[140],stage1_24[188]}
   );
   gpc615_5 gpc1017 (
      {stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356]},
      {stage0_25[24]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[45],stage1_26[62],stage1_25[141],stage1_24[189]}
   );
   gpc615_5 gpc1018 (
      {stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360], stage0_24[361]},
      {stage0_25[25]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[46],stage1_26[63],stage1_25[142],stage1_24[190]}
   );
   gpc615_5 gpc1019 (
      {stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_25[26]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[47],stage1_26[64],stage1_25[143],stage1_24[191]}
   );
   gpc615_5 gpc1020 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371]},
      {stage0_25[27]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[48],stage1_26[65],stage1_25[144],stage1_24[192]}
   );
   gpc615_5 gpc1021 (
      {stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_25[28]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[49],stage1_26[66],stage1_25[145],stage1_24[193]}
   );
   gpc615_5 gpc1022 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381]},
      {stage0_25[29]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[50],stage1_26[67],stage1_25[146],stage1_24[194]}
   );
   gpc615_5 gpc1023 (
      {stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386]},
      {stage0_25[30]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[51],stage1_26[68],stage1_25[147],stage1_24[195]}
   );
   gpc615_5 gpc1024 (
      {stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390], stage0_24[391]},
      {stage0_25[31]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[52],stage1_26[69],stage1_25[148],stage1_24[196]}
   );
   gpc615_5 gpc1025 (
      {stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_25[32]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[53],stage1_26[70],stage1_25[149],stage1_24[197]}
   );
   gpc615_5 gpc1026 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401]},
      {stage0_25[33]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[54],stage1_26[71],stage1_25[150],stage1_24[198]}
   );
   gpc615_5 gpc1027 (
      {stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_25[34]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[55],stage1_26[72],stage1_25[151],stage1_24[199]}
   );
   gpc615_5 gpc1028 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411]},
      {stage0_25[35]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[56],stage1_26[73],stage1_25[152],stage1_24[200]}
   );
   gpc615_5 gpc1029 (
      {stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416]},
      {stage0_25[36]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[57],stage1_26[74],stage1_25[153],stage1_24[201]}
   );
   gpc615_5 gpc1030 (
      {stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420], stage0_24[421]},
      {stage0_25[37]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[58],stage1_26[75],stage1_25[154],stage1_24[202]}
   );
   gpc615_5 gpc1031 (
      {stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_25[38]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[59],stage1_26[76],stage1_25[155],stage1_24[203]}
   );
   gpc615_5 gpc1032 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431]},
      {stage0_25[39]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[60],stage1_26[77],stage1_25[156],stage1_24[204]}
   );
   gpc615_5 gpc1033 (
      {stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_25[40]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[61],stage1_26[78],stage1_25[157],stage1_24[205]}
   );
   gpc615_5 gpc1034 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441]},
      {stage0_25[41]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[62],stage1_26[79],stage1_25[158],stage1_24[206]}
   );
   gpc615_5 gpc1035 (
      {stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446]},
      {stage0_25[42]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[63],stage1_26[80],stage1_25[159],stage1_24[207]}
   );
   gpc615_5 gpc1036 (
      {stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450], stage0_24[451]},
      {stage0_25[43]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[64],stage1_26[81],stage1_25[160],stage1_24[208]}
   );
   gpc615_5 gpc1037 (
      {stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_25[44]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[65],stage1_26[82],stage1_25[161],stage1_24[209]}
   );
   gpc615_5 gpc1038 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461]},
      {stage0_25[45]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[66],stage1_26[83],stage1_25[162],stage1_24[210]}
   );
   gpc615_5 gpc1039 (
      {stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_25[46]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[67],stage1_26[84],stage1_25[163],stage1_24[211]}
   );
   gpc615_5 gpc1040 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471]},
      {stage0_25[47]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[68],stage1_26[85],stage1_25[164],stage1_24[212]}
   );
   gpc615_5 gpc1041 (
      {stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476]},
      {stage0_25[48]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[69],stage1_26[86],stage1_25[165],stage1_24[213]}
   );
   gpc615_5 gpc1042 (
      {stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480], stage0_24[481]},
      {stage0_25[49]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[70],stage1_26[87],stage1_25[166],stage1_24[214]}
   );
   gpc615_5 gpc1043 (
      {stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_25[50]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[71],stage1_26[88],stage1_25[167],stage1_24[215]}
   );
   gpc615_5 gpc1044 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491]},
      {stage0_25[51]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[72],stage1_26[89],stage1_25[168],stage1_24[216]}
   );
   gpc615_5 gpc1045 (
      {stage0_24[492], stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496]},
      {stage0_25[52]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[73],stage1_26[90],stage1_25[169],stage1_24[217]}
   );
   gpc615_5 gpc1046 (
      {stage0_24[497], stage0_24[498], stage0_24[499], stage0_24[500], stage0_24[501]},
      {stage0_25[53]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[74],stage1_26[91],stage1_25[170],stage1_24[218]}
   );
   gpc615_5 gpc1047 (
      {stage0_24[502], stage0_24[503], stage0_24[504], stage0_24[505], stage0_24[506]},
      {stage0_25[54]},
      {stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429], stage0_26[430], stage0_26[431]},
      {stage1_28[71],stage1_27[75],stage1_26[92],stage1_25[171],stage1_24[219]}
   );
   gpc615_5 gpc1048 (
      {stage0_24[507], stage0_24[508], stage0_24[509], stage0_24[510], stage0_24[511]},
      {stage0_25[55]},
      {stage0_26[432], stage0_26[433], stage0_26[434], stage0_26[435], stage0_26[436], stage0_26[437]},
      {stage1_28[72],stage1_27[76],stage1_26[93],stage1_25[172],stage1_24[220]}
   );
   gpc606_5 gpc1049 (
      {stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[73],stage1_27[77],stage1_26[94],stage1_25[173]}
   );
   gpc606_5 gpc1050 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66], stage0_25[67]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[74],stage1_27[78],stage1_26[95],stage1_25[174]}
   );
   gpc606_5 gpc1051 (
      {stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71], stage0_25[72], stage0_25[73]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[75],stage1_27[79],stage1_26[96],stage1_25[175]}
   );
   gpc606_5 gpc1052 (
      {stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77], stage0_25[78], stage0_25[79]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[76],stage1_27[80],stage1_26[97],stage1_25[176]}
   );
   gpc606_5 gpc1053 (
      {stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[77],stage1_27[81],stage1_26[98],stage1_25[177]}
   );
   gpc606_5 gpc1054 (
      {stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[78],stage1_27[82],stage1_26[99],stage1_25[178]}
   );
   gpc606_5 gpc1055 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96], stage0_25[97]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[79],stage1_27[83],stage1_26[100],stage1_25[179]}
   );
   gpc606_5 gpc1056 (
      {stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101], stage0_25[102], stage0_25[103]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[80],stage1_27[84],stage1_26[101],stage1_25[180]}
   );
   gpc606_5 gpc1057 (
      {stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107], stage0_25[108], stage0_25[109]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[81],stage1_27[85],stage1_26[102],stage1_25[181]}
   );
   gpc606_5 gpc1058 (
      {stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[82],stage1_27[86],stage1_26[103],stage1_25[182]}
   );
   gpc606_5 gpc1059 (
      {stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[83],stage1_27[87],stage1_26[104],stage1_25[183]}
   );
   gpc606_5 gpc1060 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[84],stage1_27[88],stage1_26[105],stage1_25[184]}
   );
   gpc606_5 gpc1061 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[85],stage1_27[89],stage1_26[106],stage1_25[185]}
   );
   gpc606_5 gpc1062 (
      {stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[86],stage1_27[90],stage1_26[107],stage1_25[186]}
   );
   gpc606_5 gpc1063 (
      {stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[87],stage1_27[91],stage1_26[108],stage1_25[187]}
   );
   gpc606_5 gpc1064 (
      {stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[88],stage1_27[92],stage1_26[109],stage1_25[188]}
   );
   gpc606_5 gpc1065 (
      {stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[89],stage1_27[93],stage1_26[110],stage1_25[189]}
   );
   gpc606_5 gpc1066 (
      {stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[90],stage1_27[94],stage1_26[111],stage1_25[190]}
   );
   gpc606_5 gpc1067 (
      {stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[91],stage1_27[95],stage1_26[112],stage1_25[191]}
   );
   gpc606_5 gpc1068 (
      {stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[92],stage1_27[96],stage1_26[113],stage1_25[192]}
   );
   gpc606_5 gpc1069 (
      {stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[93],stage1_27[97],stage1_26[114],stage1_25[193]}
   );
   gpc606_5 gpc1070 (
      {stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[94],stage1_27[98],stage1_26[115],stage1_25[194]}
   );
   gpc606_5 gpc1071 (
      {stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[95],stage1_27[99],stage1_26[116],stage1_25[195]}
   );
   gpc606_5 gpc1072 (
      {stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[96],stage1_27[100],stage1_26[117],stage1_25[196]}
   );
   gpc606_5 gpc1073 (
      {stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[97],stage1_27[101],stage1_26[118],stage1_25[197]}
   );
   gpc606_5 gpc1074 (
      {stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[98],stage1_27[102],stage1_26[119],stage1_25[198]}
   );
   gpc606_5 gpc1075 (
      {stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[99],stage1_27[103],stage1_26[120],stage1_25[199]}
   );
   gpc606_5 gpc1076 (
      {stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[100],stage1_27[104],stage1_26[121],stage1_25[200]}
   );
   gpc606_5 gpc1077 (
      {stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[101],stage1_27[105],stage1_26[122],stage1_25[201]}
   );
   gpc606_5 gpc1078 (
      {stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[102],stage1_27[106],stage1_26[123],stage1_25[202]}
   );
   gpc606_5 gpc1079 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240], stage0_25[241]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[103],stage1_27[107],stage1_26[124],stage1_25[203]}
   );
   gpc606_5 gpc1080 (
      {stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245], stage0_25[246], stage0_25[247]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[104],stage1_27[108],stage1_26[125],stage1_25[204]}
   );
   gpc606_5 gpc1081 (
      {stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251], stage0_25[252], stage0_25[253]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[105],stage1_27[109],stage1_26[126],stage1_25[205]}
   );
   gpc606_5 gpc1082 (
      {stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[106],stage1_27[110],stage1_26[127],stage1_25[206]}
   );
   gpc606_5 gpc1083 (
      {stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[107],stage1_27[111],stage1_26[128],stage1_25[207]}
   );
   gpc606_5 gpc1084 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270], stage0_25[271]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[108],stage1_27[112],stage1_26[129],stage1_25[208]}
   );
   gpc606_5 gpc1085 (
      {stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275], stage0_25[276], stage0_25[277]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[109],stage1_27[113],stage1_26[130],stage1_25[209]}
   );
   gpc606_5 gpc1086 (
      {stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281], stage0_25[282], stage0_25[283]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[110],stage1_27[114],stage1_26[131],stage1_25[210]}
   );
   gpc606_5 gpc1087 (
      {stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[111],stage1_27[115],stage1_26[132],stage1_25[211]}
   );
   gpc606_5 gpc1088 (
      {stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[112],stage1_27[116],stage1_26[133],stage1_25[212]}
   );
   gpc606_5 gpc1089 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300], stage0_25[301]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[113],stage1_27[117],stage1_26[134],stage1_25[213]}
   );
   gpc606_5 gpc1090 (
      {stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305], stage0_25[306], stage0_25[307]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[114],stage1_27[118],stage1_26[135],stage1_25[214]}
   );
   gpc606_5 gpc1091 (
      {stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311], stage0_25[312], stage0_25[313]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[115],stage1_27[119],stage1_26[136],stage1_25[215]}
   );
   gpc606_5 gpc1092 (
      {stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[116],stage1_27[120],stage1_26[137],stage1_25[216]}
   );
   gpc606_5 gpc1093 (
      {stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[117],stage1_27[121],stage1_26[138],stage1_25[217]}
   );
   gpc606_5 gpc1094 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330], stage0_25[331]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[118],stage1_27[122],stage1_26[139],stage1_25[218]}
   );
   gpc606_5 gpc1095 (
      {stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335], stage0_25[336], stage0_25[337]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[119],stage1_27[123],stage1_26[140],stage1_25[219]}
   );
   gpc606_5 gpc1096 (
      {stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341], stage0_25[342], stage0_25[343]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[120],stage1_27[124],stage1_26[141],stage1_25[220]}
   );
   gpc606_5 gpc1097 (
      {stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[121],stage1_27[125],stage1_26[142],stage1_25[221]}
   );
   gpc606_5 gpc1098 (
      {stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[122],stage1_27[126],stage1_26[143],stage1_25[222]}
   );
   gpc606_5 gpc1099 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360], stage0_25[361]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[123],stage1_27[127],stage1_26[144],stage1_25[223]}
   );
   gpc606_5 gpc1100 (
      {stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365], stage0_25[366], stage0_25[367]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[124],stage1_27[128],stage1_26[145],stage1_25[224]}
   );
   gpc606_5 gpc1101 (
      {stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371], stage0_25[372], stage0_25[373]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[125],stage1_27[129],stage1_26[146],stage1_25[225]}
   );
   gpc606_5 gpc1102 (
      {stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[126],stage1_27[130],stage1_26[147],stage1_25[226]}
   );
   gpc606_5 gpc1103 (
      {stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[127],stage1_27[131],stage1_26[148],stage1_25[227]}
   );
   gpc606_5 gpc1104 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390], stage0_25[391]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[128],stage1_27[132],stage1_26[149],stage1_25[228]}
   );
   gpc606_5 gpc1105 (
      {stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395], stage0_25[396], stage0_25[397]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[129],stage1_27[133],stage1_26[150],stage1_25[229]}
   );
   gpc606_5 gpc1106 (
      {stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401], stage0_25[402], stage0_25[403]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[130],stage1_27[134],stage1_26[151],stage1_25[230]}
   );
   gpc606_5 gpc1107 (
      {stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[131],stage1_27[135],stage1_26[152],stage1_25[231]}
   );
   gpc606_5 gpc1108 (
      {stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[132],stage1_27[136],stage1_26[153],stage1_25[232]}
   );
   gpc606_5 gpc1109 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420], stage0_25[421]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[133],stage1_27[137],stage1_26[154],stage1_25[233]}
   );
   gpc606_5 gpc1110 (
      {stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425], stage0_25[426], stage0_25[427]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[134],stage1_27[138],stage1_26[155],stage1_25[234]}
   );
   gpc606_5 gpc1111 (
      {stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431], stage0_25[432], stage0_25[433]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[135],stage1_27[139],stage1_26[156],stage1_25[235]}
   );
   gpc606_5 gpc1112 (
      {stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[136],stage1_27[140],stage1_26[157],stage1_25[236]}
   );
   gpc606_5 gpc1113 (
      {stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[137],stage1_27[141],stage1_26[158],stage1_25[237]}
   );
   gpc606_5 gpc1114 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450], stage0_25[451]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[138],stage1_27[142],stage1_26[159],stage1_25[238]}
   );
   gpc606_5 gpc1115 (
      {stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455], stage0_25[456], stage0_25[457]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[139],stage1_27[143],stage1_26[160],stage1_25[239]}
   );
   gpc606_5 gpc1116 (
      {stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461], stage0_25[462], stage0_25[463]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[140],stage1_27[144],stage1_26[161],stage1_25[240]}
   );
   gpc606_5 gpc1117 (
      {stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[141],stage1_27[145],stage1_26[162],stage1_25[241]}
   );
   gpc606_5 gpc1118 (
      {stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[142],stage1_27[146],stage1_26[163],stage1_25[242]}
   );
   gpc606_5 gpc1119 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480], stage0_25[481]},
      {stage0_27[420], stage0_27[421], stage0_27[422], stage0_27[423], stage0_27[424], stage0_27[425]},
      {stage1_29[70],stage1_28[143],stage1_27[147],stage1_26[164],stage1_25[243]}
   );
   gpc615_5 gpc1120 (
      {stage0_26[438], stage0_26[439], stage0_26[440], stage0_26[441], stage0_26[442]},
      {stage0_27[426]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[71],stage1_28[144],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1121 (
      {stage0_26[443], stage0_26[444], stage0_26[445], stage0_26[446], stage0_26[447]},
      {stage0_27[427]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[72],stage1_28[145],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1122 (
      {stage0_26[448], stage0_26[449], stage0_26[450], stage0_26[451], stage0_26[452]},
      {stage0_27[428]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[73],stage1_28[146],stage1_27[150],stage1_26[167]}
   );
   gpc615_5 gpc1123 (
      {stage0_26[453], stage0_26[454], stage0_26[455], stage0_26[456], stage0_26[457]},
      {stage0_27[429]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[74],stage1_28[147],stage1_27[151],stage1_26[168]}
   );
   gpc615_5 gpc1124 (
      {stage0_26[458], stage0_26[459], stage0_26[460], stage0_26[461], stage0_26[462]},
      {stage0_27[430]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[75],stage1_28[148],stage1_27[152],stage1_26[169]}
   );
   gpc615_5 gpc1125 (
      {stage0_26[463], stage0_26[464], stage0_26[465], stage0_26[466], stage0_26[467]},
      {stage0_27[431]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[76],stage1_28[149],stage1_27[153],stage1_26[170]}
   );
   gpc615_5 gpc1126 (
      {stage0_26[468], stage0_26[469], stage0_26[470], stage0_26[471], stage0_26[472]},
      {stage0_27[432]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[77],stage1_28[150],stage1_27[154],stage1_26[171]}
   );
   gpc615_5 gpc1127 (
      {stage0_26[473], stage0_26[474], stage0_26[475], stage0_26[476], stage0_26[477]},
      {stage0_27[433]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[78],stage1_28[151],stage1_27[155],stage1_26[172]}
   );
   gpc615_5 gpc1128 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[434]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[79],stage1_28[152],stage1_27[156],stage1_26[173]}
   );
   gpc615_5 gpc1129 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[435]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[80],stage1_28[153],stage1_27[157],stage1_26[174]}
   );
   gpc615_5 gpc1130 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[436]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[81],stage1_28[154],stage1_27[158],stage1_26[175]}
   );
   gpc615_5 gpc1131 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[437]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[82],stage1_28[155],stage1_27[159],stage1_26[176]}
   );
   gpc606_5 gpc1132 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442], stage0_27[443]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[83],stage1_28[156],stage1_27[160]}
   );
   gpc606_5 gpc1133 (
      {stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447], stage0_27[448], stage0_27[449]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[84],stage1_28[157],stage1_27[161]}
   );
   gpc606_5 gpc1134 (
      {stage0_27[450], stage0_27[451], stage0_27[452], stage0_27[453], stage0_27[454], stage0_27[455]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[85],stage1_28[158],stage1_27[162]}
   );
   gpc606_5 gpc1135 (
      {stage0_27[456], stage0_27[457], stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[86],stage1_28[159],stage1_27[163]}
   );
   gpc606_5 gpc1136 (
      {stage0_27[462], stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[87],stage1_28[160],stage1_27[164]}
   );
   gpc606_5 gpc1137 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472], stage0_27[473]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[88],stage1_28[161],stage1_27[165]}
   );
   gpc615_5 gpc1138 (
      {stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477], stage0_27[478]},
      {stage0_28[72]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[89],stage1_28[162],stage1_27[166]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[19],stage1_29[90],stage1_28[163]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[20],stage1_29[91],stage1_28[164]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[21],stage1_29[92],stage1_28[165]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[22],stage1_29[93],stage1_28[166]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[23],stage1_29[94],stage1_28[167]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[24],stage1_29[95],stage1_28[168]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[25],stage1_29[96],stage1_28[169]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[26],stage1_29[97],stage1_28[170]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[27],stage1_29[98],stage1_28[171]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[28],stage1_29[99],stage1_28[172]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[29],stage1_29[100],stage1_28[173]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[30],stage1_29[101],stage1_28[174]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[31],stage1_29[102],stage1_28[175]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[32],stage1_29[103],stage1_28[176]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[33],stage1_29[104],stage1_28[177]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[34],stage1_29[105],stage1_28[178]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[35],stage1_29[106],stage1_28[179]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[36],stage1_29[107],stage1_28[180]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[37],stage1_29[108],stage1_28[181]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[38],stage1_29[109],stage1_28[182]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[39],stage1_29[110],stage1_28[183]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[40],stage1_29[111],stage1_28[184]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[41],stage1_29[112],stage1_28[185]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[42],stage1_29[113],stage1_28[186]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[43],stage1_29[114],stage1_28[187]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[44],stage1_29[115],stage1_28[188]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[45],stage1_29[116],stage1_28[189]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[46],stage1_29[117],stage1_28[190]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[47],stage1_29[118],stage1_28[191]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[48],stage1_29[119],stage1_28[192]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[49],stage1_29[120],stage1_28[193]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[50],stage1_29[121],stage1_28[194]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[51],stage1_29[122],stage1_28[195]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[52],stage1_29[123],stage1_28[196]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[53],stage1_29[124],stage1_28[197]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[54],stage1_29[125],stage1_28[198]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[55],stage1_29[126],stage1_28[199]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[56],stage1_29[127],stage1_28[200]}
   );
   gpc615_5 gpc1177 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_29[42]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[57],stage1_29[128],stage1_28[201]}
   );
   gpc615_5 gpc1178 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310]},
      {stage0_29[43]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[58],stage1_29[129],stage1_28[202]}
   );
   gpc615_5 gpc1179 (
      {stage0_28[311], stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315]},
      {stage0_29[44]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[47],stage1_30[59],stage1_29[130],stage1_28[203]}
   );
   gpc615_5 gpc1180 (
      {stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319], stage0_28[320]},
      {stage0_29[45]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[48],stage1_30[60],stage1_29[131],stage1_28[204]}
   );
   gpc615_5 gpc1181 (
      {stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_29[46]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[49],stage1_30[61],stage1_29[132],stage1_28[205]}
   );
   gpc615_5 gpc1182 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_29[47]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[50],stage1_30[62],stage1_29[133],stage1_28[206]}
   );
   gpc615_5 gpc1183 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_29[48]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[51],stage1_30[63],stage1_29[134],stage1_28[207]}
   );
   gpc615_5 gpc1184 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340]},
      {stage0_29[49]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[52],stage1_30[64],stage1_29[135],stage1_28[208]}
   );
   gpc615_5 gpc1185 (
      {stage0_28[341], stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345]},
      {stage0_29[50]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[53],stage1_30[65],stage1_29[136],stage1_28[209]}
   );
   gpc615_5 gpc1186 (
      {stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349], stage0_28[350]},
      {stage0_29[51]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[54],stage1_30[66],stage1_29[137],stage1_28[210]}
   );
   gpc615_5 gpc1187 (
      {stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_29[52]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[55],stage1_30[67],stage1_29[138],stage1_28[211]}
   );
   gpc615_5 gpc1188 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_29[53]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[56],stage1_30[68],stage1_29[139],stage1_28[212]}
   );
   gpc615_5 gpc1189 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_29[54]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[57],stage1_30[69],stage1_29[140],stage1_28[213]}
   );
   gpc615_5 gpc1190 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370]},
      {stage0_29[55]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[58],stage1_30[70],stage1_29[141],stage1_28[214]}
   );
   gpc615_5 gpc1191 (
      {stage0_28[371], stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375]},
      {stage0_29[56]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[59],stage1_30[71],stage1_29[142],stage1_28[215]}
   );
   gpc615_5 gpc1192 (
      {stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379], stage0_28[380]},
      {stage0_29[57]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[60],stage1_30[72],stage1_29[143],stage1_28[216]}
   );
   gpc615_5 gpc1193 (
      {stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_29[58]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[61],stage1_30[73],stage1_29[144],stage1_28[217]}
   );
   gpc615_5 gpc1194 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_29[59]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[62],stage1_30[74],stage1_29[145],stage1_28[218]}
   );
   gpc615_5 gpc1195 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_29[60]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[63],stage1_30[75],stage1_29[146],stage1_28[219]}
   );
   gpc615_5 gpc1196 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400]},
      {stage0_29[61]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[64],stage1_30[76],stage1_29[147],stage1_28[220]}
   );
   gpc615_5 gpc1197 (
      {stage0_28[401], stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405]},
      {stage0_29[62]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[65],stage1_30[77],stage1_29[148],stage1_28[221]}
   );
   gpc615_5 gpc1198 (
      {stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409], stage0_28[410]},
      {stage0_29[63]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[66],stage1_30[78],stage1_29[149],stage1_28[222]}
   );
   gpc615_5 gpc1199 (
      {stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_29[64]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[67],stage1_30[79],stage1_29[150],stage1_28[223]}
   );
   gpc615_5 gpc1200 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_29[65]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[68],stage1_30[80],stage1_29[151],stage1_28[224]}
   );
   gpc615_5 gpc1201 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_29[66]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[69],stage1_30[81],stage1_29[152],stage1_28[225]}
   );
   gpc615_5 gpc1202 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430]},
      {stage0_29[67]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[70],stage1_30[82],stage1_29[153],stage1_28[226]}
   );
   gpc615_5 gpc1203 (
      {stage0_28[431], stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435]},
      {stage0_29[68]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[71],stage1_30[83],stage1_29[154],stage1_28[227]}
   );
   gpc615_5 gpc1204 (
      {stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439], stage0_28[440]},
      {stage0_29[69]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[72],stage1_30[84],stage1_29[155],stage1_28[228]}
   );
   gpc615_5 gpc1205 (
      {stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_29[70]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[73],stage1_30[85],stage1_29[156],stage1_28[229]}
   );
   gpc615_5 gpc1206 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_29[71]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[74],stage1_30[86],stage1_29[157],stage1_28[230]}
   );
   gpc615_5 gpc1207 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455]},
      {stage0_29[72]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[75],stage1_30[87],stage1_29[158],stage1_28[231]}
   );
   gpc615_5 gpc1208 (
      {stage0_28[456], stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460]},
      {stage0_29[73]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[76],stage1_30[88],stage1_29[159],stage1_28[232]}
   );
   gpc615_5 gpc1209 (
      {stage0_28[461], stage0_28[462], stage0_28[463], stage0_28[464], stage0_28[465]},
      {stage0_29[74]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[77],stage1_30[89],stage1_29[160],stage1_28[233]}
   );
   gpc615_5 gpc1210 (
      {stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469], stage0_28[470]},
      {stage0_29[75]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[78],stage1_30[90],stage1_29[161],stage1_28[234]}
   );
   gpc615_5 gpc1211 (
      {stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_29[76]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[79],stage1_30[91],stage1_29[162],stage1_28[235]}
   );
   gpc615_5 gpc1212 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480]},
      {stage0_29[77]},
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443]},
      {stage1_32[73],stage1_31[80],stage1_30[92],stage1_29[163],stage1_28[236]}
   );
   gpc615_5 gpc1213 (
      {stage0_28[481], stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485]},
      {stage0_29[78]},
      {stage0_30[444], stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage1_32[74],stage1_31[81],stage1_30[93],stage1_29[164],stage1_28[237]}
   );
   gpc615_5 gpc1214 (
      {stage0_28[486], stage0_28[487], stage0_28[488], stage0_28[489], stage0_28[490]},
      {stage0_29[79]},
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454], stage0_30[455]},
      {stage1_32[75],stage1_31[82],stage1_30[94],stage1_29[165],stage1_28[238]}
   );
   gpc615_5 gpc1215 (
      {stage0_28[491], stage0_28[492], stage0_28[493], stage0_28[494], stage0_28[495]},
      {stage0_29[80]},
      {stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459], stage0_30[460], stage0_30[461]},
      {stage1_32[76],stage1_31[83],stage1_30[95],stage1_29[166],stage1_28[239]}
   );
   gpc615_5 gpc1216 (
      {stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499], stage0_28[500]},
      {stage0_29[81]},
      {stage0_30[462], stage0_30[463], stage0_30[464], stage0_30[465], stage0_30[466], stage0_30[467]},
      {stage1_32[77],stage1_31[84],stage1_30[96],stage1_29[167],stage1_28[240]}
   );
   gpc615_5 gpc1217 (
      {stage0_28[501], stage0_28[502], stage0_28[503], stage0_28[504], stage0_28[505]},
      {stage0_29[82]},
      {stage0_30[468], stage0_30[469], stage0_30[470], stage0_30[471], stage0_30[472], stage0_30[473]},
      {stage1_32[78],stage1_31[85],stage1_30[97],stage1_29[168],stage1_28[241]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[79],stage1_31[86],stage1_30[98],stage1_29[169]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[80],stage1_31[87],stage1_30[99],stage1_29[170]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[81],stage1_31[88],stage1_30[100],stage1_29[171]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[82],stage1_31[89],stage1_30[101],stage1_29[172]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[83],stage1_31[90],stage1_30[102],stage1_29[173]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[84],stage1_31[91],stage1_30[103],stage1_29[174]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[85],stage1_31[92],stage1_30[104],stage1_29[175]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[86],stage1_31[93],stage1_30[105],stage1_29[176]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[87],stage1_31[94],stage1_30[106],stage1_29[177]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[88],stage1_31[95],stage1_30[107],stage1_29[178]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[89],stage1_31[96],stage1_30[108],stage1_29[179]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[90],stage1_31[97],stage1_30[109],stage1_29[180]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[91],stage1_31[98],stage1_30[110],stage1_29[181]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[161], stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[92],stage1_31[99],stage1_30[111],stage1_29[182]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[167], stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[93],stage1_31[100],stage1_30[112],stage1_29[183]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[173], stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[94],stage1_31[101],stage1_30[113],stage1_29[184]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[179], stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[95],stage1_31[102],stage1_30[114],stage1_29[185]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[185], stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[96],stage1_31[103],stage1_30[115],stage1_29[186]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[97],stage1_31[104],stage1_30[116],stage1_29[187]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[98],stage1_31[105],stage1_30[117],stage1_29[188]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[203], stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[99],stage1_31[106],stage1_30[118],stage1_29[189]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[209], stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[100],stage1_31[107],stage1_30[119],stage1_29[190]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[215], stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[101],stage1_31[108],stage1_30[120],stage1_29[191]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[102],stage1_31[109],stage1_30[121],stage1_29[192]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[103],stage1_31[110],stage1_30[122],stage1_29[193]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[233], stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[104],stage1_31[111],stage1_30[123],stage1_29[194]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[239], stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[105],stage1_31[112],stage1_30[124],stage1_29[195]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[245], stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[106],stage1_31[113],stage1_30[125],stage1_29[196]}
   );
   gpc606_5 gpc1246 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[107],stage1_31[114],stage1_30[126],stage1_29[197]}
   );
   gpc606_5 gpc1247 (
      {stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[108],stage1_31[115],stage1_30[127],stage1_29[198]}
   );
   gpc606_5 gpc1248 (
      {stage0_29[263], stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[109],stage1_31[116],stage1_30[128],stage1_29[199]}
   );
   gpc606_5 gpc1249 (
      {stage0_29[269], stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[110],stage1_31[117],stage1_30[129],stage1_29[200]}
   );
   gpc606_5 gpc1250 (
      {stage0_29[275], stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[111],stage1_31[118],stage1_30[130],stage1_29[201]}
   );
   gpc606_5 gpc1251 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[112],stage1_31[119],stage1_30[131],stage1_29[202]}
   );
   gpc606_5 gpc1252 (
      {stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[113],stage1_31[120],stage1_30[132],stage1_29[203]}
   );
   gpc606_5 gpc1253 (
      {stage0_29[293], stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[114],stage1_31[121],stage1_30[133],stage1_29[204]}
   );
   gpc606_5 gpc1254 (
      {stage0_29[299], stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[115],stage1_31[122],stage1_30[134],stage1_29[205]}
   );
   gpc606_5 gpc1255 (
      {stage0_29[305], stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[116],stage1_31[123],stage1_30[135],stage1_29[206]}
   );
   gpc606_5 gpc1256 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[117],stage1_31[124],stage1_30[136],stage1_29[207]}
   );
   gpc606_5 gpc1257 (
      {stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[118],stage1_31[125],stage1_30[137],stage1_29[208]}
   );
   gpc606_5 gpc1258 (
      {stage0_29[323], stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[119],stage1_31[126],stage1_30[138],stage1_29[209]}
   );
   gpc606_5 gpc1259 (
      {stage0_29[329], stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[120],stage1_31[127],stage1_30[139],stage1_29[210]}
   );
   gpc606_5 gpc1260 (
      {stage0_29[335], stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[121],stage1_31[128],stage1_30[140],stage1_29[211]}
   );
   gpc606_5 gpc1261 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[122],stage1_31[129],stage1_30[141],stage1_29[212]}
   );
   gpc606_5 gpc1262 (
      {stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[123],stage1_31[130],stage1_30[142],stage1_29[213]}
   );
   gpc606_5 gpc1263 (
      {stage0_29[353], stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[124],stage1_31[131],stage1_30[143],stage1_29[214]}
   );
   gpc606_5 gpc1264 (
      {stage0_29[359], stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[125],stage1_31[132],stage1_30[144],stage1_29[215]}
   );
   gpc606_5 gpc1265 (
      {stage0_29[365], stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[126],stage1_31[133],stage1_30[145],stage1_29[216]}
   );
   gpc606_5 gpc1266 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[127],stage1_31[134],stage1_30[146],stage1_29[217]}
   );
   gpc606_5 gpc1267 (
      {stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[128],stage1_31[135],stage1_30[147],stage1_29[218]}
   );
   gpc606_5 gpc1268 (
      {stage0_29[383], stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[129],stage1_31[136],stage1_30[148],stage1_29[219]}
   );
   gpc606_5 gpc1269 (
      {stage0_29[389], stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[130],stage1_31[137],stage1_30[149],stage1_29[220]}
   );
   gpc606_5 gpc1270 (
      {stage0_29[395], stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[131],stage1_31[138],stage1_30[150],stage1_29[221]}
   );
   gpc606_5 gpc1271 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[132],stage1_31[139],stage1_30[151],stage1_29[222]}
   );
   gpc606_5 gpc1272 (
      {stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[133],stage1_31[140],stage1_30[152],stage1_29[223]}
   );
   gpc606_5 gpc1273 (
      {stage0_29[413], stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[134],stage1_31[141],stage1_30[153],stage1_29[224]}
   );
   gpc606_5 gpc1274 (
      {stage0_29[419], stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[135],stage1_31[142],stage1_30[154],stage1_29[225]}
   );
   gpc606_5 gpc1275 (
      {stage0_29[425], stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[136],stage1_31[143],stage1_30[155],stage1_29[226]}
   );
   gpc606_5 gpc1276 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[137],stage1_31[144],stage1_30[156],stage1_29[227]}
   );
   gpc606_5 gpc1277 (
      {stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[138],stage1_31[145],stage1_30[157],stage1_29[228]}
   );
   gpc606_5 gpc1278 (
      {stage0_29[443], stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[139],stage1_31[146],stage1_30[158],stage1_29[229]}
   );
   gpc606_5 gpc1279 (
      {stage0_29[449], stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[140],stage1_31[147],stage1_30[159],stage1_29[230]}
   );
   gpc606_5 gpc1280 (
      {stage0_29[455], stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[141],stage1_31[148],stage1_30[160],stage1_29[231]}
   );
   gpc606_5 gpc1281 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[142],stage1_31[149],stage1_30[161],stage1_29[232]}
   );
   gpc606_5 gpc1282 (
      {stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[143],stage1_31[150],stage1_30[162],stage1_29[233]}
   );
   gpc606_5 gpc1283 (
      {stage0_29[473], stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[144],stage1_31[151],stage1_30[163],stage1_29[234]}
   );
   gpc606_5 gpc1284 (
      {stage0_29[479], stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[145],stage1_31[152],stage1_30[164],stage1_29[235]}
   );
   gpc606_5 gpc1285 (
      {stage0_29[485], stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[146],stage1_31[153],stage1_30[165],stage1_29[236]}
   );
   gpc606_5 gpc1286 (
      {stage0_29[491], stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[147],stage1_31[154],stage1_30[166],stage1_29[237]}
   );
   gpc606_5 gpc1287 (
      {stage0_29[497], stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[148],stage1_31[155],stage1_30[167],stage1_29[238]}
   );
   gpc606_5 gpc1288 (
      {stage0_29[503], stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[149],stage1_31[156],stage1_30[168],stage1_29[239]}
   );
   gpc1_1 gpc1289 (
      {stage0_0[502]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1290 (
      {stage0_0[503]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1291 (
      {stage0_0[504]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1292 (
      {stage0_0[505]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1293 (
      {stage0_0[506]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1294 (
      {stage0_0[507]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1295 (
      {stage0_0[508]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1296 (
      {stage0_0[509]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1297 (
      {stage0_0[510]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1298 (
      {stage0_0[511]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1299 (
      {stage0_1[453]},
      {stage1_1[140]}
   );
   gpc1_1 gpc1300 (
      {stage0_1[454]},
      {stage1_1[141]}
   );
   gpc1_1 gpc1301 (
      {stage0_1[455]},
      {stage1_1[142]}
   );
   gpc1_1 gpc1302 (
      {stage0_1[456]},
      {stage1_1[143]}
   );
   gpc1_1 gpc1303 (
      {stage0_1[457]},
      {stage1_1[144]}
   );
   gpc1_1 gpc1304 (
      {stage0_1[458]},
      {stage1_1[145]}
   );
   gpc1_1 gpc1305 (
      {stage0_1[459]},
      {stage1_1[146]}
   );
   gpc1_1 gpc1306 (
      {stage0_1[460]},
      {stage1_1[147]}
   );
   gpc1_1 gpc1307 (
      {stage0_1[461]},
      {stage1_1[148]}
   );
   gpc1_1 gpc1308 (
      {stage0_1[462]},
      {stage1_1[149]}
   );
   gpc1_1 gpc1309 (
      {stage0_1[463]},
      {stage1_1[150]}
   );
   gpc1_1 gpc1310 (
      {stage0_1[464]},
      {stage1_1[151]}
   );
   gpc1_1 gpc1311 (
      {stage0_1[465]},
      {stage1_1[152]}
   );
   gpc1_1 gpc1312 (
      {stage0_1[466]},
      {stage1_1[153]}
   );
   gpc1_1 gpc1313 (
      {stage0_1[467]},
      {stage1_1[154]}
   );
   gpc1_1 gpc1314 (
      {stage0_1[468]},
      {stage1_1[155]}
   );
   gpc1_1 gpc1315 (
      {stage0_1[469]},
      {stage1_1[156]}
   );
   gpc1_1 gpc1316 (
      {stage0_1[470]},
      {stage1_1[157]}
   );
   gpc1_1 gpc1317 (
      {stage0_1[471]},
      {stage1_1[158]}
   );
   gpc1_1 gpc1318 (
      {stage0_1[472]},
      {stage1_1[159]}
   );
   gpc1_1 gpc1319 (
      {stage0_1[473]},
      {stage1_1[160]}
   );
   gpc1_1 gpc1320 (
      {stage0_1[474]},
      {stage1_1[161]}
   );
   gpc1_1 gpc1321 (
      {stage0_1[475]},
      {stage1_1[162]}
   );
   gpc1_1 gpc1322 (
      {stage0_1[476]},
      {stage1_1[163]}
   );
   gpc1_1 gpc1323 (
      {stage0_1[477]},
      {stage1_1[164]}
   );
   gpc1_1 gpc1324 (
      {stage0_1[478]},
      {stage1_1[165]}
   );
   gpc1_1 gpc1325 (
      {stage0_1[479]},
      {stage1_1[166]}
   );
   gpc1_1 gpc1326 (
      {stage0_1[480]},
      {stage1_1[167]}
   );
   gpc1_1 gpc1327 (
      {stage0_1[481]},
      {stage1_1[168]}
   );
   gpc1_1 gpc1328 (
      {stage0_1[482]},
      {stage1_1[169]}
   );
   gpc1_1 gpc1329 (
      {stage0_1[483]},
      {stage1_1[170]}
   );
   gpc1_1 gpc1330 (
      {stage0_1[484]},
      {stage1_1[171]}
   );
   gpc1_1 gpc1331 (
      {stage0_1[485]},
      {stage1_1[172]}
   );
   gpc1_1 gpc1332 (
      {stage0_1[486]},
      {stage1_1[173]}
   );
   gpc1_1 gpc1333 (
      {stage0_1[487]},
      {stage1_1[174]}
   );
   gpc1_1 gpc1334 (
      {stage0_1[488]},
      {stage1_1[175]}
   );
   gpc1_1 gpc1335 (
      {stage0_1[489]},
      {stage1_1[176]}
   );
   gpc1_1 gpc1336 (
      {stage0_1[490]},
      {stage1_1[177]}
   );
   gpc1_1 gpc1337 (
      {stage0_1[491]},
      {stage1_1[178]}
   );
   gpc1_1 gpc1338 (
      {stage0_1[492]},
      {stage1_1[179]}
   );
   gpc1_1 gpc1339 (
      {stage0_1[493]},
      {stage1_1[180]}
   );
   gpc1_1 gpc1340 (
      {stage0_1[494]},
      {stage1_1[181]}
   );
   gpc1_1 gpc1341 (
      {stage0_1[495]},
      {stage1_1[182]}
   );
   gpc1_1 gpc1342 (
      {stage0_1[496]},
      {stage1_1[183]}
   );
   gpc1_1 gpc1343 (
      {stage0_1[497]},
      {stage1_1[184]}
   );
   gpc1_1 gpc1344 (
      {stage0_1[498]},
      {stage1_1[185]}
   );
   gpc1_1 gpc1345 (
      {stage0_1[499]},
      {stage1_1[186]}
   );
   gpc1_1 gpc1346 (
      {stage0_1[500]},
      {stage1_1[187]}
   );
   gpc1_1 gpc1347 (
      {stage0_1[501]},
      {stage1_1[188]}
   );
   gpc1_1 gpc1348 (
      {stage0_1[502]},
      {stage1_1[189]}
   );
   gpc1_1 gpc1349 (
      {stage0_1[503]},
      {stage1_1[190]}
   );
   gpc1_1 gpc1350 (
      {stage0_1[504]},
      {stage1_1[191]}
   );
   gpc1_1 gpc1351 (
      {stage0_1[505]},
      {stage1_1[192]}
   );
   gpc1_1 gpc1352 (
      {stage0_1[506]},
      {stage1_1[193]}
   );
   gpc1_1 gpc1353 (
      {stage0_1[507]},
      {stage1_1[194]}
   );
   gpc1_1 gpc1354 (
      {stage0_1[508]},
      {stage1_1[195]}
   );
   gpc1_1 gpc1355 (
      {stage0_1[509]},
      {stage1_1[196]}
   );
   gpc1_1 gpc1356 (
      {stage0_1[510]},
      {stage1_1[197]}
   );
   gpc1_1 gpc1357 (
      {stage0_1[511]},
      {stage1_1[198]}
   );
   gpc1_1 gpc1358 (
      {stage0_2[481]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1359 (
      {stage0_2[482]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1360 (
      {stage0_2[483]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1361 (
      {stage0_2[484]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1362 (
      {stage0_2[485]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1363 (
      {stage0_2[486]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1364 (
      {stage0_2[487]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1365 (
      {stage0_2[488]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1366 (
      {stage0_2[489]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1367 (
      {stage0_2[490]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1368 (
      {stage0_2[491]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1369 (
      {stage0_2[492]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1370 (
      {stage0_2[493]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1371 (
      {stage0_2[494]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1372 (
      {stage0_2[495]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1373 (
      {stage0_2[496]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1374 (
      {stage0_2[497]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1375 (
      {stage0_2[498]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1376 (
      {stage0_2[499]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1377 (
      {stage0_2[500]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1378 (
      {stage0_2[501]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1379 (
      {stage0_2[502]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1380 (
      {stage0_2[503]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1381 (
      {stage0_2[504]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1382 (
      {stage0_2[505]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1383 (
      {stage0_2[506]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1384 (
      {stage0_2[507]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1385 (
      {stage0_2[508]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1386 (
      {stage0_2[509]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1387 (
      {stage0_2[510]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1388 (
      {stage0_2[511]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1389 (
      {stage0_3[414]},
      {stage1_3[179]}
   );
   gpc1_1 gpc1390 (
      {stage0_3[415]},
      {stage1_3[180]}
   );
   gpc1_1 gpc1391 (
      {stage0_3[416]},
      {stage1_3[181]}
   );
   gpc1_1 gpc1392 (
      {stage0_3[417]},
      {stage1_3[182]}
   );
   gpc1_1 gpc1393 (
      {stage0_3[418]},
      {stage1_3[183]}
   );
   gpc1_1 gpc1394 (
      {stage0_3[419]},
      {stage1_3[184]}
   );
   gpc1_1 gpc1395 (
      {stage0_3[420]},
      {stage1_3[185]}
   );
   gpc1_1 gpc1396 (
      {stage0_3[421]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1397 (
      {stage0_3[422]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1398 (
      {stage0_3[423]},
      {stage1_3[188]}
   );
   gpc1_1 gpc1399 (
      {stage0_3[424]},
      {stage1_3[189]}
   );
   gpc1_1 gpc1400 (
      {stage0_3[425]},
      {stage1_3[190]}
   );
   gpc1_1 gpc1401 (
      {stage0_3[426]},
      {stage1_3[191]}
   );
   gpc1_1 gpc1402 (
      {stage0_3[427]},
      {stage1_3[192]}
   );
   gpc1_1 gpc1403 (
      {stage0_3[428]},
      {stage1_3[193]}
   );
   gpc1_1 gpc1404 (
      {stage0_3[429]},
      {stage1_3[194]}
   );
   gpc1_1 gpc1405 (
      {stage0_3[430]},
      {stage1_3[195]}
   );
   gpc1_1 gpc1406 (
      {stage0_3[431]},
      {stage1_3[196]}
   );
   gpc1_1 gpc1407 (
      {stage0_3[432]},
      {stage1_3[197]}
   );
   gpc1_1 gpc1408 (
      {stage0_3[433]},
      {stage1_3[198]}
   );
   gpc1_1 gpc1409 (
      {stage0_3[434]},
      {stage1_3[199]}
   );
   gpc1_1 gpc1410 (
      {stage0_3[435]},
      {stage1_3[200]}
   );
   gpc1_1 gpc1411 (
      {stage0_3[436]},
      {stage1_3[201]}
   );
   gpc1_1 gpc1412 (
      {stage0_3[437]},
      {stage1_3[202]}
   );
   gpc1_1 gpc1413 (
      {stage0_3[438]},
      {stage1_3[203]}
   );
   gpc1_1 gpc1414 (
      {stage0_3[439]},
      {stage1_3[204]}
   );
   gpc1_1 gpc1415 (
      {stage0_3[440]},
      {stage1_3[205]}
   );
   gpc1_1 gpc1416 (
      {stage0_3[441]},
      {stage1_3[206]}
   );
   gpc1_1 gpc1417 (
      {stage0_3[442]},
      {stage1_3[207]}
   );
   gpc1_1 gpc1418 (
      {stage0_3[443]},
      {stage1_3[208]}
   );
   gpc1_1 gpc1419 (
      {stage0_3[444]},
      {stage1_3[209]}
   );
   gpc1_1 gpc1420 (
      {stage0_3[445]},
      {stage1_3[210]}
   );
   gpc1_1 gpc1421 (
      {stage0_3[446]},
      {stage1_3[211]}
   );
   gpc1_1 gpc1422 (
      {stage0_3[447]},
      {stage1_3[212]}
   );
   gpc1_1 gpc1423 (
      {stage0_3[448]},
      {stage1_3[213]}
   );
   gpc1_1 gpc1424 (
      {stage0_3[449]},
      {stage1_3[214]}
   );
   gpc1_1 gpc1425 (
      {stage0_3[450]},
      {stage1_3[215]}
   );
   gpc1_1 gpc1426 (
      {stage0_3[451]},
      {stage1_3[216]}
   );
   gpc1_1 gpc1427 (
      {stage0_3[452]},
      {stage1_3[217]}
   );
   gpc1_1 gpc1428 (
      {stage0_3[453]},
      {stage1_3[218]}
   );
   gpc1_1 gpc1429 (
      {stage0_3[454]},
      {stage1_3[219]}
   );
   gpc1_1 gpc1430 (
      {stage0_3[455]},
      {stage1_3[220]}
   );
   gpc1_1 gpc1431 (
      {stage0_3[456]},
      {stage1_3[221]}
   );
   gpc1_1 gpc1432 (
      {stage0_3[457]},
      {stage1_3[222]}
   );
   gpc1_1 gpc1433 (
      {stage0_3[458]},
      {stage1_3[223]}
   );
   gpc1_1 gpc1434 (
      {stage0_3[459]},
      {stage1_3[224]}
   );
   gpc1_1 gpc1435 (
      {stage0_3[460]},
      {stage1_3[225]}
   );
   gpc1_1 gpc1436 (
      {stage0_3[461]},
      {stage1_3[226]}
   );
   gpc1_1 gpc1437 (
      {stage0_3[462]},
      {stage1_3[227]}
   );
   gpc1_1 gpc1438 (
      {stage0_3[463]},
      {stage1_3[228]}
   );
   gpc1_1 gpc1439 (
      {stage0_3[464]},
      {stage1_3[229]}
   );
   gpc1_1 gpc1440 (
      {stage0_3[465]},
      {stage1_3[230]}
   );
   gpc1_1 gpc1441 (
      {stage0_3[466]},
      {stage1_3[231]}
   );
   gpc1_1 gpc1442 (
      {stage0_3[467]},
      {stage1_3[232]}
   );
   gpc1_1 gpc1443 (
      {stage0_3[468]},
      {stage1_3[233]}
   );
   gpc1_1 gpc1444 (
      {stage0_3[469]},
      {stage1_3[234]}
   );
   gpc1_1 gpc1445 (
      {stage0_3[470]},
      {stage1_3[235]}
   );
   gpc1_1 gpc1446 (
      {stage0_3[471]},
      {stage1_3[236]}
   );
   gpc1_1 gpc1447 (
      {stage0_3[472]},
      {stage1_3[237]}
   );
   gpc1_1 gpc1448 (
      {stage0_3[473]},
      {stage1_3[238]}
   );
   gpc1_1 gpc1449 (
      {stage0_3[474]},
      {stage1_3[239]}
   );
   gpc1_1 gpc1450 (
      {stage0_3[475]},
      {stage1_3[240]}
   );
   gpc1_1 gpc1451 (
      {stage0_3[476]},
      {stage1_3[241]}
   );
   gpc1_1 gpc1452 (
      {stage0_3[477]},
      {stage1_3[242]}
   );
   gpc1_1 gpc1453 (
      {stage0_3[478]},
      {stage1_3[243]}
   );
   gpc1_1 gpc1454 (
      {stage0_3[479]},
      {stage1_3[244]}
   );
   gpc1_1 gpc1455 (
      {stage0_3[480]},
      {stage1_3[245]}
   );
   gpc1_1 gpc1456 (
      {stage0_3[481]},
      {stage1_3[246]}
   );
   gpc1_1 gpc1457 (
      {stage0_3[482]},
      {stage1_3[247]}
   );
   gpc1_1 gpc1458 (
      {stage0_3[483]},
      {stage1_3[248]}
   );
   gpc1_1 gpc1459 (
      {stage0_3[484]},
      {stage1_3[249]}
   );
   gpc1_1 gpc1460 (
      {stage0_3[485]},
      {stage1_3[250]}
   );
   gpc1_1 gpc1461 (
      {stage0_3[486]},
      {stage1_3[251]}
   );
   gpc1_1 gpc1462 (
      {stage0_3[487]},
      {stage1_3[252]}
   );
   gpc1_1 gpc1463 (
      {stage0_3[488]},
      {stage1_3[253]}
   );
   gpc1_1 gpc1464 (
      {stage0_3[489]},
      {stage1_3[254]}
   );
   gpc1_1 gpc1465 (
      {stage0_3[490]},
      {stage1_3[255]}
   );
   gpc1_1 gpc1466 (
      {stage0_3[491]},
      {stage1_3[256]}
   );
   gpc1_1 gpc1467 (
      {stage0_3[492]},
      {stage1_3[257]}
   );
   gpc1_1 gpc1468 (
      {stage0_3[493]},
      {stage1_3[258]}
   );
   gpc1_1 gpc1469 (
      {stage0_3[494]},
      {stage1_3[259]}
   );
   gpc1_1 gpc1470 (
      {stage0_3[495]},
      {stage1_3[260]}
   );
   gpc1_1 gpc1471 (
      {stage0_3[496]},
      {stage1_3[261]}
   );
   gpc1_1 gpc1472 (
      {stage0_3[497]},
      {stage1_3[262]}
   );
   gpc1_1 gpc1473 (
      {stage0_3[498]},
      {stage1_3[263]}
   );
   gpc1_1 gpc1474 (
      {stage0_3[499]},
      {stage1_3[264]}
   );
   gpc1_1 gpc1475 (
      {stage0_3[500]},
      {stage1_3[265]}
   );
   gpc1_1 gpc1476 (
      {stage0_3[501]},
      {stage1_3[266]}
   );
   gpc1_1 gpc1477 (
      {stage0_3[502]},
      {stage1_3[267]}
   );
   gpc1_1 gpc1478 (
      {stage0_3[503]},
      {stage1_3[268]}
   );
   gpc1_1 gpc1479 (
      {stage0_3[504]},
      {stage1_3[269]}
   );
   gpc1_1 gpc1480 (
      {stage0_3[505]},
      {stage1_3[270]}
   );
   gpc1_1 gpc1481 (
      {stage0_3[506]},
      {stage1_3[271]}
   );
   gpc1_1 gpc1482 (
      {stage0_3[507]},
      {stage1_3[272]}
   );
   gpc1_1 gpc1483 (
      {stage0_3[508]},
      {stage1_3[273]}
   );
   gpc1_1 gpc1484 (
      {stage0_3[509]},
      {stage1_3[274]}
   );
   gpc1_1 gpc1485 (
      {stage0_3[510]},
      {stage1_3[275]}
   );
   gpc1_1 gpc1486 (
      {stage0_3[511]},
      {stage1_3[276]}
   );
   gpc1_1 gpc1487 (
      {stage0_6[446]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1488 (
      {stage0_6[447]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1489 (
      {stage0_6[448]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1490 (
      {stage0_6[449]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1491 (
      {stage0_6[450]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1492 (
      {stage0_6[451]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1493 (
      {stage0_6[452]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1494 (
      {stage0_6[453]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1495 (
      {stage0_6[454]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1496 (
      {stage0_6[455]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1497 (
      {stage0_6[456]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1498 (
      {stage0_6[457]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1499 (
      {stage0_6[458]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1500 (
      {stage0_6[459]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1501 (
      {stage0_6[460]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1502 (
      {stage0_6[461]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1503 (
      {stage0_6[462]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1504 (
      {stage0_6[463]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1505 (
      {stage0_6[464]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1506 (
      {stage0_6[465]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1507 (
      {stage0_6[466]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1508 (
      {stage0_6[467]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1509 (
      {stage0_6[468]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1510 (
      {stage0_6[469]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1511 (
      {stage0_6[470]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1512 (
      {stage0_6[471]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1513 (
      {stage0_6[472]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1514 (
      {stage0_6[473]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1515 (
      {stage0_6[474]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1516 (
      {stage0_6[475]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1517 (
      {stage0_6[476]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1518 (
      {stage0_6[477]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1519 (
      {stage0_6[478]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1520 (
      {stage0_6[479]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1521 (
      {stage0_6[480]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1522 (
      {stage0_6[481]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1523 (
      {stage0_6[482]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1524 (
      {stage0_6[483]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1525 (
      {stage0_6[484]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1526 (
      {stage0_6[485]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1527 (
      {stage0_6[486]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1528 (
      {stage0_6[487]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1529 (
      {stage0_6[488]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1530 (
      {stage0_6[489]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1531 (
      {stage0_6[490]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1532 (
      {stage0_6[491]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1533 (
      {stage0_6[492]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1534 (
      {stage0_6[493]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1535 (
      {stage0_6[494]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1536 (
      {stage0_6[495]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1537 (
      {stage0_6[496]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1538 (
      {stage0_6[497]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1539 (
      {stage0_6[498]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1540 (
      {stage0_6[499]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1541 (
      {stage0_6[500]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1542 (
      {stage0_6[501]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1543 (
      {stage0_6[502]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1544 (
      {stage0_6[503]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1545 (
      {stage0_6[504]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1546 (
      {stage0_6[505]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1547 (
      {stage0_6[506]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1548 (
      {stage0_6[507]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1549 (
      {stage0_6[508]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1550 (
      {stage0_6[509]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1551 (
      {stage0_6[510]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1552 (
      {stage0_6[511]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1553 (
      {stage0_8[377]},
      {stage1_8[214]}
   );
   gpc1_1 gpc1554 (
      {stage0_8[378]},
      {stage1_8[215]}
   );
   gpc1_1 gpc1555 (
      {stage0_8[379]},
      {stage1_8[216]}
   );
   gpc1_1 gpc1556 (
      {stage0_8[380]},
      {stage1_8[217]}
   );
   gpc1_1 gpc1557 (
      {stage0_8[381]},
      {stage1_8[218]}
   );
   gpc1_1 gpc1558 (
      {stage0_8[382]},
      {stage1_8[219]}
   );
   gpc1_1 gpc1559 (
      {stage0_8[383]},
      {stage1_8[220]}
   );
   gpc1_1 gpc1560 (
      {stage0_8[384]},
      {stage1_8[221]}
   );
   gpc1_1 gpc1561 (
      {stage0_8[385]},
      {stage1_8[222]}
   );
   gpc1_1 gpc1562 (
      {stage0_8[386]},
      {stage1_8[223]}
   );
   gpc1_1 gpc1563 (
      {stage0_8[387]},
      {stage1_8[224]}
   );
   gpc1_1 gpc1564 (
      {stage0_8[388]},
      {stage1_8[225]}
   );
   gpc1_1 gpc1565 (
      {stage0_8[389]},
      {stage1_8[226]}
   );
   gpc1_1 gpc1566 (
      {stage0_8[390]},
      {stage1_8[227]}
   );
   gpc1_1 gpc1567 (
      {stage0_8[391]},
      {stage1_8[228]}
   );
   gpc1_1 gpc1568 (
      {stage0_8[392]},
      {stage1_8[229]}
   );
   gpc1_1 gpc1569 (
      {stage0_8[393]},
      {stage1_8[230]}
   );
   gpc1_1 gpc1570 (
      {stage0_8[394]},
      {stage1_8[231]}
   );
   gpc1_1 gpc1571 (
      {stage0_8[395]},
      {stage1_8[232]}
   );
   gpc1_1 gpc1572 (
      {stage0_8[396]},
      {stage1_8[233]}
   );
   gpc1_1 gpc1573 (
      {stage0_8[397]},
      {stage1_8[234]}
   );
   gpc1_1 gpc1574 (
      {stage0_8[398]},
      {stage1_8[235]}
   );
   gpc1_1 gpc1575 (
      {stage0_8[399]},
      {stage1_8[236]}
   );
   gpc1_1 gpc1576 (
      {stage0_8[400]},
      {stage1_8[237]}
   );
   gpc1_1 gpc1577 (
      {stage0_8[401]},
      {stage1_8[238]}
   );
   gpc1_1 gpc1578 (
      {stage0_8[402]},
      {stage1_8[239]}
   );
   gpc1_1 gpc1579 (
      {stage0_8[403]},
      {stage1_8[240]}
   );
   gpc1_1 gpc1580 (
      {stage0_8[404]},
      {stage1_8[241]}
   );
   gpc1_1 gpc1581 (
      {stage0_8[405]},
      {stage1_8[242]}
   );
   gpc1_1 gpc1582 (
      {stage0_8[406]},
      {stage1_8[243]}
   );
   gpc1_1 gpc1583 (
      {stage0_8[407]},
      {stage1_8[244]}
   );
   gpc1_1 gpc1584 (
      {stage0_8[408]},
      {stage1_8[245]}
   );
   gpc1_1 gpc1585 (
      {stage0_8[409]},
      {stage1_8[246]}
   );
   gpc1_1 gpc1586 (
      {stage0_8[410]},
      {stage1_8[247]}
   );
   gpc1_1 gpc1587 (
      {stage0_8[411]},
      {stage1_8[248]}
   );
   gpc1_1 gpc1588 (
      {stage0_8[412]},
      {stage1_8[249]}
   );
   gpc1_1 gpc1589 (
      {stage0_8[413]},
      {stage1_8[250]}
   );
   gpc1_1 gpc1590 (
      {stage0_8[414]},
      {stage1_8[251]}
   );
   gpc1_1 gpc1591 (
      {stage0_8[415]},
      {stage1_8[252]}
   );
   gpc1_1 gpc1592 (
      {stage0_8[416]},
      {stage1_8[253]}
   );
   gpc1_1 gpc1593 (
      {stage0_8[417]},
      {stage1_8[254]}
   );
   gpc1_1 gpc1594 (
      {stage0_8[418]},
      {stage1_8[255]}
   );
   gpc1_1 gpc1595 (
      {stage0_8[419]},
      {stage1_8[256]}
   );
   gpc1_1 gpc1596 (
      {stage0_8[420]},
      {stage1_8[257]}
   );
   gpc1_1 gpc1597 (
      {stage0_8[421]},
      {stage1_8[258]}
   );
   gpc1_1 gpc1598 (
      {stage0_8[422]},
      {stage1_8[259]}
   );
   gpc1_1 gpc1599 (
      {stage0_8[423]},
      {stage1_8[260]}
   );
   gpc1_1 gpc1600 (
      {stage0_8[424]},
      {stage1_8[261]}
   );
   gpc1_1 gpc1601 (
      {stage0_8[425]},
      {stage1_8[262]}
   );
   gpc1_1 gpc1602 (
      {stage0_8[426]},
      {stage1_8[263]}
   );
   gpc1_1 gpc1603 (
      {stage0_8[427]},
      {stage1_8[264]}
   );
   gpc1_1 gpc1604 (
      {stage0_8[428]},
      {stage1_8[265]}
   );
   gpc1_1 gpc1605 (
      {stage0_8[429]},
      {stage1_8[266]}
   );
   gpc1_1 gpc1606 (
      {stage0_8[430]},
      {stage1_8[267]}
   );
   gpc1_1 gpc1607 (
      {stage0_8[431]},
      {stage1_8[268]}
   );
   gpc1_1 gpc1608 (
      {stage0_8[432]},
      {stage1_8[269]}
   );
   gpc1_1 gpc1609 (
      {stage0_8[433]},
      {stage1_8[270]}
   );
   gpc1_1 gpc1610 (
      {stage0_8[434]},
      {stage1_8[271]}
   );
   gpc1_1 gpc1611 (
      {stage0_8[435]},
      {stage1_8[272]}
   );
   gpc1_1 gpc1612 (
      {stage0_8[436]},
      {stage1_8[273]}
   );
   gpc1_1 gpc1613 (
      {stage0_8[437]},
      {stage1_8[274]}
   );
   gpc1_1 gpc1614 (
      {stage0_8[438]},
      {stage1_8[275]}
   );
   gpc1_1 gpc1615 (
      {stage0_8[439]},
      {stage1_8[276]}
   );
   gpc1_1 gpc1616 (
      {stage0_8[440]},
      {stage1_8[277]}
   );
   gpc1_1 gpc1617 (
      {stage0_8[441]},
      {stage1_8[278]}
   );
   gpc1_1 gpc1618 (
      {stage0_8[442]},
      {stage1_8[279]}
   );
   gpc1_1 gpc1619 (
      {stage0_8[443]},
      {stage1_8[280]}
   );
   gpc1_1 gpc1620 (
      {stage0_8[444]},
      {stage1_8[281]}
   );
   gpc1_1 gpc1621 (
      {stage0_8[445]},
      {stage1_8[282]}
   );
   gpc1_1 gpc1622 (
      {stage0_8[446]},
      {stage1_8[283]}
   );
   gpc1_1 gpc1623 (
      {stage0_8[447]},
      {stage1_8[284]}
   );
   gpc1_1 gpc1624 (
      {stage0_8[448]},
      {stage1_8[285]}
   );
   gpc1_1 gpc1625 (
      {stage0_8[449]},
      {stage1_8[286]}
   );
   gpc1_1 gpc1626 (
      {stage0_8[450]},
      {stage1_8[287]}
   );
   gpc1_1 gpc1627 (
      {stage0_8[451]},
      {stage1_8[288]}
   );
   gpc1_1 gpc1628 (
      {stage0_8[452]},
      {stage1_8[289]}
   );
   gpc1_1 gpc1629 (
      {stage0_8[453]},
      {stage1_8[290]}
   );
   gpc1_1 gpc1630 (
      {stage0_8[454]},
      {stage1_8[291]}
   );
   gpc1_1 gpc1631 (
      {stage0_8[455]},
      {stage1_8[292]}
   );
   gpc1_1 gpc1632 (
      {stage0_8[456]},
      {stage1_8[293]}
   );
   gpc1_1 gpc1633 (
      {stage0_8[457]},
      {stage1_8[294]}
   );
   gpc1_1 gpc1634 (
      {stage0_8[458]},
      {stage1_8[295]}
   );
   gpc1_1 gpc1635 (
      {stage0_8[459]},
      {stage1_8[296]}
   );
   gpc1_1 gpc1636 (
      {stage0_8[460]},
      {stage1_8[297]}
   );
   gpc1_1 gpc1637 (
      {stage0_8[461]},
      {stage1_8[298]}
   );
   gpc1_1 gpc1638 (
      {stage0_8[462]},
      {stage1_8[299]}
   );
   gpc1_1 gpc1639 (
      {stage0_8[463]},
      {stage1_8[300]}
   );
   gpc1_1 gpc1640 (
      {stage0_8[464]},
      {stage1_8[301]}
   );
   gpc1_1 gpc1641 (
      {stage0_8[465]},
      {stage1_8[302]}
   );
   gpc1_1 gpc1642 (
      {stage0_8[466]},
      {stage1_8[303]}
   );
   gpc1_1 gpc1643 (
      {stage0_8[467]},
      {stage1_8[304]}
   );
   gpc1_1 gpc1644 (
      {stage0_8[468]},
      {stage1_8[305]}
   );
   gpc1_1 gpc1645 (
      {stage0_8[469]},
      {stage1_8[306]}
   );
   gpc1_1 gpc1646 (
      {stage0_8[470]},
      {stage1_8[307]}
   );
   gpc1_1 gpc1647 (
      {stage0_8[471]},
      {stage1_8[308]}
   );
   gpc1_1 gpc1648 (
      {stage0_8[472]},
      {stage1_8[309]}
   );
   gpc1_1 gpc1649 (
      {stage0_8[473]},
      {stage1_8[310]}
   );
   gpc1_1 gpc1650 (
      {stage0_8[474]},
      {stage1_8[311]}
   );
   gpc1_1 gpc1651 (
      {stage0_8[475]},
      {stage1_8[312]}
   );
   gpc1_1 gpc1652 (
      {stage0_8[476]},
      {stage1_8[313]}
   );
   gpc1_1 gpc1653 (
      {stage0_8[477]},
      {stage1_8[314]}
   );
   gpc1_1 gpc1654 (
      {stage0_8[478]},
      {stage1_8[315]}
   );
   gpc1_1 gpc1655 (
      {stage0_8[479]},
      {stage1_8[316]}
   );
   gpc1_1 gpc1656 (
      {stage0_8[480]},
      {stage1_8[317]}
   );
   gpc1_1 gpc1657 (
      {stage0_8[481]},
      {stage1_8[318]}
   );
   gpc1_1 gpc1658 (
      {stage0_8[482]},
      {stage1_8[319]}
   );
   gpc1_1 gpc1659 (
      {stage0_8[483]},
      {stage1_8[320]}
   );
   gpc1_1 gpc1660 (
      {stage0_8[484]},
      {stage1_8[321]}
   );
   gpc1_1 gpc1661 (
      {stage0_8[485]},
      {stage1_8[322]}
   );
   gpc1_1 gpc1662 (
      {stage0_8[486]},
      {stage1_8[323]}
   );
   gpc1_1 gpc1663 (
      {stage0_8[487]},
      {stage1_8[324]}
   );
   gpc1_1 gpc1664 (
      {stage0_8[488]},
      {stage1_8[325]}
   );
   gpc1_1 gpc1665 (
      {stage0_8[489]},
      {stage1_8[326]}
   );
   gpc1_1 gpc1666 (
      {stage0_8[490]},
      {stage1_8[327]}
   );
   gpc1_1 gpc1667 (
      {stage0_8[491]},
      {stage1_8[328]}
   );
   gpc1_1 gpc1668 (
      {stage0_8[492]},
      {stage1_8[329]}
   );
   gpc1_1 gpc1669 (
      {stage0_8[493]},
      {stage1_8[330]}
   );
   gpc1_1 gpc1670 (
      {stage0_8[494]},
      {stage1_8[331]}
   );
   gpc1_1 gpc1671 (
      {stage0_8[495]},
      {stage1_8[332]}
   );
   gpc1_1 gpc1672 (
      {stage0_8[496]},
      {stage1_8[333]}
   );
   gpc1_1 gpc1673 (
      {stage0_8[497]},
      {stage1_8[334]}
   );
   gpc1_1 gpc1674 (
      {stage0_8[498]},
      {stage1_8[335]}
   );
   gpc1_1 gpc1675 (
      {stage0_8[499]},
      {stage1_8[336]}
   );
   gpc1_1 gpc1676 (
      {stage0_8[500]},
      {stage1_8[337]}
   );
   gpc1_1 gpc1677 (
      {stage0_8[501]},
      {stage1_8[338]}
   );
   gpc1_1 gpc1678 (
      {stage0_8[502]},
      {stage1_8[339]}
   );
   gpc1_1 gpc1679 (
      {stage0_8[503]},
      {stage1_8[340]}
   );
   gpc1_1 gpc1680 (
      {stage0_8[504]},
      {stage1_8[341]}
   );
   gpc1_1 gpc1681 (
      {stage0_8[505]},
      {stage1_8[342]}
   );
   gpc1_1 gpc1682 (
      {stage0_8[506]},
      {stage1_8[343]}
   );
   gpc1_1 gpc1683 (
      {stage0_8[507]},
      {stage1_8[344]}
   );
   gpc1_1 gpc1684 (
      {stage0_8[508]},
      {stage1_8[345]}
   );
   gpc1_1 gpc1685 (
      {stage0_8[509]},
      {stage1_8[346]}
   );
   gpc1_1 gpc1686 (
      {stage0_8[510]},
      {stage1_8[347]}
   );
   gpc1_1 gpc1687 (
      {stage0_8[511]},
      {stage1_8[348]}
   );
   gpc1_1 gpc1688 (
      {stage0_9[509]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1689 (
      {stage0_9[510]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1690 (
      {stage0_9[511]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1691 (
      {stage0_11[501]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1692 (
      {stage0_11[502]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1693 (
      {stage0_11[503]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1694 (
      {stage0_11[504]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1695 (
      {stage0_11[505]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1696 (
      {stage0_11[506]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1697 (
      {stage0_11[507]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1698 (
      {stage0_11[508]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1699 (
      {stage0_11[509]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1700 (
      {stage0_11[510]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1701 (
      {stage0_11[511]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1702 (
      {stage0_13[507]},
      {stage1_13[227]}
   );
   gpc1_1 gpc1703 (
      {stage0_13[508]},
      {stage1_13[228]}
   );
   gpc1_1 gpc1704 (
      {stage0_13[509]},
      {stage1_13[229]}
   );
   gpc1_1 gpc1705 (
      {stage0_13[510]},
      {stage1_13[230]}
   );
   gpc1_1 gpc1706 (
      {stage0_13[511]},
      {stage1_13[231]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[472]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[473]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[474]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[475]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[476]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[477]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[478]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[479]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[480]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[481]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[482]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[483]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[484]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[485]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[486]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[487]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[488]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[489]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[490]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[491]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[492]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[493]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[494]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[495]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[496]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[497]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[498]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[499]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[500]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[501]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[502]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[503]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[504]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[505]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[506]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[507]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[508]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[509]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[510]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[511]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1747 (
      {stage0_15[456]},
      {stage1_15[181]}
   );
   gpc1_1 gpc1748 (
      {stage0_15[457]},
      {stage1_15[182]}
   );
   gpc1_1 gpc1749 (
      {stage0_15[458]},
      {stage1_15[183]}
   );
   gpc1_1 gpc1750 (
      {stage0_15[459]},
      {stage1_15[184]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[460]},
      {stage1_15[185]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[461]},
      {stage1_15[186]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[462]},
      {stage1_15[187]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[463]},
      {stage1_15[188]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[464]},
      {stage1_15[189]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[465]},
      {stage1_15[190]}
   );
   gpc1_1 gpc1757 (
      {stage0_15[466]},
      {stage1_15[191]}
   );
   gpc1_1 gpc1758 (
      {stage0_15[467]},
      {stage1_15[192]}
   );
   gpc1_1 gpc1759 (
      {stage0_15[468]},
      {stage1_15[193]}
   );
   gpc1_1 gpc1760 (
      {stage0_15[469]},
      {stage1_15[194]}
   );
   gpc1_1 gpc1761 (
      {stage0_15[470]},
      {stage1_15[195]}
   );
   gpc1_1 gpc1762 (
      {stage0_15[471]},
      {stage1_15[196]}
   );
   gpc1_1 gpc1763 (
      {stage0_15[472]},
      {stage1_15[197]}
   );
   gpc1_1 gpc1764 (
      {stage0_15[473]},
      {stage1_15[198]}
   );
   gpc1_1 gpc1765 (
      {stage0_15[474]},
      {stage1_15[199]}
   );
   gpc1_1 gpc1766 (
      {stage0_15[475]},
      {stage1_15[200]}
   );
   gpc1_1 gpc1767 (
      {stage0_15[476]},
      {stage1_15[201]}
   );
   gpc1_1 gpc1768 (
      {stage0_15[477]},
      {stage1_15[202]}
   );
   gpc1_1 gpc1769 (
      {stage0_15[478]},
      {stage1_15[203]}
   );
   gpc1_1 gpc1770 (
      {stage0_15[479]},
      {stage1_15[204]}
   );
   gpc1_1 gpc1771 (
      {stage0_15[480]},
      {stage1_15[205]}
   );
   gpc1_1 gpc1772 (
      {stage0_15[481]},
      {stage1_15[206]}
   );
   gpc1_1 gpc1773 (
      {stage0_15[482]},
      {stage1_15[207]}
   );
   gpc1_1 gpc1774 (
      {stage0_15[483]},
      {stage1_15[208]}
   );
   gpc1_1 gpc1775 (
      {stage0_15[484]},
      {stage1_15[209]}
   );
   gpc1_1 gpc1776 (
      {stage0_15[485]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1777 (
      {stage0_15[486]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1778 (
      {stage0_15[487]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1779 (
      {stage0_15[488]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1780 (
      {stage0_15[489]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1781 (
      {stage0_15[490]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1782 (
      {stage0_15[491]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1783 (
      {stage0_15[492]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1784 (
      {stage0_15[493]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1785 (
      {stage0_15[494]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1786 (
      {stage0_15[495]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1787 (
      {stage0_15[496]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1788 (
      {stage0_15[497]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1789 (
      {stage0_15[498]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1790 (
      {stage0_15[499]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1791 (
      {stage0_15[500]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1792 (
      {stage0_15[501]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1793 (
      {stage0_15[502]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1794 (
      {stage0_15[503]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1795 (
      {stage0_15[504]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1796 (
      {stage0_15[505]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1797 (
      {stage0_15[506]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1798 (
      {stage0_15[507]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1799 (
      {stage0_15[508]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1800 (
      {stage0_15[509]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1801 (
      {stage0_15[510]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1802 (
      {stage0_15[511]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1803 (
      {stage0_17[510]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1804 (
      {stage0_17[511]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1805 (
      {stage0_18[511]},
      {stage1_18[202]}
   );
   gpc1_1 gpc1806 (
      {stage0_19[431]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1807 (
      {stage0_19[432]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1808 (
      {stage0_19[433]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1809 (
      {stage0_19[434]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1810 (
      {stage0_19[435]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1811 (
      {stage0_19[436]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1812 (
      {stage0_19[437]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1813 (
      {stage0_19[438]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1814 (
      {stage0_19[439]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1815 (
      {stage0_19[440]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1816 (
      {stage0_19[441]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1817 (
      {stage0_19[442]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1818 (
      {stage0_19[443]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1819 (
      {stage0_19[444]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1820 (
      {stage0_19[445]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1821 (
      {stage0_19[446]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1822 (
      {stage0_19[447]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1823 (
      {stage0_19[448]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1824 (
      {stage0_19[449]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1825 (
      {stage0_19[450]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1826 (
      {stage0_19[451]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1827 (
      {stage0_19[452]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1828 (
      {stage0_19[453]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1829 (
      {stage0_19[454]},
      {stage1_19[205]}
   );
   gpc1_1 gpc1830 (
      {stage0_19[455]},
      {stage1_19[206]}
   );
   gpc1_1 gpc1831 (
      {stage0_19[456]},
      {stage1_19[207]}
   );
   gpc1_1 gpc1832 (
      {stage0_19[457]},
      {stage1_19[208]}
   );
   gpc1_1 gpc1833 (
      {stage0_19[458]},
      {stage1_19[209]}
   );
   gpc1_1 gpc1834 (
      {stage0_19[459]},
      {stage1_19[210]}
   );
   gpc1_1 gpc1835 (
      {stage0_19[460]},
      {stage1_19[211]}
   );
   gpc1_1 gpc1836 (
      {stage0_19[461]},
      {stage1_19[212]}
   );
   gpc1_1 gpc1837 (
      {stage0_19[462]},
      {stage1_19[213]}
   );
   gpc1_1 gpc1838 (
      {stage0_19[463]},
      {stage1_19[214]}
   );
   gpc1_1 gpc1839 (
      {stage0_19[464]},
      {stage1_19[215]}
   );
   gpc1_1 gpc1840 (
      {stage0_19[465]},
      {stage1_19[216]}
   );
   gpc1_1 gpc1841 (
      {stage0_19[466]},
      {stage1_19[217]}
   );
   gpc1_1 gpc1842 (
      {stage0_19[467]},
      {stage1_19[218]}
   );
   gpc1_1 gpc1843 (
      {stage0_19[468]},
      {stage1_19[219]}
   );
   gpc1_1 gpc1844 (
      {stage0_19[469]},
      {stage1_19[220]}
   );
   gpc1_1 gpc1845 (
      {stage0_19[470]},
      {stage1_19[221]}
   );
   gpc1_1 gpc1846 (
      {stage0_19[471]},
      {stage1_19[222]}
   );
   gpc1_1 gpc1847 (
      {stage0_19[472]},
      {stage1_19[223]}
   );
   gpc1_1 gpc1848 (
      {stage0_19[473]},
      {stage1_19[224]}
   );
   gpc1_1 gpc1849 (
      {stage0_19[474]},
      {stage1_19[225]}
   );
   gpc1_1 gpc1850 (
      {stage0_19[475]},
      {stage1_19[226]}
   );
   gpc1_1 gpc1851 (
      {stage0_19[476]},
      {stage1_19[227]}
   );
   gpc1_1 gpc1852 (
      {stage0_19[477]},
      {stage1_19[228]}
   );
   gpc1_1 gpc1853 (
      {stage0_19[478]},
      {stage1_19[229]}
   );
   gpc1_1 gpc1854 (
      {stage0_19[479]},
      {stage1_19[230]}
   );
   gpc1_1 gpc1855 (
      {stage0_19[480]},
      {stage1_19[231]}
   );
   gpc1_1 gpc1856 (
      {stage0_19[481]},
      {stage1_19[232]}
   );
   gpc1_1 gpc1857 (
      {stage0_19[482]},
      {stage1_19[233]}
   );
   gpc1_1 gpc1858 (
      {stage0_19[483]},
      {stage1_19[234]}
   );
   gpc1_1 gpc1859 (
      {stage0_19[484]},
      {stage1_19[235]}
   );
   gpc1_1 gpc1860 (
      {stage0_19[485]},
      {stage1_19[236]}
   );
   gpc1_1 gpc1861 (
      {stage0_19[486]},
      {stage1_19[237]}
   );
   gpc1_1 gpc1862 (
      {stage0_19[487]},
      {stage1_19[238]}
   );
   gpc1_1 gpc1863 (
      {stage0_19[488]},
      {stage1_19[239]}
   );
   gpc1_1 gpc1864 (
      {stage0_19[489]},
      {stage1_19[240]}
   );
   gpc1_1 gpc1865 (
      {stage0_19[490]},
      {stage1_19[241]}
   );
   gpc1_1 gpc1866 (
      {stage0_19[491]},
      {stage1_19[242]}
   );
   gpc1_1 gpc1867 (
      {stage0_19[492]},
      {stage1_19[243]}
   );
   gpc1_1 gpc1868 (
      {stage0_19[493]},
      {stage1_19[244]}
   );
   gpc1_1 gpc1869 (
      {stage0_19[494]},
      {stage1_19[245]}
   );
   gpc1_1 gpc1870 (
      {stage0_19[495]},
      {stage1_19[246]}
   );
   gpc1_1 gpc1871 (
      {stage0_19[496]},
      {stage1_19[247]}
   );
   gpc1_1 gpc1872 (
      {stage0_19[497]},
      {stage1_19[248]}
   );
   gpc1_1 gpc1873 (
      {stage0_19[498]},
      {stage1_19[249]}
   );
   gpc1_1 gpc1874 (
      {stage0_19[499]},
      {stage1_19[250]}
   );
   gpc1_1 gpc1875 (
      {stage0_19[500]},
      {stage1_19[251]}
   );
   gpc1_1 gpc1876 (
      {stage0_19[501]},
      {stage1_19[252]}
   );
   gpc1_1 gpc1877 (
      {stage0_19[502]},
      {stage1_19[253]}
   );
   gpc1_1 gpc1878 (
      {stage0_19[503]},
      {stage1_19[254]}
   );
   gpc1_1 gpc1879 (
      {stage0_19[504]},
      {stage1_19[255]}
   );
   gpc1_1 gpc1880 (
      {stage0_19[505]},
      {stage1_19[256]}
   );
   gpc1_1 gpc1881 (
      {stage0_19[506]},
      {stage1_19[257]}
   );
   gpc1_1 gpc1882 (
      {stage0_19[507]},
      {stage1_19[258]}
   );
   gpc1_1 gpc1883 (
      {stage0_19[508]},
      {stage1_19[259]}
   );
   gpc1_1 gpc1884 (
      {stage0_19[509]},
      {stage1_19[260]}
   );
   gpc1_1 gpc1885 (
      {stage0_19[510]},
      {stage1_19[261]}
   );
   gpc1_1 gpc1886 (
      {stage0_19[511]},
      {stage1_19[262]}
   );
   gpc1_1 gpc1887 (
      {stage0_20[504]},
      {stage1_20[206]}
   );
   gpc1_1 gpc1888 (
      {stage0_20[505]},
      {stage1_20[207]}
   );
   gpc1_1 gpc1889 (
      {stage0_20[506]},
      {stage1_20[208]}
   );
   gpc1_1 gpc1890 (
      {stage0_20[507]},
      {stage1_20[209]}
   );
   gpc1_1 gpc1891 (
      {stage0_20[508]},
      {stage1_20[210]}
   );
   gpc1_1 gpc1892 (
      {stage0_20[509]},
      {stage1_20[211]}
   );
   gpc1_1 gpc1893 (
      {stage0_20[510]},
      {stage1_20[212]}
   );
   gpc1_1 gpc1894 (
      {stage0_20[511]},
      {stage1_20[213]}
   );
   gpc1_1 gpc1895 (
      {stage0_21[471]},
      {stage1_21[229]}
   );
   gpc1_1 gpc1896 (
      {stage0_21[472]},
      {stage1_21[230]}
   );
   gpc1_1 gpc1897 (
      {stage0_21[473]},
      {stage1_21[231]}
   );
   gpc1_1 gpc1898 (
      {stage0_21[474]},
      {stage1_21[232]}
   );
   gpc1_1 gpc1899 (
      {stage0_21[475]},
      {stage1_21[233]}
   );
   gpc1_1 gpc1900 (
      {stage0_21[476]},
      {stage1_21[234]}
   );
   gpc1_1 gpc1901 (
      {stage0_21[477]},
      {stage1_21[235]}
   );
   gpc1_1 gpc1902 (
      {stage0_21[478]},
      {stage1_21[236]}
   );
   gpc1_1 gpc1903 (
      {stage0_21[479]},
      {stage1_21[237]}
   );
   gpc1_1 gpc1904 (
      {stage0_21[480]},
      {stage1_21[238]}
   );
   gpc1_1 gpc1905 (
      {stage0_21[481]},
      {stage1_21[239]}
   );
   gpc1_1 gpc1906 (
      {stage0_21[482]},
      {stage1_21[240]}
   );
   gpc1_1 gpc1907 (
      {stage0_21[483]},
      {stage1_21[241]}
   );
   gpc1_1 gpc1908 (
      {stage0_21[484]},
      {stage1_21[242]}
   );
   gpc1_1 gpc1909 (
      {stage0_21[485]},
      {stage1_21[243]}
   );
   gpc1_1 gpc1910 (
      {stage0_21[486]},
      {stage1_21[244]}
   );
   gpc1_1 gpc1911 (
      {stage0_21[487]},
      {stage1_21[245]}
   );
   gpc1_1 gpc1912 (
      {stage0_21[488]},
      {stage1_21[246]}
   );
   gpc1_1 gpc1913 (
      {stage0_21[489]},
      {stage1_21[247]}
   );
   gpc1_1 gpc1914 (
      {stage0_21[490]},
      {stage1_21[248]}
   );
   gpc1_1 gpc1915 (
      {stage0_21[491]},
      {stage1_21[249]}
   );
   gpc1_1 gpc1916 (
      {stage0_21[492]},
      {stage1_21[250]}
   );
   gpc1_1 gpc1917 (
      {stage0_21[493]},
      {stage1_21[251]}
   );
   gpc1_1 gpc1918 (
      {stage0_21[494]},
      {stage1_21[252]}
   );
   gpc1_1 gpc1919 (
      {stage0_21[495]},
      {stage1_21[253]}
   );
   gpc1_1 gpc1920 (
      {stage0_21[496]},
      {stage1_21[254]}
   );
   gpc1_1 gpc1921 (
      {stage0_21[497]},
      {stage1_21[255]}
   );
   gpc1_1 gpc1922 (
      {stage0_21[498]},
      {stage1_21[256]}
   );
   gpc1_1 gpc1923 (
      {stage0_21[499]},
      {stage1_21[257]}
   );
   gpc1_1 gpc1924 (
      {stage0_21[500]},
      {stage1_21[258]}
   );
   gpc1_1 gpc1925 (
      {stage0_21[501]},
      {stage1_21[259]}
   );
   gpc1_1 gpc1926 (
      {stage0_21[502]},
      {stage1_21[260]}
   );
   gpc1_1 gpc1927 (
      {stage0_21[503]},
      {stage1_21[261]}
   );
   gpc1_1 gpc1928 (
      {stage0_21[504]},
      {stage1_21[262]}
   );
   gpc1_1 gpc1929 (
      {stage0_21[505]},
      {stage1_21[263]}
   );
   gpc1_1 gpc1930 (
      {stage0_21[506]},
      {stage1_21[264]}
   );
   gpc1_1 gpc1931 (
      {stage0_21[507]},
      {stage1_21[265]}
   );
   gpc1_1 gpc1932 (
      {stage0_21[508]},
      {stage1_21[266]}
   );
   gpc1_1 gpc1933 (
      {stage0_21[509]},
      {stage1_21[267]}
   );
   gpc1_1 gpc1934 (
      {stage0_21[510]},
      {stage1_21[268]}
   );
   gpc1_1 gpc1935 (
      {stage0_21[511]},
      {stage1_21[269]}
   );
   gpc1_1 gpc1936 (
      {stage0_22[423]},
      {stage1_22[185]}
   );
   gpc1_1 gpc1937 (
      {stage0_22[424]},
      {stage1_22[186]}
   );
   gpc1_1 gpc1938 (
      {stage0_22[425]},
      {stage1_22[187]}
   );
   gpc1_1 gpc1939 (
      {stage0_22[426]},
      {stage1_22[188]}
   );
   gpc1_1 gpc1940 (
      {stage0_22[427]},
      {stage1_22[189]}
   );
   gpc1_1 gpc1941 (
      {stage0_22[428]},
      {stage1_22[190]}
   );
   gpc1_1 gpc1942 (
      {stage0_22[429]},
      {stage1_22[191]}
   );
   gpc1_1 gpc1943 (
      {stage0_22[430]},
      {stage1_22[192]}
   );
   gpc1_1 gpc1944 (
      {stage0_22[431]},
      {stage1_22[193]}
   );
   gpc1_1 gpc1945 (
      {stage0_22[432]},
      {stage1_22[194]}
   );
   gpc1_1 gpc1946 (
      {stage0_22[433]},
      {stage1_22[195]}
   );
   gpc1_1 gpc1947 (
      {stage0_22[434]},
      {stage1_22[196]}
   );
   gpc1_1 gpc1948 (
      {stage0_22[435]},
      {stage1_22[197]}
   );
   gpc1_1 gpc1949 (
      {stage0_22[436]},
      {stage1_22[198]}
   );
   gpc1_1 gpc1950 (
      {stage0_22[437]},
      {stage1_22[199]}
   );
   gpc1_1 gpc1951 (
      {stage0_22[438]},
      {stage1_22[200]}
   );
   gpc1_1 gpc1952 (
      {stage0_22[439]},
      {stage1_22[201]}
   );
   gpc1_1 gpc1953 (
      {stage0_22[440]},
      {stage1_22[202]}
   );
   gpc1_1 gpc1954 (
      {stage0_22[441]},
      {stage1_22[203]}
   );
   gpc1_1 gpc1955 (
      {stage0_22[442]},
      {stage1_22[204]}
   );
   gpc1_1 gpc1956 (
      {stage0_22[443]},
      {stage1_22[205]}
   );
   gpc1_1 gpc1957 (
      {stage0_22[444]},
      {stage1_22[206]}
   );
   gpc1_1 gpc1958 (
      {stage0_22[445]},
      {stage1_22[207]}
   );
   gpc1_1 gpc1959 (
      {stage0_22[446]},
      {stage1_22[208]}
   );
   gpc1_1 gpc1960 (
      {stage0_22[447]},
      {stage1_22[209]}
   );
   gpc1_1 gpc1961 (
      {stage0_22[448]},
      {stage1_22[210]}
   );
   gpc1_1 gpc1962 (
      {stage0_22[449]},
      {stage1_22[211]}
   );
   gpc1_1 gpc1963 (
      {stage0_22[450]},
      {stage1_22[212]}
   );
   gpc1_1 gpc1964 (
      {stage0_22[451]},
      {stage1_22[213]}
   );
   gpc1_1 gpc1965 (
      {stage0_22[452]},
      {stage1_22[214]}
   );
   gpc1_1 gpc1966 (
      {stage0_22[453]},
      {stage1_22[215]}
   );
   gpc1_1 gpc1967 (
      {stage0_22[454]},
      {stage1_22[216]}
   );
   gpc1_1 gpc1968 (
      {stage0_22[455]},
      {stage1_22[217]}
   );
   gpc1_1 gpc1969 (
      {stage0_22[456]},
      {stage1_22[218]}
   );
   gpc1_1 gpc1970 (
      {stage0_22[457]},
      {stage1_22[219]}
   );
   gpc1_1 gpc1971 (
      {stage0_22[458]},
      {stage1_22[220]}
   );
   gpc1_1 gpc1972 (
      {stage0_22[459]},
      {stage1_22[221]}
   );
   gpc1_1 gpc1973 (
      {stage0_22[460]},
      {stage1_22[222]}
   );
   gpc1_1 gpc1974 (
      {stage0_22[461]},
      {stage1_22[223]}
   );
   gpc1_1 gpc1975 (
      {stage0_22[462]},
      {stage1_22[224]}
   );
   gpc1_1 gpc1976 (
      {stage0_22[463]},
      {stage1_22[225]}
   );
   gpc1_1 gpc1977 (
      {stage0_22[464]},
      {stage1_22[226]}
   );
   gpc1_1 gpc1978 (
      {stage0_22[465]},
      {stage1_22[227]}
   );
   gpc1_1 gpc1979 (
      {stage0_22[466]},
      {stage1_22[228]}
   );
   gpc1_1 gpc1980 (
      {stage0_22[467]},
      {stage1_22[229]}
   );
   gpc1_1 gpc1981 (
      {stage0_22[468]},
      {stage1_22[230]}
   );
   gpc1_1 gpc1982 (
      {stage0_22[469]},
      {stage1_22[231]}
   );
   gpc1_1 gpc1983 (
      {stage0_22[470]},
      {stage1_22[232]}
   );
   gpc1_1 gpc1984 (
      {stage0_22[471]},
      {stage1_22[233]}
   );
   gpc1_1 gpc1985 (
      {stage0_22[472]},
      {stage1_22[234]}
   );
   gpc1_1 gpc1986 (
      {stage0_22[473]},
      {stage1_22[235]}
   );
   gpc1_1 gpc1987 (
      {stage0_22[474]},
      {stage1_22[236]}
   );
   gpc1_1 gpc1988 (
      {stage0_22[475]},
      {stage1_22[237]}
   );
   gpc1_1 gpc1989 (
      {stage0_22[476]},
      {stage1_22[238]}
   );
   gpc1_1 gpc1990 (
      {stage0_22[477]},
      {stage1_22[239]}
   );
   gpc1_1 gpc1991 (
      {stage0_22[478]},
      {stage1_22[240]}
   );
   gpc1_1 gpc1992 (
      {stage0_22[479]},
      {stage1_22[241]}
   );
   gpc1_1 gpc1993 (
      {stage0_22[480]},
      {stage1_22[242]}
   );
   gpc1_1 gpc1994 (
      {stage0_22[481]},
      {stage1_22[243]}
   );
   gpc1_1 gpc1995 (
      {stage0_22[482]},
      {stage1_22[244]}
   );
   gpc1_1 gpc1996 (
      {stage0_22[483]},
      {stage1_22[245]}
   );
   gpc1_1 gpc1997 (
      {stage0_22[484]},
      {stage1_22[246]}
   );
   gpc1_1 gpc1998 (
      {stage0_22[485]},
      {stage1_22[247]}
   );
   gpc1_1 gpc1999 (
      {stage0_22[486]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2000 (
      {stage0_22[487]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2001 (
      {stage0_22[488]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2002 (
      {stage0_22[489]},
      {stage1_22[251]}
   );
   gpc1_1 gpc2003 (
      {stage0_22[490]},
      {stage1_22[252]}
   );
   gpc1_1 gpc2004 (
      {stage0_22[491]},
      {stage1_22[253]}
   );
   gpc1_1 gpc2005 (
      {stage0_22[492]},
      {stage1_22[254]}
   );
   gpc1_1 gpc2006 (
      {stage0_22[493]},
      {stage1_22[255]}
   );
   gpc1_1 gpc2007 (
      {stage0_22[494]},
      {stage1_22[256]}
   );
   gpc1_1 gpc2008 (
      {stage0_22[495]},
      {stage1_22[257]}
   );
   gpc1_1 gpc2009 (
      {stage0_22[496]},
      {stage1_22[258]}
   );
   gpc1_1 gpc2010 (
      {stage0_22[497]},
      {stage1_22[259]}
   );
   gpc1_1 gpc2011 (
      {stage0_22[498]},
      {stage1_22[260]}
   );
   gpc1_1 gpc2012 (
      {stage0_22[499]},
      {stage1_22[261]}
   );
   gpc1_1 gpc2013 (
      {stage0_22[500]},
      {stage1_22[262]}
   );
   gpc1_1 gpc2014 (
      {stage0_22[501]},
      {stage1_22[263]}
   );
   gpc1_1 gpc2015 (
      {stage0_22[502]},
      {stage1_22[264]}
   );
   gpc1_1 gpc2016 (
      {stage0_22[503]},
      {stage1_22[265]}
   );
   gpc1_1 gpc2017 (
      {stage0_22[504]},
      {stage1_22[266]}
   );
   gpc1_1 gpc2018 (
      {stage0_22[505]},
      {stage1_22[267]}
   );
   gpc1_1 gpc2019 (
      {stage0_22[506]},
      {stage1_22[268]}
   );
   gpc1_1 gpc2020 (
      {stage0_22[507]},
      {stage1_22[269]}
   );
   gpc1_1 gpc2021 (
      {stage0_22[508]},
      {stage1_22[270]}
   );
   gpc1_1 gpc2022 (
      {stage0_22[509]},
      {stage1_22[271]}
   );
   gpc1_1 gpc2023 (
      {stage0_22[510]},
      {stage1_22[272]}
   );
   gpc1_1 gpc2024 (
      {stage0_22[511]},
      {stage1_22[273]}
   );
   gpc1_1 gpc2025 (
      {stage0_23[500]},
      {stage1_23[154]}
   );
   gpc1_1 gpc2026 (
      {stage0_23[501]},
      {stage1_23[155]}
   );
   gpc1_1 gpc2027 (
      {stage0_23[502]},
      {stage1_23[156]}
   );
   gpc1_1 gpc2028 (
      {stage0_23[503]},
      {stage1_23[157]}
   );
   gpc1_1 gpc2029 (
      {stage0_23[504]},
      {stage1_23[158]}
   );
   gpc1_1 gpc2030 (
      {stage0_23[505]},
      {stage1_23[159]}
   );
   gpc1_1 gpc2031 (
      {stage0_23[506]},
      {stage1_23[160]}
   );
   gpc1_1 gpc2032 (
      {stage0_23[507]},
      {stage1_23[161]}
   );
   gpc1_1 gpc2033 (
      {stage0_23[508]},
      {stage1_23[162]}
   );
   gpc1_1 gpc2034 (
      {stage0_23[509]},
      {stage1_23[163]}
   );
   gpc1_1 gpc2035 (
      {stage0_23[510]},
      {stage1_23[164]}
   );
   gpc1_1 gpc2036 (
      {stage0_23[511]},
      {stage1_23[165]}
   );
   gpc1_1 gpc2037 (
      {stage0_25[482]},
      {stage1_25[244]}
   );
   gpc1_1 gpc2038 (
      {stage0_25[483]},
      {stage1_25[245]}
   );
   gpc1_1 gpc2039 (
      {stage0_25[484]},
      {stage1_25[246]}
   );
   gpc1_1 gpc2040 (
      {stage0_25[485]},
      {stage1_25[247]}
   );
   gpc1_1 gpc2041 (
      {stage0_25[486]},
      {stage1_25[248]}
   );
   gpc1_1 gpc2042 (
      {stage0_25[487]},
      {stage1_25[249]}
   );
   gpc1_1 gpc2043 (
      {stage0_25[488]},
      {stage1_25[250]}
   );
   gpc1_1 gpc2044 (
      {stage0_25[489]},
      {stage1_25[251]}
   );
   gpc1_1 gpc2045 (
      {stage0_25[490]},
      {stage1_25[252]}
   );
   gpc1_1 gpc2046 (
      {stage0_25[491]},
      {stage1_25[253]}
   );
   gpc1_1 gpc2047 (
      {stage0_25[492]},
      {stage1_25[254]}
   );
   gpc1_1 gpc2048 (
      {stage0_25[493]},
      {stage1_25[255]}
   );
   gpc1_1 gpc2049 (
      {stage0_25[494]},
      {stage1_25[256]}
   );
   gpc1_1 gpc2050 (
      {stage0_25[495]},
      {stage1_25[257]}
   );
   gpc1_1 gpc2051 (
      {stage0_25[496]},
      {stage1_25[258]}
   );
   gpc1_1 gpc2052 (
      {stage0_25[497]},
      {stage1_25[259]}
   );
   gpc1_1 gpc2053 (
      {stage0_25[498]},
      {stage1_25[260]}
   );
   gpc1_1 gpc2054 (
      {stage0_25[499]},
      {stage1_25[261]}
   );
   gpc1_1 gpc2055 (
      {stage0_25[500]},
      {stage1_25[262]}
   );
   gpc1_1 gpc2056 (
      {stage0_25[501]},
      {stage1_25[263]}
   );
   gpc1_1 gpc2057 (
      {stage0_25[502]},
      {stage1_25[264]}
   );
   gpc1_1 gpc2058 (
      {stage0_25[503]},
      {stage1_25[265]}
   );
   gpc1_1 gpc2059 (
      {stage0_25[504]},
      {stage1_25[266]}
   );
   gpc1_1 gpc2060 (
      {stage0_25[505]},
      {stage1_25[267]}
   );
   gpc1_1 gpc2061 (
      {stage0_25[506]},
      {stage1_25[268]}
   );
   gpc1_1 gpc2062 (
      {stage0_25[507]},
      {stage1_25[269]}
   );
   gpc1_1 gpc2063 (
      {stage0_25[508]},
      {stage1_25[270]}
   );
   gpc1_1 gpc2064 (
      {stage0_25[509]},
      {stage1_25[271]}
   );
   gpc1_1 gpc2065 (
      {stage0_25[510]},
      {stage1_25[272]}
   );
   gpc1_1 gpc2066 (
      {stage0_25[511]},
      {stage1_25[273]}
   );
   gpc1_1 gpc2067 (
      {stage0_26[498]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2068 (
      {stage0_26[499]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2069 (
      {stage0_26[500]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2070 (
      {stage0_26[501]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2071 (
      {stage0_26[502]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2072 (
      {stage0_26[503]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2073 (
      {stage0_26[504]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2074 (
      {stage0_26[505]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2075 (
      {stage0_26[506]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2076 (
      {stage0_26[507]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2077 (
      {stage0_26[508]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2078 (
      {stage0_26[509]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2079 (
      {stage0_26[510]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2080 (
      {stage0_26[511]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2081 (
      {stage0_27[479]},
      {stage1_27[167]}
   );
   gpc1_1 gpc2082 (
      {stage0_27[480]},
      {stage1_27[168]}
   );
   gpc1_1 gpc2083 (
      {stage0_27[481]},
      {stage1_27[169]}
   );
   gpc1_1 gpc2084 (
      {stage0_27[482]},
      {stage1_27[170]}
   );
   gpc1_1 gpc2085 (
      {stage0_27[483]},
      {stage1_27[171]}
   );
   gpc1_1 gpc2086 (
      {stage0_27[484]},
      {stage1_27[172]}
   );
   gpc1_1 gpc2087 (
      {stage0_27[485]},
      {stage1_27[173]}
   );
   gpc1_1 gpc2088 (
      {stage0_27[486]},
      {stage1_27[174]}
   );
   gpc1_1 gpc2089 (
      {stage0_27[487]},
      {stage1_27[175]}
   );
   gpc1_1 gpc2090 (
      {stage0_27[488]},
      {stage1_27[176]}
   );
   gpc1_1 gpc2091 (
      {stage0_27[489]},
      {stage1_27[177]}
   );
   gpc1_1 gpc2092 (
      {stage0_27[490]},
      {stage1_27[178]}
   );
   gpc1_1 gpc2093 (
      {stage0_27[491]},
      {stage1_27[179]}
   );
   gpc1_1 gpc2094 (
      {stage0_27[492]},
      {stage1_27[180]}
   );
   gpc1_1 gpc2095 (
      {stage0_27[493]},
      {stage1_27[181]}
   );
   gpc1_1 gpc2096 (
      {stage0_27[494]},
      {stage1_27[182]}
   );
   gpc1_1 gpc2097 (
      {stage0_27[495]},
      {stage1_27[183]}
   );
   gpc1_1 gpc2098 (
      {stage0_27[496]},
      {stage1_27[184]}
   );
   gpc1_1 gpc2099 (
      {stage0_27[497]},
      {stage1_27[185]}
   );
   gpc1_1 gpc2100 (
      {stage0_27[498]},
      {stage1_27[186]}
   );
   gpc1_1 gpc2101 (
      {stage0_27[499]},
      {stage1_27[187]}
   );
   gpc1_1 gpc2102 (
      {stage0_27[500]},
      {stage1_27[188]}
   );
   gpc1_1 gpc2103 (
      {stage0_27[501]},
      {stage1_27[189]}
   );
   gpc1_1 gpc2104 (
      {stage0_27[502]},
      {stage1_27[190]}
   );
   gpc1_1 gpc2105 (
      {stage0_27[503]},
      {stage1_27[191]}
   );
   gpc1_1 gpc2106 (
      {stage0_27[504]},
      {stage1_27[192]}
   );
   gpc1_1 gpc2107 (
      {stage0_27[505]},
      {stage1_27[193]}
   );
   gpc1_1 gpc2108 (
      {stage0_27[506]},
      {stage1_27[194]}
   );
   gpc1_1 gpc2109 (
      {stage0_27[507]},
      {stage1_27[195]}
   );
   gpc1_1 gpc2110 (
      {stage0_27[508]},
      {stage1_27[196]}
   );
   gpc1_1 gpc2111 (
      {stage0_27[509]},
      {stage1_27[197]}
   );
   gpc1_1 gpc2112 (
      {stage0_27[510]},
      {stage1_27[198]}
   );
   gpc1_1 gpc2113 (
      {stage0_27[511]},
      {stage1_27[199]}
   );
   gpc1_1 gpc2114 (
      {stage0_28[506]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2115 (
      {stage0_28[507]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2116 (
      {stage0_28[508]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2117 (
      {stage0_28[509]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2118 (
      {stage0_28[510]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2119 (
      {stage0_28[511]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2120 (
      {stage0_29[509]},
      {stage1_29[240]}
   );
   gpc1_1 gpc2121 (
      {stage0_29[510]},
      {stage1_29[241]}
   );
   gpc1_1 gpc2122 (
      {stage0_29[511]},
      {stage1_29[242]}
   );
   gpc1_1 gpc2123 (
      {stage0_30[474]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2124 (
      {stage0_30[475]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2125 (
      {stage0_30[476]},
      {stage1_30[171]}
   );
   gpc1_1 gpc2126 (
      {stage0_30[477]},
      {stage1_30[172]}
   );
   gpc1_1 gpc2127 (
      {stage0_30[478]},
      {stage1_30[173]}
   );
   gpc1_1 gpc2128 (
      {stage0_30[479]},
      {stage1_30[174]}
   );
   gpc1_1 gpc2129 (
      {stage0_30[480]},
      {stage1_30[175]}
   );
   gpc1_1 gpc2130 (
      {stage0_30[481]},
      {stage1_30[176]}
   );
   gpc1_1 gpc2131 (
      {stage0_30[482]},
      {stage1_30[177]}
   );
   gpc1_1 gpc2132 (
      {stage0_30[483]},
      {stage1_30[178]}
   );
   gpc1_1 gpc2133 (
      {stage0_30[484]},
      {stage1_30[179]}
   );
   gpc1_1 gpc2134 (
      {stage0_30[485]},
      {stage1_30[180]}
   );
   gpc1_1 gpc2135 (
      {stage0_30[486]},
      {stage1_30[181]}
   );
   gpc1_1 gpc2136 (
      {stage0_30[487]},
      {stage1_30[182]}
   );
   gpc1_1 gpc2137 (
      {stage0_30[488]},
      {stage1_30[183]}
   );
   gpc1_1 gpc2138 (
      {stage0_30[489]},
      {stage1_30[184]}
   );
   gpc1_1 gpc2139 (
      {stage0_30[490]},
      {stage1_30[185]}
   );
   gpc1_1 gpc2140 (
      {stage0_30[491]},
      {stage1_30[186]}
   );
   gpc1_1 gpc2141 (
      {stage0_30[492]},
      {stage1_30[187]}
   );
   gpc1_1 gpc2142 (
      {stage0_30[493]},
      {stage1_30[188]}
   );
   gpc1_1 gpc2143 (
      {stage0_30[494]},
      {stage1_30[189]}
   );
   gpc1_1 gpc2144 (
      {stage0_30[495]},
      {stage1_30[190]}
   );
   gpc1_1 gpc2145 (
      {stage0_30[496]},
      {stage1_30[191]}
   );
   gpc1_1 gpc2146 (
      {stage0_30[497]},
      {stage1_30[192]}
   );
   gpc1_1 gpc2147 (
      {stage0_30[498]},
      {stage1_30[193]}
   );
   gpc1_1 gpc2148 (
      {stage0_30[499]},
      {stage1_30[194]}
   );
   gpc1_1 gpc2149 (
      {stage0_30[500]},
      {stage1_30[195]}
   );
   gpc1_1 gpc2150 (
      {stage0_30[501]},
      {stage1_30[196]}
   );
   gpc1_1 gpc2151 (
      {stage0_30[502]},
      {stage1_30[197]}
   );
   gpc1_1 gpc2152 (
      {stage0_30[503]},
      {stage1_30[198]}
   );
   gpc1_1 gpc2153 (
      {stage0_30[504]},
      {stage1_30[199]}
   );
   gpc1_1 gpc2154 (
      {stage0_30[505]},
      {stage1_30[200]}
   );
   gpc1_1 gpc2155 (
      {stage0_30[506]},
      {stage1_30[201]}
   );
   gpc1_1 gpc2156 (
      {stage0_30[507]},
      {stage1_30[202]}
   );
   gpc1_1 gpc2157 (
      {stage0_30[508]},
      {stage1_30[203]}
   );
   gpc1_1 gpc2158 (
      {stage0_30[509]},
      {stage1_30[204]}
   );
   gpc1_1 gpc2159 (
      {stage0_30[510]},
      {stage1_30[205]}
   );
   gpc1_1 gpc2160 (
      {stage0_30[511]},
      {stage1_30[206]}
   );
   gpc1_1 gpc2161 (
      {stage0_31[426]},
      {stage1_31[157]}
   );
   gpc1_1 gpc2162 (
      {stage0_31[427]},
      {stage1_31[158]}
   );
   gpc1_1 gpc2163 (
      {stage0_31[428]},
      {stage1_31[159]}
   );
   gpc1_1 gpc2164 (
      {stage0_31[429]},
      {stage1_31[160]}
   );
   gpc1_1 gpc2165 (
      {stage0_31[430]},
      {stage1_31[161]}
   );
   gpc1_1 gpc2166 (
      {stage0_31[431]},
      {stage1_31[162]}
   );
   gpc1_1 gpc2167 (
      {stage0_31[432]},
      {stage1_31[163]}
   );
   gpc1_1 gpc2168 (
      {stage0_31[433]},
      {stage1_31[164]}
   );
   gpc1_1 gpc2169 (
      {stage0_31[434]},
      {stage1_31[165]}
   );
   gpc1_1 gpc2170 (
      {stage0_31[435]},
      {stage1_31[166]}
   );
   gpc1_1 gpc2171 (
      {stage0_31[436]},
      {stage1_31[167]}
   );
   gpc1_1 gpc2172 (
      {stage0_31[437]},
      {stage1_31[168]}
   );
   gpc1_1 gpc2173 (
      {stage0_31[438]},
      {stage1_31[169]}
   );
   gpc1_1 gpc2174 (
      {stage0_31[439]},
      {stage1_31[170]}
   );
   gpc1_1 gpc2175 (
      {stage0_31[440]},
      {stage1_31[171]}
   );
   gpc1_1 gpc2176 (
      {stage0_31[441]},
      {stage1_31[172]}
   );
   gpc1_1 gpc2177 (
      {stage0_31[442]},
      {stage1_31[173]}
   );
   gpc1_1 gpc2178 (
      {stage0_31[443]},
      {stage1_31[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_31[444]},
      {stage1_31[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_31[445]},
      {stage1_31[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_31[446]},
      {stage1_31[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_31[447]},
      {stage1_31[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_31[448]},
      {stage1_31[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_31[449]},
      {stage1_31[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_31[450]},
      {stage1_31[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_31[451]},
      {stage1_31[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_31[452]},
      {stage1_31[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_31[453]},
      {stage1_31[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_31[454]},
      {stage1_31[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_31[455]},
      {stage1_31[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_31[456]},
      {stage1_31[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_31[457]},
      {stage1_31[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_31[458]},
      {stage1_31[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_31[459]},
      {stage1_31[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_31[460]},
      {stage1_31[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_31[461]},
      {stage1_31[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_31[462]},
      {stage1_31[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_31[463]},
      {stage1_31[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_31[464]},
      {stage1_31[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_31[465]},
      {stage1_31[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_31[466]},
      {stage1_31[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_31[467]},
      {stage1_31[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_31[468]},
      {stage1_31[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_31[469]},
      {stage1_31[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_31[470]},
      {stage1_31[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_31[471]},
      {stage1_31[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_31[472]},
      {stage1_31[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_31[473]},
      {stage1_31[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_31[474]},
      {stage1_31[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_31[475]},
      {stage1_31[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_31[476]},
      {stage1_31[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_31[477]},
      {stage1_31[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_31[478]},
      {stage1_31[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_31[479]},
      {stage1_31[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_31[480]},
      {stage1_31[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_31[481]},
      {stage1_31[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_31[482]},
      {stage1_31[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_31[483]},
      {stage1_31[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_31[484]},
      {stage1_31[215]}
   );
   gpc1_1 gpc2220 (
      {stage0_31[485]},
      {stage1_31[216]}
   );
   gpc1_1 gpc2221 (
      {stage0_31[486]},
      {stage1_31[217]}
   );
   gpc1_1 gpc2222 (
      {stage0_31[487]},
      {stage1_31[218]}
   );
   gpc1_1 gpc2223 (
      {stage0_31[488]},
      {stage1_31[219]}
   );
   gpc1_1 gpc2224 (
      {stage0_31[489]},
      {stage1_31[220]}
   );
   gpc1_1 gpc2225 (
      {stage0_31[490]},
      {stage1_31[221]}
   );
   gpc1_1 gpc2226 (
      {stage0_31[491]},
      {stage1_31[222]}
   );
   gpc1_1 gpc2227 (
      {stage0_31[492]},
      {stage1_31[223]}
   );
   gpc1_1 gpc2228 (
      {stage0_31[493]},
      {stage1_31[224]}
   );
   gpc1_1 gpc2229 (
      {stage0_31[494]},
      {stage1_31[225]}
   );
   gpc1_1 gpc2230 (
      {stage0_31[495]},
      {stage1_31[226]}
   );
   gpc1_1 gpc2231 (
      {stage0_31[496]},
      {stage1_31[227]}
   );
   gpc1_1 gpc2232 (
      {stage0_31[497]},
      {stage1_31[228]}
   );
   gpc1_1 gpc2233 (
      {stage0_31[498]},
      {stage1_31[229]}
   );
   gpc1_1 gpc2234 (
      {stage0_31[499]},
      {stage1_31[230]}
   );
   gpc1_1 gpc2235 (
      {stage0_31[500]},
      {stage1_31[231]}
   );
   gpc1_1 gpc2236 (
      {stage0_31[501]},
      {stage1_31[232]}
   );
   gpc1_1 gpc2237 (
      {stage0_31[502]},
      {stage1_31[233]}
   );
   gpc1_1 gpc2238 (
      {stage0_31[503]},
      {stage1_31[234]}
   );
   gpc1_1 gpc2239 (
      {stage0_31[504]},
      {stage1_31[235]}
   );
   gpc1_1 gpc2240 (
      {stage0_31[505]},
      {stage1_31[236]}
   );
   gpc1_1 gpc2241 (
      {stage0_31[506]},
      {stage1_31[237]}
   );
   gpc1_1 gpc2242 (
      {stage0_31[507]},
      {stage1_31[238]}
   );
   gpc1_1 gpc2243 (
      {stage0_31[508]},
      {stage1_31[239]}
   );
   gpc1_1 gpc2244 (
      {stage0_31[509]},
      {stage1_31[240]}
   );
   gpc1_1 gpc2245 (
      {stage0_31[510]},
      {stage1_31[241]}
   );
   gpc1_1 gpc2246 (
      {stage0_31[511]},
      {stage1_31[242]}
   );
   gpc2135_5 gpc2247 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc2248 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc2249 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc2250 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc2251 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[12]},
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2252 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2253 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[14]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc2254 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[15]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc2255 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[16]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc2256 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[17]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc2257 (
      {stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54]},
      {stage1_1[18]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc2258 (
      {stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[19]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2259 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[0],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc2260 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage2_5[1],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc2261 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25]},
      {stage2_5[2],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc2262 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage2_5[3],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc2263 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage2_5[4],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc2264 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage2_5[5],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc2265 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage2_5[6],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc2266 (
      {stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65], stage1_1[66], stage1_1[67]},
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage2_5[7],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc606_5 gpc2267 (
      {stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71], stage1_1[72], stage1_1[73]},
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage2_5[8],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc606_5 gpc2268 (
      {stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78], stage1_1[79]},
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage2_5[9],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc2269 (
      {stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84], stage1_1[85]},
      {stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage2_5[10],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2270 (
      {stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90], stage1_1[91]},
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79]},
      {stage2_5[11],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2271 (
      {stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96], stage1_1[97]},
      {stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage2_5[12],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2272 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage2_5[13],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2273 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage2_5[14],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2274 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage2_5[15],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2275 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109]},
      {stage2_5[16],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2276 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage2_5[17],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2277 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121]},
      {stage2_5[18],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2278 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage2_5[19],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc2279 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage2_5[20],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc2280 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139]},
      {stage2_5[21],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc2281 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage2_5[22],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc2282 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150], stage1_3[151]},
      {stage2_5[23],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc2283 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], stage1_1[169]},
      {stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157]},
      {stage2_5[24],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc2284 (
      {stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174], stage1_1[175]},
      {stage1_3[158], stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage2_5[25],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc2285 (
      {stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], stage1_1[180], stage1_1[181]},
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169]},
      {stage2_5[26],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc615_5 gpc2286 (
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56]},
      {stage1_3[170]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[27],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc2287 (
      {stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_3[171]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[28],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc2288 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage1_3[172]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[29],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc2289 (
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_3[173]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[30],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc2290 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76]},
      {stage1_3[174]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[31],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2291 (
      {stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage1_3[175]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[32],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2292 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86]},
      {stage1_3[176]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[33],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2293 (
      {stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91]},
      {stage1_3[177]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[34],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2294 (
      {stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage1_3[178]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[35],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc2295 (
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage1_3[179]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[36],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc2296 (
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106]},
      {stage1_3[180]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[37],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc2297 (
      {stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_3[181]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[38],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc2298 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116]},
      {stage1_3[182]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[39],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc2299 (
      {stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121]},
      {stage1_3[183]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[40],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc2300 (
      {stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage1_3[184]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[41],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc2301 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_3[185]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[42],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc2302 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136]},
      {stage1_3[186]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[43],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc2303 (
      {stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_3[187]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[44],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc2304 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146]},
      {stage1_3[188]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[45],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc2305 (
      {stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151]},
      {stage1_3[189]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[46],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc2306 (
      {stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194]},
      {stage1_4[120]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[20],stage2_5[47],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2307 (
      {stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199]},
      {stage1_4[121]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[21],stage2_5[48],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2308 (
      {stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204]},
      {stage1_4[122]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[22],stage2_5[49],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2309 (
      {stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209]},
      {stage1_4[123]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[23],stage2_5[50],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2310 (
      {stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214]},
      {stage1_4[124]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[24],stage2_5[51],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2311 (
      {stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219]},
      {stage1_4[125]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[25],stage2_5[52],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2312 (
      {stage1_3[220], stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224]},
      {stage1_4[126]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[26],stage2_5[53],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2313 (
      {stage1_3[225], stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229]},
      {stage1_4[127]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[27],stage2_5[54],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2314 (
      {stage1_3[230], stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234]},
      {stage1_4[128]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[28],stage2_5[55],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2315 (
      {stage1_3[235], stage1_3[236], stage1_3[237], stage1_3[238], stage1_3[239]},
      {stage1_4[129]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[29],stage2_5[56],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc2316 (
      {stage1_3[240], stage1_3[241], stage1_3[242], stage1_3[243], stage1_3[244]},
      {stage1_4[130]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[30],stage2_5[57],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[245], stage1_3[246], stage1_3[247], stage1_3[248], stage1_3[249]},
      {stage1_4[131]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[31],stage2_5[58],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[250], stage1_3[251], stage1_3[252], stage1_3[253], stage1_3[254]},
      {stage1_4[132]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[32],stage2_5[59],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[255], stage1_3[256], stage1_3[257], stage1_3[258], stage1_3[259]},
      {stage1_4[133]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[33],stage2_5[60],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[260], stage1_3[261], stage1_3[262], stage1_3[263], stage1_3[264]},
      {stage1_4[134]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[34],stage2_5[61],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[265], stage1_3[266], stage1_3[267], stage1_3[268], stage1_3[269]},
      {stage1_4[135]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[35],stage2_5[62],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[270], stage1_3[271], stage1_3[272], stage1_3[273], stage1_3[274]},
      {stage1_4[136]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[36],stage2_5[63],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[275], stage1_3[276], 1'b0, 1'b0, 1'b0},
      {stage1_4[137]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[37],stage2_5[64],stage2_4[76],stage2_3[76]}
   );
   gpc1163_5 gpc2324 (
      {stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[18],stage2_6[38],stage2_5[65],stage2_4[77]}
   );
   gpc606_5 gpc2325 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[19],stage2_6[39],stage2_5[66],stage2_4[78]}
   );
   gpc606_5 gpc2326 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[20],stage2_6[40],stage2_5[67],stage2_4[79]}
   );
   gpc606_5 gpc2327 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[21],stage2_6[41],stage2_5[68],stage2_4[80]}
   );
   gpc606_5 gpc2328 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[22],stage2_6[42],stage2_5[69],stage2_4[81]}
   );
   gpc606_5 gpc2329 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[23],stage2_6[43],stage2_5[70],stage2_4[82]}
   );
   gpc606_5 gpc2330 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[24],stage2_6[44],stage2_5[71],stage2_4[83]}
   );
   gpc606_5 gpc2331 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[25],stage2_6[45],stage2_5[72],stage2_4[84]}
   );
   gpc606_5 gpc2332 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[26],stage2_6[46],stage2_5[73],stage2_4[85]}
   );
   gpc606_5 gpc2333 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[27],stage2_6[47],stage2_5[74],stage2_4[86]}
   );
   gpc606_5 gpc2334 (
      {stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[28],stage2_6[48],stage2_5[75],stage2_4[87]}
   );
   gpc606_5 gpc2335 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[29],stage2_6[49],stage2_5[76],stage2_4[88]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[114]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[30],stage2_6[50],stage2_5[77],stage2_4[89]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[115]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[31],stage2_6[51],stage2_5[78],stage2_4[90]}
   );
   gpc606_5 gpc2338 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[14],stage2_7[32],stage2_6[52],stage2_5[79]}
   );
   gpc606_5 gpc2339 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[15],stage2_7[33],stage2_6[53],stage2_5[80]}
   );
   gpc606_5 gpc2340 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[16],stage2_7[34],stage2_6[54],stage2_5[81]}
   );
   gpc606_5 gpc2341 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[17],stage2_7[35],stage2_6[55],stage2_5[82]}
   );
   gpc606_5 gpc2342 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[18],stage2_7[36],stage2_6[56],stage2_5[83]}
   );
   gpc606_5 gpc2343 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[19],stage2_7[37],stage2_6[57],stage2_5[84]}
   );
   gpc606_5 gpc2344 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[20],stage2_7[38],stage2_6[58],stage2_5[85]}
   );
   gpc606_5 gpc2345 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[21],stage2_7[39],stage2_6[59],stage2_5[86]}
   );
   gpc606_5 gpc2346 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[22],stage2_7[40],stage2_6[60],stage2_5[87]}
   );
   gpc606_5 gpc2347 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[23],stage2_7[41],stage2_6[61],stage2_5[88]}
   );
   gpc606_5 gpc2348 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage2_9[10],stage2_8[24],stage2_7[42],stage2_6[62],stage2_5[89]}
   );
   gpc606_5 gpc2349 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72]},
      {stage2_9[11],stage2_8[25],stage2_7[43],stage2_6[63],stage2_5[90]}
   );
   gpc606_5 gpc2350 (
      {stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193]},
      {stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78]},
      {stage2_9[12],stage2_8[26],stage2_7[44],stage2_6[64],stage2_5[91]}
   );
   gpc606_5 gpc2351 (
      {stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199]},
      {stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84]},
      {stage2_9[13],stage2_8[27],stage2_7[45],stage2_6[65],stage2_5[92]}
   );
   gpc606_5 gpc2352 (
      {stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205]},
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90]},
      {stage2_9[14],stage2_8[28],stage2_7[46],stage2_6[66],stage2_5[93]}
   );
   gpc606_5 gpc2353 (
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[29],stage2_7[47],stage2_6[67]}
   );
   gpc606_5 gpc2354 (
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[30],stage2_7[48],stage2_6[68]}
   );
   gpc606_5 gpc2355 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[31],stage2_7[49],stage2_6[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[32],stage2_7[50],stage2_6[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[33],stage2_7[51],stage2_6[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[20],stage2_8[34],stage2_7[52],stage2_6[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[21],stage2_8[35],stage2_7[53],stage2_6[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[22],stage2_8[36],stage2_7[54],stage2_6[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[23],stage2_8[37],stage2_7[55],stage2_6[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[24],stage2_8[38],stage2_7[56],stage2_6[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[25],stage2_8[39],stage2_7[57],stage2_6[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[26],stage2_8[40],stage2_7[58],stage2_6[78]}
   );
   gpc606_5 gpc2365 (
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[27],stage2_8[41],stage2_7[59],stage2_6[79]}
   );
   gpc606_5 gpc2366 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[28],stage2_8[42],stage2_7[60],stage2_6[80]}
   );
   gpc606_5 gpc2367 (
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[29],stage2_8[43],stage2_7[61],stage2_6[81]}
   );
   gpc606_5 gpc2368 (
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[30],stage2_8[44],stage2_7[62],stage2_6[82]}
   );
   gpc606_5 gpc2369 (
      {stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[31],stage2_8[45],stage2_7[63],stage2_6[83]}
   );
   gpc606_5 gpc2370 (
      {stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[32],stage2_8[46],stage2_7[64],stage2_6[84]}
   );
   gpc606_5 gpc2371 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191], stage1_6[192]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[33],stage2_8[47],stage2_7[65],stage2_6[85]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196], stage1_6[197]},
      {stage1_7[91]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[34],stage2_8[48],stage2_7[66],stage2_6[86]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201], stage1_6[202]},
      {stage1_7[92]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[35],stage2_8[49],stage2_7[67],stage2_6[87]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206], stage1_6[207]},
      {stage1_7[93]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[36],stage2_8[50],stage2_7[68],stage2_6[88]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211], stage1_6[212]},
      {stage1_7[94]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[37],stage2_8[51],stage2_7[69],stage2_6[89]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216], stage1_6[217]},
      {stage1_7[95]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[38],stage2_8[52],stage2_7[70],stage2_6[90]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221], stage1_6[222]},
      {stage1_7[96]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[39],stage2_8[53],stage2_7[71],stage2_6[91]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226], stage1_6[227]},
      {stage1_7[97]},
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage2_10[25],stage2_9[40],stage2_8[54],stage2_7[72],stage2_6[92]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231], stage1_6[232]},
      {stage1_7[98]},
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage2_10[26],stage2_9[41],stage2_8[55],stage2_7[73],stage2_6[93]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236], stage1_6[237]},
      {stage1_7[99]},
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage2_10[27],stage2_9[42],stage2_8[56],stage2_7[74],stage2_6[94]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241], stage1_6[242]},
      {stage1_7[100]},
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage2_10[28],stage2_9[43],stage2_8[57],stage2_7[75],stage2_6[95]}
   );
   gpc615_5 gpc2382 (
      {stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105]},
      {stage1_8[174]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[29],stage2_9[44],stage2_8[58],stage2_7[76]}
   );
   gpc615_5 gpc2383 (
      {stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110]},
      {stage1_8[175]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[30],stage2_9[45],stage2_8[59],stage2_7[77]}
   );
   gpc615_5 gpc2384 (
      {stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage1_8[176]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[31],stage2_9[46],stage2_8[60],stage2_7[78]}
   );
   gpc615_5 gpc2385 (
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_8[177]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[32],stage2_9[47],stage2_8[61],stage2_7[79]}
   );
   gpc615_5 gpc2386 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage1_8[178]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[33],stage2_9[48],stage2_8[62],stage2_7[80]}
   );
   gpc615_5 gpc2387 (
      {stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130]},
      {stage1_8[179]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[34],stage2_9[49],stage2_8[63],stage2_7[81]}
   );
   gpc615_5 gpc2388 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[180]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[35],stage2_9[50],stage2_8[64],stage2_7[82]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[181]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[36],stage2_9[51],stage2_8[65],stage2_7[83]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[182]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[37],stage2_9[52],stage2_8[66],stage2_7[84]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[183]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[38],stage2_9[53],stage2_8[67],stage2_7[85]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[184]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[39],stage2_9[54],stage2_8[68],stage2_7[86]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[185]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[40],stage2_9[55],stage2_8[69],stage2_7[87]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[186]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[41],stage2_9[56],stage2_8[70],stage2_7[88]}
   );
   gpc606_5 gpc2395 (
      {stage1_8[187], stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[13],stage2_10[42],stage2_9[57],stage2_8[71]}
   );
   gpc606_5 gpc2396 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197], stage1_8[198]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[14],stage2_10[43],stage2_9[58],stage2_8[72]}
   );
   gpc606_5 gpc2397 (
      {stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202], stage1_8[203], stage1_8[204]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[15],stage2_10[44],stage2_9[59],stage2_8[73]}
   );
   gpc606_5 gpc2398 (
      {stage1_8[205], stage1_8[206], stage1_8[207], stage1_8[208], stage1_8[209], stage1_8[210]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[16],stage2_10[45],stage2_9[60],stage2_8[74]}
   );
   gpc606_5 gpc2399 (
      {stage1_8[211], stage1_8[212], stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[17],stage2_10[46],stage2_9[61],stage2_8[75]}
   );
   gpc606_5 gpc2400 (
      {stage1_8[217], stage1_8[218], stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[18],stage2_10[47],stage2_9[62],stage2_8[76]}
   );
   gpc606_5 gpc2401 (
      {stage1_8[223], stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[19],stage2_10[48],stage2_9[63],stage2_8[77]}
   );
   gpc606_5 gpc2402 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233], stage1_8[234]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[20],stage2_10[49],stage2_9[64],stage2_8[78]}
   );
   gpc606_5 gpc2403 (
      {stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238], stage1_8[239], stage1_8[240]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[21],stage2_10[50],stage2_9[65],stage2_8[79]}
   );
   gpc606_5 gpc2404 (
      {stage1_8[241], stage1_8[242], stage1_8[243], stage1_8[244], stage1_8[245], stage1_8[246]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[22],stage2_10[51],stage2_9[66],stage2_8[80]}
   );
   gpc606_5 gpc2405 (
      {stage1_8[247], stage1_8[248], stage1_8[249], stage1_8[250], stage1_8[251], stage1_8[252]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[23],stage2_10[52],stage2_9[67],stage2_8[81]}
   );
   gpc606_5 gpc2406 (
      {stage1_8[253], stage1_8[254], stage1_8[255], stage1_8[256], stage1_8[257], stage1_8[258]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[24],stage2_10[53],stage2_9[68],stage2_8[82]}
   );
   gpc606_5 gpc2407 (
      {stage1_8[259], stage1_8[260], stage1_8[261], stage1_8[262], stage1_8[263], stage1_8[264]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[25],stage2_10[54],stage2_9[69],stage2_8[83]}
   );
   gpc606_5 gpc2408 (
      {stage1_8[265], stage1_8[266], stage1_8[267], stage1_8[268], stage1_8[269], stage1_8[270]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[26],stage2_10[55],stage2_9[70],stage2_8[84]}
   );
   gpc606_5 gpc2409 (
      {stage1_8[271], stage1_8[272], stage1_8[273], stage1_8[274], stage1_8[275], stage1_8[276]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[27],stage2_10[56],stage2_9[71],stage2_8[85]}
   );
   gpc606_5 gpc2410 (
      {stage1_8[277], stage1_8[278], stage1_8[279], stage1_8[280], stage1_8[281], stage1_8[282]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[28],stage2_10[57],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc2411 (
      {stage1_8[283], stage1_8[284], stage1_8[285], stage1_8[286], stage1_8[287], stage1_8[288]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[29],stage2_10[58],stage2_9[73],stage2_8[87]}
   );
   gpc606_5 gpc2412 (
      {stage1_8[289], stage1_8[290], stage1_8[291], stage1_8[292], stage1_8[293], stage1_8[294]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[30],stage2_10[59],stage2_9[74],stage2_8[88]}
   );
   gpc606_5 gpc2413 (
      {stage1_8[295], stage1_8[296], stage1_8[297], stage1_8[298], stage1_8[299], stage1_8[300]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[31],stage2_10[60],stage2_9[75],stage2_8[89]}
   );
   gpc606_5 gpc2414 (
      {stage1_8[301], stage1_8[302], stage1_8[303], stage1_8[304], stage1_8[305], stage1_8[306]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[32],stage2_10[61],stage2_9[76],stage2_8[90]}
   );
   gpc606_5 gpc2415 (
      {stage1_8[307], stage1_8[308], stage1_8[309], stage1_8[310], stage1_8[311], stage1_8[312]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[33],stage2_10[62],stage2_9[77],stage2_8[91]}
   );
   gpc606_5 gpc2416 (
      {stage1_8[313], stage1_8[314], stage1_8[315], stage1_8[316], stage1_8[317], stage1_8[318]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[34],stage2_10[63],stage2_9[78],stage2_8[92]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[319], stage1_8[320], stage1_8[321], stage1_8[322], stage1_8[323], stage1_8[324]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[35],stage2_10[64],stage2_9[79],stage2_8[93]}
   );
   gpc606_5 gpc2418 (
      {stage1_8[325], stage1_8[326], stage1_8[327], stage1_8[328], stage1_8[329], stage1_8[330]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[36],stage2_10[65],stage2_9[80],stage2_8[94]}
   );
   gpc606_5 gpc2419 (
      {stage1_8[331], stage1_8[332], stage1_8[333], stage1_8[334], stage1_8[335], stage1_8[336]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[37],stage2_10[66],stage2_9[81],stage2_8[95]}
   );
   gpc606_5 gpc2420 (
      {stage1_8[337], stage1_8[338], stage1_8[339], stage1_8[340], stage1_8[341], stage1_8[342]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[38],stage2_10[67],stage2_9[82],stage2_8[96]}
   );
   gpc606_5 gpc2421 (
      {stage1_8[343], stage1_8[344], stage1_8[345], stage1_8[346], stage1_8[347], stage1_8[348]},
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage2_12[26],stage2_11[39],stage2_10[68],stage2_9[83],stage2_8[97]}
   );
   gpc606_5 gpc2422 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[27],stage2_11[40],stage2_10[69],stage2_9[84]}
   );
   gpc606_5 gpc2423 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[28],stage2_11[41],stage2_10[70],stage2_9[85]}
   );
   gpc606_5 gpc2424 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[29],stage2_11[42],stage2_10[71],stage2_9[86]}
   );
   gpc606_5 gpc2425 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[30],stage2_11[43],stage2_10[72],stage2_9[87]}
   );
   gpc606_5 gpc2426 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[31],stage2_11[44],stage2_10[73],stage2_9[88]}
   );
   gpc606_5 gpc2427 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[32],stage2_11[45],stage2_10[74],stage2_9[89]}
   );
   gpc606_5 gpc2428 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[33],stage2_11[46],stage2_10[75],stage2_9[90]}
   );
   gpc606_5 gpc2429 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[34],stage2_11[47],stage2_10[76],stage2_9[91]}
   );
   gpc606_5 gpc2430 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[35],stage2_11[48],stage2_10[77],stage2_9[92]}
   );
   gpc606_5 gpc2431 (
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[36],stage2_11[49],stage2_10[78],stage2_9[93]}
   );
   gpc606_5 gpc2432 (
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[37],stage2_11[50],stage2_10[79],stage2_9[94]}
   );
   gpc606_5 gpc2433 (
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[38],stage2_11[51],stage2_10[80],stage2_9[95]}
   );
   gpc606_5 gpc2434 (
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[39],stage2_11[52],stage2_10[81],stage2_9[96]}
   );
   gpc606_5 gpc2435 (
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[40],stage2_11[53],stage2_10[82],stage2_9[97]}
   );
   gpc606_5 gpc2436 (
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[41],stage2_11[54],stage2_10[83],stage2_9[98]}
   );
   gpc606_5 gpc2437 (
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[42],stage2_11[55],stage2_10[84],stage2_9[99]}
   );
   gpc606_5 gpc2438 (
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[43],stage2_11[56],stage2_10[85],stage2_9[100]}
   );
   gpc606_5 gpc2439 (
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[44],stage2_11[57],stage2_10[86],stage2_9[101]}
   );
   gpc606_5 gpc2440 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage2_13[18],stage2_12[45],stage2_11[58],stage2_10[87],stage2_9[102]}
   );
   gpc606_5 gpc2441 (
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage2_13[19],stage2_12[46],stage2_11[59],stage2_10[88],stage2_9[103]}
   );
   gpc606_5 gpc2442 (
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125]},
      {stage2_13[20],stage2_12[47],stage2_11[60],stage2_10[89],stage2_9[104]}
   );
   gpc606_5 gpc2443 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131]},
      {stage2_13[21],stage2_12[48],stage2_11[61],stage2_10[90],stage2_9[105]}
   );
   gpc615_5 gpc2444 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_11[132]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[22],stage2_12[49],stage2_11[62],stage2_10[91]}
   );
   gpc615_5 gpc2445 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171]},
      {stage1_11[133]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[23],stage2_12[50],stage2_11[63],stage2_10[92]}
   );
   gpc615_5 gpc2446 (
      {stage1_10[172], stage1_10[173], stage1_10[174], stage1_10[175], stage1_10[176]},
      {stage1_11[134]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[24],stage2_12[51],stage2_11[64],stage2_10[93]}
   );
   gpc615_5 gpc2447 (
      {stage1_10[177], stage1_10[178], stage1_10[179], stage1_10[180], stage1_10[181]},
      {stage1_11[135]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[25],stage2_12[52],stage2_11[65],stage2_10[94]}
   );
   gpc615_5 gpc2448 (
      {stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139], stage1_11[140]},
      {stage1_12[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[4],stage2_13[26],stage2_12[53],stage2_11[66]}
   );
   gpc615_5 gpc2449 (
      {stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144], stage1_11[145]},
      {stage1_12[25]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[5],stage2_13[27],stage2_12[54],stage2_11[67]}
   );
   gpc615_5 gpc2450 (
      {stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[26]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[6],stage2_13[28],stage2_12[55],stage2_11[68]}
   );
   gpc615_5 gpc2451 (
      {stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154], stage1_11[155]},
      {stage1_12[27]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[7],stage2_13[29],stage2_12[56],stage2_11[69]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159], stage1_11[160]},
      {stage1_12[28]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[8],stage2_13[30],stage2_12[57],stage2_11[70]}
   );
   gpc606_5 gpc2453 (
      {stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[5],stage2_14[9],stage2_13[31],stage2_12[58]}
   );
   gpc615_5 gpc2454 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39]},
      {stage1_13[30]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[6],stage2_14[10],stage2_13[32],stage2_12[59]}
   );
   gpc615_5 gpc2455 (
      {stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_13[31]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[7],stage2_14[11],stage2_13[33],stage2_12[60]}
   );
   gpc615_5 gpc2456 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_13[32]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[8],stage2_14[12],stage2_13[34],stage2_12[61]}
   );
   gpc615_5 gpc2457 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54]},
      {stage1_13[33]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[9],stage2_14[13],stage2_13[35],stage2_12[62]}
   );
   gpc615_5 gpc2458 (
      {stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[34]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[10],stage2_14[14],stage2_13[36],stage2_12[63]}
   );
   gpc615_5 gpc2459 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64]},
      {stage1_13[35]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[11],stage2_14[15],stage2_13[37],stage2_12[64]}
   );
   gpc615_5 gpc2460 (
      {stage1_12[65], stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69]},
      {stage1_13[36]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[12],stage2_14[16],stage2_13[38],stage2_12[65]}
   );
   gpc615_5 gpc2461 (
      {stage1_12[70], stage1_12[71], stage1_12[72], stage1_12[73], stage1_12[74]},
      {stage1_13[37]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[13],stage2_14[17],stage2_13[39],stage2_12[66]}
   );
   gpc615_5 gpc2462 (
      {stage1_12[75], stage1_12[76], stage1_12[77], stage1_12[78], stage1_12[79]},
      {stage1_13[38]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[14],stage2_14[18],stage2_13[40],stage2_12[67]}
   );
   gpc615_5 gpc2463 (
      {stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_13[39]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[15],stage2_14[19],stage2_13[41],stage2_12[68]}
   );
   gpc615_5 gpc2464 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[40]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[16],stage2_14[20],stage2_13[42],stage2_12[69]}
   );
   gpc615_5 gpc2465 (
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94]},
      {stage1_13[41]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[17],stage2_14[21],stage2_13[43],stage2_12[70]}
   );
   gpc615_5 gpc2466 (
      {stage1_12[95], stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99]},
      {stage1_13[42]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[18],stage2_14[22],stage2_13[44],stage2_12[71]}
   );
   gpc615_5 gpc2467 (
      {stage1_12[100], stage1_12[101], stage1_12[102], stage1_12[103], stage1_12[104]},
      {stage1_13[43]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[19],stage2_14[23],stage2_13[45],stage2_12[72]}
   );
   gpc615_5 gpc2468 (
      {stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108], stage1_12[109]},
      {stage1_13[44]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[20],stage2_14[24],stage2_13[46],stage2_12[73]}
   );
   gpc615_5 gpc2469 (
      {stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_13[45]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[21],stage2_14[25],stage2_13[47],stage2_12[74]}
   );
   gpc615_5 gpc2470 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[46]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[22],stage2_14[26],stage2_13[48],stage2_12[75]}
   );
   gpc615_5 gpc2471 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_13[47]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[23],stage2_14[27],stage2_13[49],stage2_12[76]}
   );
   gpc615_5 gpc2472 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129]},
      {stage1_13[48]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[24],stage2_14[28],stage2_13[50],stage2_12[77]}
   );
   gpc615_5 gpc2473 (
      {stage1_12[130], stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134]},
      {stage1_13[49]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[25],stage2_14[29],stage2_13[51],stage2_12[78]}
   );
   gpc615_5 gpc2474 (
      {stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138], stage1_12[139]},
      {stage1_13[50]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[26],stage2_14[30],stage2_13[52],stage2_12[79]}
   );
   gpc615_5 gpc2475 (
      {stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_13[51]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[27],stage2_14[31],stage2_13[53],stage2_12[80]}
   );
   gpc615_5 gpc2476 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_13[52]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[28],stage2_14[32],stage2_13[54],stage2_12[81]}
   );
   gpc615_5 gpc2477 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_13[53]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[29],stage2_14[33],stage2_13[55],stage2_12[82]}
   );
   gpc615_5 gpc2478 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159]},
      {stage1_13[54]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[30],stage2_14[34],stage2_13[56],stage2_12[83]}
   );
   gpc615_5 gpc2479 (
      {stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_13[55]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[31],stage2_14[35],stage2_13[57],stage2_12[84]}
   );
   gpc615_5 gpc2480 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169]},
      {stage1_13[56]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[32],stage2_14[36],stage2_13[58],stage2_12[85]}
   );
   gpc615_5 gpc2481 (
      {stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_13[57]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[33],stage2_14[37],stage2_13[59],stage2_12[86]}
   );
   gpc615_5 gpc2482 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_13[58]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[34],stage2_14[38],stage2_13[60],stage2_12[87]}
   );
   gpc615_5 gpc2483 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184]},
      {stage1_13[59]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[35],stage2_14[39],stage2_13[61],stage2_12[88]}
   );
   gpc615_5 gpc2484 (
      {stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189]},
      {stage1_13[60]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[36],stage2_14[40],stage2_13[62],stage2_12[89]}
   );
   gpc615_5 gpc2485 (
      {stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_13[61]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[37],stage2_14[41],stage2_13[63],stage2_12[90]}
   );
   gpc615_5 gpc2486 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199]},
      {stage1_13[62]},
      {stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203]},
      {stage2_16[33],stage2_15[38],stage2_14[42],stage2_13[64],stage2_12[91]}
   );
   gpc615_5 gpc2487 (
      {stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_13[63]},
      {stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209]},
      {stage2_16[34],stage2_15[39],stage2_14[43],stage2_13[65],stage2_12[92]}
   );
   gpc615_5 gpc2488 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_13[64]},
      {stage1_14[210], stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage2_16[35],stage2_15[40],stage2_14[44],stage2_13[66],stage2_12[93]}
   );
   gpc615_5 gpc2489 (
      {stage1_12[210], stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214]},
      {stage1_13[65]},
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221]},
      {stage2_16[36],stage2_15[41],stage2_14[45],stage2_13[67],stage2_12[94]}
   );
   gpc606_5 gpc2490 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[37],stage2_15[42],stage2_14[46],stage2_13[68]}
   );
   gpc606_5 gpc2491 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[38],stage2_15[43],stage2_14[47],stage2_13[69]}
   );
   gpc606_5 gpc2492 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[39],stage2_15[44],stage2_14[48],stage2_13[70]}
   );
   gpc606_5 gpc2493 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[40],stage2_15[45],stage2_14[49],stage2_13[71]}
   );
   gpc606_5 gpc2494 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[41],stage2_15[46],stage2_14[50],stage2_13[72]}
   );
   gpc606_5 gpc2495 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[42],stage2_15[47],stage2_14[51],stage2_13[73]}
   );
   gpc606_5 gpc2496 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[43],stage2_15[48],stage2_14[52],stage2_13[74]}
   );
   gpc606_5 gpc2497 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[44],stage2_15[49],stage2_14[53],stage2_13[75]}
   );
   gpc606_5 gpc2498 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[45],stage2_15[50],stage2_14[54],stage2_13[76]}
   );
   gpc606_5 gpc2499 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[46],stage2_15[51],stage2_14[55],stage2_13[77]}
   );
   gpc606_5 gpc2500 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[47],stage2_15[52],stage2_14[56],stage2_13[78]}
   );
   gpc606_5 gpc2501 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[48],stage2_15[53],stage2_14[57],stage2_13[79]}
   );
   gpc606_5 gpc2502 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[49],stage2_15[54],stage2_14[58],stage2_13[80]}
   );
   gpc606_5 gpc2503 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[50],stage2_15[55],stage2_14[59],stage2_13[81]}
   );
   gpc606_5 gpc2504 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[51],stage2_15[56],stage2_14[60],stage2_13[82]}
   );
   gpc606_5 gpc2505 (
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[52],stage2_15[57],stage2_14[61],stage2_13[83]}
   );
   gpc606_5 gpc2506 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[53],stage2_15[58],stage2_14[62],stage2_13[84]}
   );
   gpc606_5 gpc2507 (
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[54],stage2_15[59],stage2_14[63],stage2_13[85]}
   );
   gpc606_5 gpc2508 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[55],stage2_15[60],stage2_14[64],stage2_13[86]}
   );
   gpc606_5 gpc2509 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[56],stage2_15[61],stage2_14[65],stage2_13[87]}
   );
   gpc606_5 gpc2510 (
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[57],stage2_15[62],stage2_14[66],stage2_13[88]}
   );
   gpc606_5 gpc2511 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[58],stage2_15[63],stage2_14[67],stage2_13[89]}
   );
   gpc615_5 gpc2512 (
      {stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226]},
      {stage1_15[132]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[22],stage2_16[59],stage2_15[64],stage2_14[68]}
   );
   gpc615_5 gpc2513 (
      {stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231]},
      {stage1_15[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[23],stage2_16[60],stage2_15[65],stage2_14[69]}
   );
   gpc606_5 gpc2514 (
      {stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137], stage1_15[138], stage1_15[139]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[24],stage2_16[61],stage2_15[66]}
   );
   gpc606_5 gpc2515 (
      {stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143], stage1_15[144], stage1_15[145]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[25],stage2_16[62],stage2_15[67]}
   );
   gpc606_5 gpc2516 (
      {stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149], stage1_15[150], stage1_15[151]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[26],stage2_16[63],stage2_15[68]}
   );
   gpc615_5 gpc2517 (
      {stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155], stage1_15[156]},
      {stage1_16[12]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[27],stage2_16[64],stage2_15[69]}
   );
   gpc615_5 gpc2518 (
      {stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[13]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[28],stage2_16[65],stage2_15[70]}
   );
   gpc615_5 gpc2519 (
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166]},
      {stage1_16[14]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[29],stage2_16[66],stage2_15[71]}
   );
   gpc615_5 gpc2520 (
      {stage1_15[167], stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171]},
      {stage1_16[15]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[30],stage2_16[67],stage2_15[72]}
   );
   gpc615_5 gpc2521 (
      {stage1_15[172], stage1_15[173], stage1_15[174], stage1_15[175], stage1_15[176]},
      {stage1_16[16]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[31],stage2_16[68],stage2_15[73]}
   );
   gpc615_5 gpc2522 (
      {stage1_15[177], stage1_15[178], stage1_15[179], stage1_15[180], stage1_15[181]},
      {stage1_16[17]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[32],stage2_16[69],stage2_15[74]}
   );
   gpc615_5 gpc2523 (
      {stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185], stage1_15[186]},
      {stage1_16[18]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[33],stage2_16[70],stage2_15[75]}
   );
   gpc615_5 gpc2524 (
      {stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[19]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[34],stage2_16[71],stage2_15[76]}
   );
   gpc615_5 gpc2525 (
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196]},
      {stage1_16[20]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[35],stage2_16[72],stage2_15[77]}
   );
   gpc615_5 gpc2526 (
      {stage1_15[197], stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201]},
      {stage1_16[21]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[14],stage2_17[36],stage2_16[73],stage2_15[78]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[202], stage1_15[203], stage1_15[204], stage1_15[205], stage1_15[206]},
      {stage1_16[22]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[15],stage2_17[37],stage2_16[74],stage2_15[79]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211]},
      {stage1_16[23]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[16],stage2_17[38],stage2_16[75],stage2_15[80]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216]},
      {stage1_16[24]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[17],stage2_17[39],stage2_16[76],stage2_15[81]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[25]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[18],stage2_17[40],stage2_16[77],stage2_15[82]}
   );
   gpc606_5 gpc2531 (
      {stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30], stage1_16[31]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[19],stage2_17[41],stage2_16[78]}
   );
   gpc606_5 gpc2532 (
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[20],stage2_17[42],stage2_16[79]}
   );
   gpc606_5 gpc2533 (
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[21],stage2_17[43],stage2_16[80]}
   );
   gpc606_5 gpc2534 (
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[22],stage2_17[44],stage2_16[81]}
   );
   gpc606_5 gpc2535 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[23],stage2_17[45],stage2_16[82]}
   );
   gpc606_5 gpc2536 (
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[24],stage2_17[46],stage2_16[83]}
   );
   gpc606_5 gpc2537 (
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[25],stage2_17[47],stage2_16[84]}
   );
   gpc606_5 gpc2538 (
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[26],stage2_17[48],stage2_16[85]}
   );
   gpc606_5 gpc2539 (
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[27],stage2_17[49],stage2_16[86]}
   );
   gpc606_5 gpc2540 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[28],stage2_17[50],stage2_16[87]}
   );
   gpc606_5 gpc2541 (
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[29],stage2_17[51],stage2_16[88]}
   );
   gpc606_5 gpc2542 (
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[30],stage2_17[52],stage2_16[89]}
   );
   gpc606_5 gpc2543 (
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[31],stage2_17[53],stage2_16[90]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[32],stage2_17[54],stage2_16[91]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[33],stage2_17[55],stage2_16[92]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[34],stage2_17[56],stage2_16[93]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[35],stage2_17[57],stage2_16[94]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[36],stage2_17[58],stage2_16[95]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[37],stage2_17[59],stage2_16[96]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[38],stage2_17[60],stage2_16[97]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[39],stage2_17[61],stage2_16[98]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[40],stage2_17[62],stage2_16[99]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[41],stage2_17[63],stage2_16[100]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[42],stage2_17[64],stage2_16[101]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[43],stage2_17[65],stage2_16[102]}
   );
   gpc615_5 gpc2556 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180]},
      {stage1_17[102]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[44],stage2_17[66],stage2_16[103]}
   );
   gpc615_5 gpc2557 (
      {stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage1_17[103]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[45],stage2_17[67],stage2_16[104]}
   );
   gpc615_5 gpc2558 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_17[104]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[46],stage2_17[68],stage2_16[105]}
   );
   gpc615_5 gpc2559 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195]},
      {stage1_17[105]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[47],stage2_17[69],stage2_16[106]}
   );
   gpc606_5 gpc2560 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[29],stage2_19[46],stage2_18[48],stage2_17[70]}
   );
   gpc606_5 gpc2561 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[30],stage2_19[47],stage2_18[49],stage2_17[71]}
   );
   gpc606_5 gpc2562 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[31],stage2_19[48],stage2_18[50],stage2_17[72]}
   );
   gpc606_5 gpc2563 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[32],stage2_19[49],stage2_18[51],stage2_17[73]}
   );
   gpc606_5 gpc2564 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[33],stage2_19[50],stage2_18[52],stage2_17[74]}
   );
   gpc606_5 gpc2565 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[34],stage2_19[51],stage2_18[53],stage2_17[75]}
   );
   gpc606_5 gpc2566 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[35],stage2_19[52],stage2_18[54],stage2_17[76]}
   );
   gpc606_5 gpc2567 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[36],stage2_19[53],stage2_18[55],stage2_17[77]}
   );
   gpc606_5 gpc2568 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[37],stage2_19[54],stage2_18[56],stage2_17[78]}
   );
   gpc606_5 gpc2569 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[38],stage2_19[55],stage2_18[57],stage2_17[79]}
   );
   gpc606_5 gpc2570 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[39],stage2_19[56],stage2_18[58],stage2_17[80]}
   );
   gpc606_5 gpc2571 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[40],stage2_19[57],stage2_18[59],stage2_17[81]}
   );
   gpc615_5 gpc2572 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[72]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[12],stage2_20[41],stage2_19[58],stage2_18[60]}
   );
   gpc615_5 gpc2573 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[73]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[13],stage2_20[42],stage2_19[59],stage2_18[61]}
   );
   gpc615_5 gpc2574 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[74]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[14],stage2_20[43],stage2_19[60],stage2_18[62]}
   );
   gpc615_5 gpc2575 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[75]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[15],stage2_20[44],stage2_19[61],stage2_18[63]}
   );
   gpc606_5 gpc2576 (
      {stage1_19[76], stage1_19[77], stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[16],stage2_20[45],stage2_19[62]}
   );
   gpc606_5 gpc2577 (
      {stage1_19[82], stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[17],stage2_20[46],stage2_19[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[18],stage2_20[47],stage2_19[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_19[94], stage1_19[95], stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[19],stage2_20[48],stage2_19[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_19[100], stage1_19[101], stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[20],stage2_20[49],stage2_19[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_19[106], stage1_19[107], stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[9],stage2_21[21],stage2_20[50],stage2_19[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_19[112], stage1_19[113], stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[10],stage2_21[22],stage2_20[51],stage2_19[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_19[118], stage1_19[119], stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[11],stage2_21[23],stage2_20[52],stage2_19[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_19[124], stage1_19[125], stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[12],stage2_21[24],stage2_20[53],stage2_19[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_19[130], stage1_19[131], stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[13],stage2_21[25],stage2_20[54],stage2_19[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_19[136], stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[14],stage2_21[26],stage2_20[55],stage2_19[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[15],stage2_21[27],stage2_20[56],stage2_19[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[16],stage2_21[28],stage2_20[57],stage2_19[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_19[154], stage1_19[155], stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[17],stage2_21[29],stage2_20[58],stage2_19[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_19[160], stage1_19[161], stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[18],stage2_21[30],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2591 (
      {stage1_19[166], stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170]},
      {stage1_20[24]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[19],stage2_21[31],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2592 (
      {stage1_19[171], stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175]},
      {stage1_20[25]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[20],stage2_21[32],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2593 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[26]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[21],stage2_21[33],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2594 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[27]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[22],stage2_21[34],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2595 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[28]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[23],stage2_21[35],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2596 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[29]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[24],stage2_21[36],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2597 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[30]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[25],stage2_21[37],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2598 (
      {stage1_19[201], stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205]},
      {stage1_20[31]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[26],stage2_21[38],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210]},
      {stage1_20[32]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[27],stage2_21[39],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage1_20[33]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[28],stage2_21[40],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220]},
      {stage1_20[34]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[29],stage2_21[41],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[221], stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225]},
      {stage1_20[35]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[30],stage2_21[42],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[226], stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230]},
      {stage1_20[36]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[31],stage2_21[43],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[231], stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235]},
      {stage1_20[37]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[32],stage2_21[44],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[236], stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240]},
      {stage1_20[38]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[33],stage2_21[45],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[241], stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245]},
      {stage1_20[39]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[34],stage2_21[46],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[246], stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250]},
      {stage1_20[40]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[35],stage2_21[47],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[251], stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255]},
      {stage1_20[41]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[36],stage2_21[48],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[256], stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260]},
      {stage1_20[42]},
      {stage1_21[198], stage1_21[199], stage1_21[200], stage1_21[201], stage1_21[202], stage1_21[203]},
      {stage2_23[33],stage2_22[37],stage2_21[49],stage2_20[78],stage2_19[95]}
   );
   gpc606_5 gpc2610 (
      {stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47], stage1_20[48]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[34],stage2_22[38],stage2_21[50],stage2_20[79]}
   );
   gpc606_5 gpc2611 (
      {stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53], stage1_20[54]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[35],stage2_22[39],stage2_21[51],stage2_20[80]}
   );
   gpc606_5 gpc2612 (
      {stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59], stage1_20[60]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[36],stage2_22[40],stage2_21[52],stage2_20[81]}
   );
   gpc606_5 gpc2613 (
      {stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65], stage1_20[66]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[37],stage2_22[41],stage2_21[53],stage2_20[82]}
   );
   gpc606_5 gpc2614 (
      {stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71], stage1_20[72]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[38],stage2_22[42],stage2_21[54],stage2_20[83]}
   );
   gpc606_5 gpc2615 (
      {stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77], stage1_20[78]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[39],stage2_22[43],stage2_21[55],stage2_20[84]}
   );
   gpc606_5 gpc2616 (
      {stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83], stage1_20[84]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[40],stage2_22[44],stage2_21[56],stage2_20[85]}
   );
   gpc606_5 gpc2617 (
      {stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89], stage1_20[90]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[41],stage2_22[45],stage2_21[57],stage2_20[86]}
   );
   gpc606_5 gpc2618 (
      {stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95], stage1_20[96]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[42],stage2_22[46],stage2_21[58],stage2_20[87]}
   );
   gpc606_5 gpc2619 (
      {stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101], stage1_20[102]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[43],stage2_22[47],stage2_21[59],stage2_20[88]}
   );
   gpc606_5 gpc2620 (
      {stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107], stage1_20[108]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[44],stage2_22[48],stage2_21[60],stage2_20[89]}
   );
   gpc606_5 gpc2621 (
      {stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113], stage1_20[114]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[45],stage2_22[49],stage2_21[61],stage2_20[90]}
   );
   gpc606_5 gpc2622 (
      {stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119], stage1_20[120]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[46],stage2_22[50],stage2_21[62],stage2_20[91]}
   );
   gpc606_5 gpc2623 (
      {stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125], stage1_20[126]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[47],stage2_22[51],stage2_21[63],stage2_20[92]}
   );
   gpc606_5 gpc2624 (
      {stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131], stage1_20[132]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[48],stage2_22[52],stage2_21[64],stage2_20[93]}
   );
   gpc606_5 gpc2625 (
      {stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137], stage1_20[138]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[49],stage2_22[53],stage2_21[65],stage2_20[94]}
   );
   gpc606_5 gpc2626 (
      {stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143], stage1_20[144]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[50],stage2_22[54],stage2_21[66],stage2_20[95]}
   );
   gpc606_5 gpc2627 (
      {stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149], stage1_20[150]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[51],stage2_22[55],stage2_21[67],stage2_20[96]}
   );
   gpc606_5 gpc2628 (
      {stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155], stage1_20[156]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[52],stage2_22[56],stage2_21[68],stage2_20[97]}
   );
   gpc606_5 gpc2629 (
      {stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161], stage1_20[162]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[53],stage2_22[57],stage2_21[69],stage2_20[98]}
   );
   gpc606_5 gpc2630 (
      {stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167], stage1_20[168]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[54],stage2_22[58],stage2_21[70],stage2_20[99]}
   );
   gpc606_5 gpc2631 (
      {stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173], stage1_20[174]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[55],stage2_22[59],stage2_21[71],stage2_20[100]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179], stage1_20[180]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[56],stage2_22[60],stage2_21[72],stage2_20[101]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage2_24[23],stage2_23[57],stage2_22[61],stage2_21[73],stage2_20[102]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191], stage1_20[192]},
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148], stage1_22[149]},
      {stage2_24[24],stage2_23[58],stage2_22[62],stage2_21[74],stage2_20[103]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197], stage1_20[198]},
      {stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153], stage1_22[154], stage1_22[155]},
      {stage2_24[25],stage2_23[59],stage2_22[63],stage2_21[75],stage2_20[104]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203], stage1_20[204]},
      {stage1_22[156], stage1_22[157], stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161]},
      {stage2_24[26],stage2_23[60],stage2_22[64],stage2_21[76],stage2_20[105]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[205], stage1_20[206], stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210]},
      {stage1_22[162], stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage2_24[27],stage2_23[61],stage2_22[65],stage2_21[77],stage2_20[106]}
   );
   gpc606_5 gpc2638 (
      {stage1_21[204], stage1_21[205], stage1_21[206], stage1_21[207], stage1_21[208], stage1_21[209]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[28],stage2_23[62],stage2_22[66],stage2_21[78]}
   );
   gpc606_5 gpc2639 (
      {stage1_21[210], stage1_21[211], stage1_21[212], stage1_21[213], stage1_21[214], stage1_21[215]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[29],stage2_23[63],stage2_22[67],stage2_21[79]}
   );
   gpc606_5 gpc2640 (
      {stage1_21[216], stage1_21[217], stage1_21[218], stage1_21[219], stage1_21[220], stage1_21[221]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[30],stage2_23[64],stage2_22[68],stage2_21[80]}
   );
   gpc615_5 gpc2641 (
      {stage1_21[222], stage1_21[223], stage1_21[224], stage1_21[225], stage1_21[226]},
      {stage1_22[168]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[31],stage2_23[65],stage2_22[69],stage2_21[81]}
   );
   gpc606_5 gpc2642 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173], stage1_22[174]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[32],stage2_23[66],stage2_22[70]}
   );
   gpc606_5 gpc2643 (
      {stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178], stage1_22[179], stage1_22[180]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[33],stage2_23[67],stage2_22[71]}
   );
   gpc606_5 gpc2644 (
      {stage1_22[181], stage1_22[182], stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[34],stage2_23[68],stage2_22[72]}
   );
   gpc606_5 gpc2645 (
      {stage1_22[187], stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[35],stage2_23[69],stage2_22[73]}
   );
   gpc615_5 gpc2646 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[24]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[36],stage2_23[70],stage2_22[74]}
   );
   gpc615_5 gpc2647 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[25]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[37],stage2_23[71],stage2_22[75]}
   );
   gpc615_5 gpc2648 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[26]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[38],stage2_23[72],stage2_22[76]}
   );
   gpc615_5 gpc2649 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[27]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[39],stage2_23[73],stage2_22[77]}
   );
   gpc615_5 gpc2650 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[28]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[40],stage2_23[74],stage2_22[78]}
   );
   gpc615_5 gpc2651 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[29]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[41],stage2_23[75],stage2_22[79]}
   );
   gpc615_5 gpc2652 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[30]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[42],stage2_23[76],stage2_22[80]}
   );
   gpc615_5 gpc2653 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[31]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[43],stage2_23[77],stage2_22[81]}
   );
   gpc615_5 gpc2654 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[32]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[44],stage2_23[78],stage2_22[82]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[33]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[17],stage2_24[45],stage2_23[79],stage2_22[83]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[34]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[18],stage2_24[46],stage2_23[80],stage2_22[84]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[248], stage1_22[249], stage1_22[250], stage1_22[251], stage1_22[252]},
      {stage1_23[35]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[19],stage2_24[47],stage2_23[81],stage2_22[85]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[253], stage1_22[254], stage1_22[255], stage1_22[256], stage1_22[257]},
      {stage1_23[36]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[20],stage2_24[48],stage2_23[82],stage2_22[86]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[258], stage1_22[259], stage1_22[260], stage1_22[261], stage1_22[262]},
      {stage1_23[37]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[21],stage2_24[49],stage2_23[83],stage2_22[87]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[263], stage1_22[264], stage1_22[265], stage1_22[266], stage1_22[267]},
      {stage1_23[38]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[22],stage2_24[50],stage2_23[84],stage2_22[88]}
   );
   gpc606_5 gpc2661 (
      {stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42], stage1_23[43], stage1_23[44]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[19],stage2_25[23],stage2_24[51],stage2_23[85]}
   );
   gpc606_5 gpc2662 (
      {stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48], stage1_23[49], stage1_23[50]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[20],stage2_25[24],stage2_24[52],stage2_23[86]}
   );
   gpc606_5 gpc2663 (
      {stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[21],stage2_25[25],stage2_24[53],stage2_23[87]}
   );
   gpc606_5 gpc2664 (
      {stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[22],stage2_25[26],stage2_24[54],stage2_23[88]}
   );
   gpc606_5 gpc2665 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67], stage1_23[68]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[23],stage2_25[27],stage2_24[55],stage2_23[89]}
   );
   gpc606_5 gpc2666 (
      {stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72], stage1_23[73], stage1_23[74]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[24],stage2_25[28],stage2_24[56],stage2_23[90]}
   );
   gpc606_5 gpc2667 (
      {stage1_23[75], stage1_23[76], stage1_23[77], stage1_23[78], stage1_23[79], stage1_23[80]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[25],stage2_25[29],stage2_24[57],stage2_23[91]}
   );
   gpc606_5 gpc2668 (
      {stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[26],stage2_25[30],stage2_24[58],stage2_23[92]}
   );
   gpc606_5 gpc2669 (
      {stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[27],stage2_25[31],stage2_24[59],stage2_23[93]}
   );
   gpc606_5 gpc2670 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97], stage1_23[98]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[28],stage2_25[32],stage2_24[60],stage2_23[94]}
   );
   gpc606_5 gpc2671 (
      {stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102], stage1_23[103], stage1_23[104]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[29],stage2_25[33],stage2_24[61],stage2_23[95]}
   );
   gpc606_5 gpc2672 (
      {stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108], stage1_23[109], stage1_23[110]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[30],stage2_25[34],stage2_24[62],stage2_23[96]}
   );
   gpc606_5 gpc2673 (
      {stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[31],stage2_25[35],stage2_24[63],stage2_23[97]}
   );
   gpc606_5 gpc2674 (
      {stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[32],stage2_25[36],stage2_24[64],stage2_23[98]}
   );
   gpc606_5 gpc2675 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127], stage1_23[128]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[33],stage2_25[37],stage2_24[65],stage2_23[99]}
   );
   gpc606_5 gpc2676 (
      {stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132], stage1_23[133], stage1_23[134]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[34],stage2_25[38],stage2_24[66],stage2_23[100]}
   );
   gpc606_5 gpc2677 (
      {stage1_23[135], stage1_23[136], stage1_23[137], stage1_23[138], stage1_23[139], stage1_23[140]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[35],stage2_25[39],stage2_24[67],stage2_23[101]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[141], stage1_23[142], stage1_23[143], stage1_23[144], stage1_23[145]},
      {stage1_24[114]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[36],stage2_25[40],stage2_24[68],stage2_23[102]}
   );
   gpc606_5 gpc2679 (
      {stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119], stage1_24[120]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[18],stage2_26[37],stage2_25[41],stage2_24[69]}
   );
   gpc606_5 gpc2680 (
      {stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125], stage1_24[126]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[19],stage2_26[38],stage2_25[42],stage2_24[70]}
   );
   gpc606_5 gpc2681 (
      {stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[20],stage2_26[39],stage2_25[43],stage2_24[71]}
   );
   gpc606_5 gpc2682 (
      {stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[21],stage2_26[40],stage2_25[44],stage2_24[72]}
   );
   gpc606_5 gpc2683 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143], stage1_24[144]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[22],stage2_26[41],stage2_25[45],stage2_24[73]}
   );
   gpc606_5 gpc2684 (
      {stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149], stage1_24[150]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[23],stage2_26[42],stage2_25[46],stage2_24[74]}
   );
   gpc606_5 gpc2685 (
      {stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155], stage1_24[156]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[24],stage2_26[43],stage2_25[47],stage2_24[75]}
   );
   gpc606_5 gpc2686 (
      {stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[25],stage2_26[44],stage2_25[48],stage2_24[76]}
   );
   gpc606_5 gpc2687 (
      {stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[26],stage2_26[45],stage2_25[49],stage2_24[77]}
   );
   gpc606_5 gpc2688 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173], stage1_24[174]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[27],stage2_26[46],stage2_25[50],stage2_24[78]}
   );
   gpc606_5 gpc2689 (
      {stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179], stage1_24[180]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[28],stage2_26[47],stage2_25[51],stage2_24[79]}
   );
   gpc606_5 gpc2690 (
      {stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185], stage1_24[186]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[29],stage2_26[48],stage2_25[52],stage2_24[80]}
   );
   gpc606_5 gpc2691 (
      {stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[30],stage2_26[49],stage2_25[53],stage2_24[81]}
   );
   gpc606_5 gpc2692 (
      {stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[31],stage2_26[50],stage2_25[54],stage2_24[82]}
   );
   gpc606_5 gpc2693 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203], stage1_24[204]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[32],stage2_26[51],stage2_25[55],stage2_24[83]}
   );
   gpc606_5 gpc2694 (
      {stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209], stage1_24[210]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[33],stage2_26[52],stage2_25[56],stage2_24[84]}
   );
   gpc606_5 gpc2695 (
      {stage1_24[211], stage1_24[212], stage1_24[213], stage1_24[214], stage1_24[215], stage1_24[216]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[34],stage2_26[53],stage2_25[57],stage2_24[85]}
   );
   gpc606_5 gpc2696 (
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[17],stage2_27[35],stage2_26[54],stage2_25[58]}
   );
   gpc606_5 gpc2697 (
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[18],stage2_27[36],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc2698 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[19],stage2_27[37],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc2699 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[20],stage2_27[38],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc2700 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[21],stage2_27[39],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc2701 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[22],stage2_27[40],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc2702 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[23],stage2_27[41],stage2_26[60],stage2_25[64]}
   );
   gpc606_5 gpc2703 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[24],stage2_27[42],stage2_26[61],stage2_25[65]}
   );
   gpc606_5 gpc2704 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[25],stage2_27[43],stage2_26[62],stage2_25[66]}
   );
   gpc606_5 gpc2705 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[26],stage2_27[44],stage2_26[63],stage2_25[67]}
   );
   gpc606_5 gpc2706 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64], stage1_27[65]},
      {stage2_29[10],stage2_28[27],stage2_27[45],stage2_26[64],stage2_25[68]}
   );
   gpc606_5 gpc2707 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71]},
      {stage2_29[11],stage2_28[28],stage2_27[46],stage2_26[65],stage2_25[69]}
   );
   gpc606_5 gpc2708 (
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage1_27[72], stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage2_29[12],stage2_28[29],stage2_27[47],stage2_26[66],stage2_25[70]}
   );
   gpc606_5 gpc2709 (
      {stage1_25[186], stage1_25[187], stage1_25[188], stage1_25[189], stage1_25[190], stage1_25[191]},
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83]},
      {stage2_29[13],stage2_28[30],stage2_27[48],stage2_26[67],stage2_25[71]}
   );
   gpc606_5 gpc2710 (
      {stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196], stage1_25[197]},
      {stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage2_29[14],stage2_28[31],stage2_27[49],stage2_26[68],stage2_25[72]}
   );
   gpc606_5 gpc2711 (
      {stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202], stage1_25[203]},
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage2_29[15],stage2_28[32],stage2_27[50],stage2_26[69],stage2_25[73]}
   );
   gpc606_5 gpc2712 (
      {stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208], stage1_25[209]},
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101]},
      {stage2_29[16],stage2_28[33],stage2_27[51],stage2_26[70],stage2_25[74]}
   );
   gpc615_5 gpc2713 (
      {stage1_25[210], stage1_25[211], stage1_25[212], stage1_25[213], stage1_25[214]},
      {stage1_26[102]},
      {stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage2_29[17],stage2_28[34],stage2_27[52],stage2_26[71],stage2_25[75]}
   );
   gpc615_5 gpc2714 (
      {stage1_25[215], stage1_25[216], stage1_25[217], stage1_25[218], stage1_25[219]},
      {stage1_26[103]},
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113]},
      {stage2_29[18],stage2_28[35],stage2_27[53],stage2_26[72],stage2_25[76]}
   );
   gpc615_5 gpc2715 (
      {stage1_25[220], stage1_25[221], stage1_25[222], stage1_25[223], stage1_25[224]},
      {stage1_26[104]},
      {stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage2_29[19],stage2_28[36],stage2_27[54],stage2_26[73],stage2_25[77]}
   );
   gpc615_5 gpc2716 (
      {stage1_25[225], stage1_25[226], stage1_25[227], stage1_25[228], stage1_25[229]},
      {stage1_26[105]},
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage2_29[20],stage2_28[37],stage2_27[55],stage2_26[74],stage2_25[78]}
   );
   gpc615_5 gpc2717 (
      {stage1_25[230], stage1_25[231], stage1_25[232], stage1_25[233], stage1_25[234]},
      {stage1_26[106]},
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131]},
      {stage2_29[21],stage2_28[38],stage2_27[56],stage2_26[75],stage2_25[79]}
   );
   gpc615_5 gpc2718 (
      {stage1_25[235], stage1_25[236], stage1_25[237], stage1_25[238], stage1_25[239]},
      {stage1_26[107]},
      {stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage2_29[22],stage2_28[39],stage2_27[57],stage2_26[76],stage2_25[80]}
   );
   gpc615_5 gpc2719 (
      {stage1_25[240], stage1_25[241], stage1_25[242], stage1_25[243], stage1_25[244]},
      {stage1_26[108]},
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143]},
      {stage2_29[23],stage2_28[40],stage2_27[58],stage2_26[77],stage2_25[81]}
   );
   gpc615_5 gpc2720 (
      {stage1_25[245], stage1_25[246], stage1_25[247], stage1_25[248], stage1_25[249]},
      {stage1_26[109]},
      {stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage2_29[24],stage2_28[41],stage2_27[59],stage2_26[78],stage2_25[82]}
   );
   gpc615_5 gpc2721 (
      {stage1_25[250], stage1_25[251], stage1_25[252], stage1_25[253], stage1_25[254]},
      {stage1_26[110]},
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage2_29[25],stage2_28[42],stage2_27[60],stage2_26[79],stage2_25[83]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[156]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[26],stage2_28[43],stage2_27[61],stage2_26[80]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[157]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[27],stage2_28[44],stage2_27[62],stage2_26[81]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[158]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[28],stage2_28[45],stage2_27[63],stage2_26[82]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[159]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[29],stage2_28[46],stage2_27[64],stage2_26[83]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[160]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[30],stage2_28[47],stage2_27[65],stage2_26[84]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[161]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[31],stage2_28[48],stage2_27[66],stage2_26[85]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[162]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[32],stage2_28[49],stage2_27[67],stage2_26[86]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[163]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[33],stage2_28[50],stage2_27[68],stage2_26[87]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage1_27[164]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[34],stage2_28[51],stage2_27[69],stage2_26[88]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160]},
      {stage1_27[165]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[35],stage2_28[52],stage2_27[70],stage2_26[89]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165]},
      {stage1_27[166]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[36],stage2_28[53],stage2_27[71],stage2_26[90]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169], stage1_26[170]},
      {stage1_27[167]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[37],stage2_28[54],stage2_27[72],stage2_26[91]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174], stage1_26[175]},
      {stage1_27[168]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[38],stage2_28[55],stage2_27[73],stage2_26[92]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179], stage1_26[180]},
      {stage1_27[169]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[39],stage2_28[56],stage2_27[74],stage2_26[93]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage1_27[170]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[40],stage2_28[57],stage2_27[75],stage2_26[94]}
   );
   gpc615_5 gpc2737 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[90]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[15],stage2_29[41],stage2_28[58],stage2_27[76]}
   );
   gpc615_5 gpc2738 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[91]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[16],stage2_29[42],stage2_28[59],stage2_27[77]}
   );
   gpc615_5 gpc2739 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[92]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[17],stage2_29[43],stage2_28[60],stage2_27[78]}
   );
   gpc615_5 gpc2740 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[93]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[18],stage2_29[44],stage2_28[61],stage2_27[79]}
   );
   gpc615_5 gpc2741 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[94]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[19],stage2_29[45],stage2_28[62],stage2_27[80]}
   );
   gpc606_5 gpc2742 (
      {stage1_28[95], stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[5],stage2_30[20],stage2_29[46],stage2_28[63]}
   );
   gpc606_5 gpc2743 (
      {stage1_28[101], stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[6],stage2_30[21],stage2_29[47],stage2_28[64]}
   );
   gpc606_5 gpc2744 (
      {stage1_28[107], stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[7],stage2_30[22],stage2_29[48],stage2_28[65]}
   );
   gpc606_5 gpc2745 (
      {stage1_28[113], stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[8],stage2_30[23],stage2_29[49],stage2_28[66]}
   );
   gpc606_5 gpc2746 (
      {stage1_28[119], stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[9],stage2_30[24],stage2_29[50],stage2_28[67]}
   );
   gpc606_5 gpc2747 (
      {stage1_28[125], stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[10],stage2_30[25],stage2_29[51],stage2_28[68]}
   );
   gpc606_5 gpc2748 (
      {stage1_28[131], stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[11],stage2_30[26],stage2_29[52],stage2_28[69]}
   );
   gpc606_5 gpc2749 (
      {stage1_28[137], stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[12],stage2_30[27],stage2_29[53],stage2_28[70]}
   );
   gpc606_5 gpc2750 (
      {stage1_28[143], stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[13],stage2_30[28],stage2_29[54],stage2_28[71]}
   );
   gpc606_5 gpc2751 (
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[9],stage2_31[14],stage2_30[29],stage2_29[55]}
   );
   gpc606_5 gpc2752 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[10],stage2_31[15],stage2_30[30],stage2_29[56]}
   );
   gpc606_5 gpc2753 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[11],stage2_31[16],stage2_30[31],stage2_29[57]}
   );
   gpc606_5 gpc2754 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[12],stage2_31[17],stage2_30[32],stage2_29[58]}
   );
   gpc606_5 gpc2755 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[13],stage2_31[18],stage2_30[33],stage2_29[59]}
   );
   gpc606_5 gpc2756 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[14],stage2_31[19],stage2_30[34],stage2_29[60]}
   );
   gpc606_5 gpc2757 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[15],stage2_31[20],stage2_30[35],stage2_29[61]}
   );
   gpc606_5 gpc2758 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[16],stage2_31[21],stage2_30[36],stage2_29[62]}
   );
   gpc606_5 gpc2759 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[17],stage2_31[22],stage2_30[37],stage2_29[63]}
   );
   gpc606_5 gpc2760 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[18],stage2_31[23],stage2_30[38],stage2_29[64]}
   );
   gpc606_5 gpc2761 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[19],stage2_31[24],stage2_30[39],stage2_29[65]}
   );
   gpc606_5 gpc2762 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[20],stage2_31[25],stage2_30[40],stage2_29[66]}
   );
   gpc606_5 gpc2763 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[21],stage2_31[26],stage2_30[41],stage2_29[67]}
   );
   gpc606_5 gpc2764 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[22],stage2_31[27],stage2_30[42],stage2_29[68]}
   );
   gpc606_5 gpc2765 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage2_33[14],stage2_32[23],stage2_31[28],stage2_30[43],stage2_29[69]}
   );
   gpc606_5 gpc2766 (
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage2_33[15],stage2_32[24],stage2_31[29],stage2_30[44],stage2_29[70]}
   );
   gpc606_5 gpc2767 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage2_33[16],stage2_32[25],stage2_31[30],stage2_30[45],stage2_29[71]}
   );
   gpc606_5 gpc2768 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage2_33[17],stage2_32[26],stage2_31[31],stage2_30[46],stage2_29[72]}
   );
   gpc606_5 gpc2769 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage2_33[18],stage2_32[27],stage2_31[32],stage2_30[47],stage2_29[73]}
   );
   gpc606_5 gpc2770 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage2_33[19],stage2_32[28],stage2_31[33],stage2_30[48],stage2_29[74]}
   );
   gpc606_5 gpc2771 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage2_33[20],stage2_32[29],stage2_31[34],stage2_30[49],stage2_29[75]}
   );
   gpc606_5 gpc2772 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage2_33[21],stage2_32[30],stage2_31[35],stage2_30[50],stage2_29[76]}
   );
   gpc606_5 gpc2773 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage2_33[22],stage2_32[31],stage2_31[36],stage2_30[51],stage2_29[77]}
   );
   gpc606_5 gpc2774 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage2_33[23],stage2_32[32],stage2_31[37],stage2_30[52],stage2_29[78]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[144], stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage2_33[24],stage2_32[33],stage2_31[38],stage2_30[53],stage2_29[79]}
   );
   gpc606_5 gpc2776 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[25],stage2_32[34],stage2_31[39],stage2_30[54]}
   );
   gpc606_5 gpc2777 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[26],stage2_32[35],stage2_31[40],stage2_30[55]}
   );
   gpc606_5 gpc2778 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[27],stage2_32[36],stage2_31[41],stage2_30[56]}
   );
   gpc606_5 gpc2779 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[28],stage2_32[37],stage2_31[42],stage2_30[57]}
   );
   gpc606_5 gpc2780 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[29],stage2_32[38],stage2_31[43],stage2_30[58]}
   );
   gpc606_5 gpc2781 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[30],stage2_32[39],stage2_31[44],stage2_30[59]}
   );
   gpc606_5 gpc2782 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[31],stage2_32[40],stage2_31[45],stage2_30[60]}
   );
   gpc606_5 gpc2783 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[32],stage2_32[41],stage2_31[46],stage2_30[61]}
   );
   gpc606_5 gpc2784 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[33],stage2_32[42],stage2_31[47],stage2_30[62]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[34],stage2_32[43],stage2_31[48],stage2_30[63]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[35],stage2_32[44],stage2_31[49],stage2_30[64]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[36],stage2_32[45],stage2_31[50],stage2_30[65]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[37],stage2_32[46],stage2_31[51],stage2_30[66]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135], stage1_30[136], stage1_30[137]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[38],stage2_32[47],stage2_31[52],stage2_30[67]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[39],stage2_32[48],stage2_31[53],stage2_30[68]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[40],stage2_32[49],stage2_31[54],stage2_30[69]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154], stage1_30[155]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[41],stage2_32[50],stage2_31[55],stage2_30[70]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159], stage1_30[160], stage1_30[161]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[42],stage2_32[51],stage2_31[56],stage2_30[71]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165], stage1_30[166], stage1_30[167]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[43],stage2_32[52],stage2_31[57],stage2_30[72]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171], stage1_30[172], stage1_30[173]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[44],stage2_32[53],stage2_31[58],stage2_30[73]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177], stage1_30[178], stage1_30[179]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[45],stage2_32[54],stage2_31[59],stage2_30[74]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183], stage1_30[184], stage1_30[185]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[46],stage2_32[55],stage2_31[60],stage2_30[75]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189], stage1_30[190], stage1_30[191]},
      {stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136], stage1_32[137]},
      {stage2_34[22],stage2_33[47],stage2_32[56],stage2_31[61],stage2_30[76]}
   );
   gpc606_5 gpc2799 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154], stage1_31[155]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[23],stage2_33[48],stage2_32[57],stage2_31[62]}
   );
   gpc606_5 gpc2800 (
      {stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159], stage1_31[160], stage1_31[161]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[24],stage2_33[49],stage2_32[58],stage2_31[63]}
   );
   gpc606_5 gpc2801 (
      {stage1_31[162], stage1_31[163], stage1_31[164], stage1_31[165], stage1_31[166], stage1_31[167]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[25],stage2_33[50],stage2_32[59],stage2_31[64]}
   );
   gpc606_5 gpc2802 (
      {stage1_31[168], stage1_31[169], stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[26],stage2_33[51],stage2_32[60],stage2_31[65]}
   );
   gpc606_5 gpc2803 (
      {stage1_31[174], stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[27],stage2_33[52],stage2_32[61],stage2_31[66]}
   );
   gpc615_5 gpc2804 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[138]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[28],stage2_33[53],stage2_32[62],stage2_31[67]}
   );
   gpc615_5 gpc2805 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[139]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[29],stage2_33[54],stage2_32[63],stage2_31[68]}
   );
   gpc615_5 gpc2806 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[140]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[30],stage2_33[55],stage2_32[64],stage2_31[69]}
   );
   gpc615_5 gpc2807 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[141]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[31],stage2_33[56],stage2_32[65],stage2_31[70]}
   );
   gpc615_5 gpc2808 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[142]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[32],stage2_33[57],stage2_32[66],stage2_31[71]}
   );
   gpc615_5 gpc2809 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[143]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[33],stage2_33[58],stage2_32[67],stage2_31[72]}
   );
   gpc615_5 gpc2810 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[144]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], 1'b0},
      {stage2_35[11],stage2_34[34],stage2_33[59],stage2_32[68],stage2_31[73]}
   );
   gpc1_1 gpc2811 (
      {stage1_0[60]},
      {stage2_0[12]}
   );
   gpc1_1 gpc2812 (
      {stage1_0[61]},
      {stage2_0[13]}
   );
   gpc1_1 gpc2813 (
      {stage1_0[62]},
      {stage2_0[14]}
   );
   gpc1_1 gpc2814 (
      {stage1_0[63]},
      {stage2_0[15]}
   );
   gpc1_1 gpc2815 (
      {stage1_0[64]},
      {stage2_0[16]}
   );
   gpc1_1 gpc2816 (
      {stage1_0[65]},
      {stage2_0[17]}
   );
   gpc1_1 gpc2817 (
      {stage1_0[66]},
      {stage2_0[18]}
   );
   gpc1_1 gpc2818 (
      {stage1_0[67]},
      {stage2_0[19]}
   );
   gpc1_1 gpc2819 (
      {stage1_0[68]},
      {stage2_0[20]}
   );
   gpc1_1 gpc2820 (
      {stage1_0[69]},
      {stage2_0[21]}
   );
   gpc1_1 gpc2821 (
      {stage1_0[70]},
      {stage2_0[22]}
   );
   gpc1_1 gpc2822 (
      {stage1_0[71]},
      {stage2_0[23]}
   );
   gpc1_1 gpc2823 (
      {stage1_0[72]},
      {stage2_0[24]}
   );
   gpc1_1 gpc2824 (
      {stage1_0[73]},
      {stage2_0[25]}
   );
   gpc1_1 gpc2825 (
      {stage1_0[74]},
      {stage2_0[26]}
   );
   gpc1_1 gpc2826 (
      {stage1_0[75]},
      {stage2_0[27]}
   );
   gpc1_1 gpc2827 (
      {stage1_0[76]},
      {stage2_0[28]}
   );
   gpc1_1 gpc2828 (
      {stage1_0[77]},
      {stage2_0[29]}
   );
   gpc1_1 gpc2829 (
      {stage1_0[78]},
      {stage2_0[30]}
   );
   gpc1_1 gpc2830 (
      {stage1_0[79]},
      {stage2_0[31]}
   );
   gpc1_1 gpc2831 (
      {stage1_0[80]},
      {stage2_0[32]}
   );
   gpc1_1 gpc2832 (
      {stage1_0[81]},
      {stage2_0[33]}
   );
   gpc1_1 gpc2833 (
      {stage1_0[82]},
      {stage2_0[34]}
   );
   gpc1_1 gpc2834 (
      {stage1_0[83]},
      {stage2_0[35]}
   );
   gpc1_1 gpc2835 (
      {stage1_0[84]},
      {stage2_0[36]}
   );
   gpc1_1 gpc2836 (
      {stage1_0[85]},
      {stage2_0[37]}
   );
   gpc1_1 gpc2837 (
      {stage1_0[86]},
      {stage2_0[38]}
   );
   gpc1_1 gpc2838 (
      {stage1_0[87]},
      {stage2_0[39]}
   );
   gpc1_1 gpc2839 (
      {stage1_0[88]},
      {stage2_0[40]}
   );
   gpc1_1 gpc2840 (
      {stage1_0[89]},
      {stage2_0[41]}
   );
   gpc1_1 gpc2841 (
      {stage1_0[90]},
      {stage2_0[42]}
   );
   gpc1_1 gpc2842 (
      {stage1_0[91]},
      {stage2_0[43]}
   );
   gpc1_1 gpc2843 (
      {stage1_0[92]},
      {stage2_0[44]}
   );
   gpc1_1 gpc2844 (
      {stage1_0[93]},
      {stage2_0[45]}
   );
   gpc1_1 gpc2845 (
      {stage1_0[94]},
      {stage2_0[46]}
   );
   gpc1_1 gpc2846 (
      {stage1_0[95]},
      {stage2_0[47]}
   );
   gpc1_1 gpc2847 (
      {stage1_0[96]},
      {stage2_0[48]}
   );
   gpc1_1 gpc2848 (
      {stage1_0[97]},
      {stage2_0[49]}
   );
   gpc1_1 gpc2849 (
      {stage1_0[98]},
      {stage2_0[50]}
   );
   gpc1_1 gpc2850 (
      {stage1_0[99]},
      {stage2_0[51]}
   );
   gpc1_1 gpc2851 (
      {stage1_0[100]},
      {stage2_0[52]}
   );
   gpc1_1 gpc2852 (
      {stage1_0[101]},
      {stage2_0[53]}
   );
   gpc1_1 gpc2853 (
      {stage1_0[102]},
      {stage2_0[54]}
   );
   gpc1_1 gpc2854 (
      {stage1_0[103]},
      {stage2_0[55]}
   );
   gpc1_1 gpc2855 (
      {stage1_0[104]},
      {stage2_0[56]}
   );
   gpc1_1 gpc2856 (
      {stage1_0[105]},
      {stage2_0[57]}
   );
   gpc1_1 gpc2857 (
      {stage1_0[106]},
      {stage2_0[58]}
   );
   gpc1_1 gpc2858 (
      {stage1_0[107]},
      {stage2_0[59]}
   );
   gpc1_1 gpc2859 (
      {stage1_0[108]},
      {stage2_0[60]}
   );
   gpc1_1 gpc2860 (
      {stage1_0[109]},
      {stage2_0[61]}
   );
   gpc1_1 gpc2861 (
      {stage1_0[110]},
      {stage2_0[62]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[182]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[183]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[184]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[185]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[186]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[187]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[188]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[189]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[190]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[191]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[192]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[193]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[194]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[195]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[196]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[197]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[198]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2879 (
      {stage1_2[152]},
      {stage2_2[59]}
   );
   gpc1_1 gpc2880 (
      {stage1_2[153]},
      {stage2_2[60]}
   );
   gpc1_1 gpc2881 (
      {stage1_2[154]},
      {stage2_2[61]}
   );
   gpc1_1 gpc2882 (
      {stage1_2[155]},
      {stage2_2[62]}
   );
   gpc1_1 gpc2883 (
      {stage1_2[156]},
      {stage2_2[63]}
   );
   gpc1_1 gpc2884 (
      {stage1_2[157]},
      {stage2_2[64]}
   );
   gpc1_1 gpc2885 (
      {stage1_2[158]},
      {stage2_2[65]}
   );
   gpc1_1 gpc2886 (
      {stage1_2[159]},
      {stage2_2[66]}
   );
   gpc1_1 gpc2887 (
      {stage1_2[160]},
      {stage2_2[67]}
   );
   gpc1_1 gpc2888 (
      {stage1_2[161]},
      {stage2_2[68]}
   );
   gpc1_1 gpc2889 (
      {stage1_2[162]},
      {stage2_2[69]}
   );
   gpc1_1 gpc2890 (
      {stage1_2[163]},
      {stage2_2[70]}
   );
   gpc1_1 gpc2891 (
      {stage1_2[164]},
      {stage2_2[71]}
   );
   gpc1_1 gpc2892 (
      {stage1_2[165]},
      {stage2_2[72]}
   );
   gpc1_1 gpc2893 (
      {stage1_2[166]},
      {stage2_2[73]}
   );
   gpc1_1 gpc2894 (
      {stage1_2[167]},
      {stage2_2[74]}
   );
   gpc1_1 gpc2895 (
      {stage1_2[168]},
      {stage2_2[75]}
   );
   gpc1_1 gpc2896 (
      {stage1_2[169]},
      {stage2_2[76]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[170]},
      {stage2_2[77]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[171]},
      {stage2_2[78]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[172]},
      {stage2_2[79]}
   );
   gpc1_1 gpc2900 (
      {stage1_2[173]},
      {stage2_2[80]}
   );
   gpc1_1 gpc2901 (
      {stage1_2[174]},
      {stage2_2[81]}
   );
   gpc1_1 gpc2902 (
      {stage1_2[175]},
      {stage2_2[82]}
   );
   gpc1_1 gpc2903 (
      {stage1_2[176]},
      {stage2_2[83]}
   );
   gpc1_1 gpc2904 (
      {stage1_2[177]},
      {stage2_2[84]}
   );
   gpc1_1 gpc2905 (
      {stage1_2[178]},
      {stage2_2[85]}
   );
   gpc1_1 gpc2906 (
      {stage1_2[179]},
      {stage2_2[86]}
   );
   gpc1_1 gpc2907 (
      {stage1_2[180]},
      {stage2_2[87]}
   );
   gpc1_1 gpc2908 (
      {stage1_2[181]},
      {stage2_2[88]}
   );
   gpc1_1 gpc2909 (
      {stage1_2[182]},
      {stage2_2[89]}
   );
   gpc1_1 gpc2910 (
      {stage1_2[183]},
      {stage2_2[90]}
   );
   gpc1_1 gpc2911 (
      {stage1_2[184]},
      {stage2_2[91]}
   );
   gpc1_1 gpc2912 (
      {stage1_2[185]},
      {stage2_2[92]}
   );
   gpc1_1 gpc2913 (
      {stage1_2[186]},
      {stage2_2[93]}
   );
   gpc1_1 gpc2914 (
      {stage1_2[187]},
      {stage2_2[94]}
   );
   gpc1_1 gpc2915 (
      {stage1_4[217]},
      {stage2_4[91]}
   );
   gpc1_1 gpc2916 (
      {stage1_4[218]},
      {stage2_4[92]}
   );
   gpc1_1 gpc2917 (
      {stage1_4[219]},
      {stage2_4[93]}
   );
   gpc1_1 gpc2918 (
      {stage1_4[220]},
      {stage2_4[94]}
   );
   gpc1_1 gpc2919 (
      {stage1_4[221]},
      {stage2_4[95]}
   );
   gpc1_1 gpc2920 (
      {stage1_4[222]},
      {stage2_4[96]}
   );
   gpc1_1 gpc2921 (
      {stage1_4[223]},
      {stage2_4[97]}
   );
   gpc1_1 gpc2922 (
      {stage1_4[224]},
      {stage2_4[98]}
   );
   gpc1_1 gpc2923 (
      {stage1_4[225]},
      {stage2_4[99]}
   );
   gpc1_1 gpc2924 (
      {stage1_4[226]},
      {stage2_4[100]}
   );
   gpc1_1 gpc2925 (
      {stage1_4[227]},
      {stage2_4[101]}
   );
   gpc1_1 gpc2926 (
      {stage1_4[228]},
      {stage2_4[102]}
   );
   gpc1_1 gpc2927 (
      {stage1_4[229]},
      {stage2_4[103]}
   );
   gpc1_1 gpc2928 (
      {stage1_4[230]},
      {stage2_4[104]}
   );
   gpc1_1 gpc2929 (
      {stage1_4[231]},
      {stage2_4[105]}
   );
   gpc1_1 gpc2930 (
      {stage1_4[232]},
      {stage2_4[106]}
   );
   gpc1_1 gpc2931 (
      {stage1_4[233]},
      {stage2_4[107]}
   );
   gpc1_1 gpc2932 (
      {stage1_4[234]},
      {stage2_4[108]}
   );
   gpc1_1 gpc2933 (
      {stage1_4[235]},
      {stage2_4[109]}
   );
   gpc1_1 gpc2934 (
      {stage1_4[236]},
      {stage2_4[110]}
   );
   gpc1_1 gpc2935 (
      {stage1_4[237]},
      {stage2_4[111]}
   );
   gpc1_1 gpc2936 (
      {stage1_4[238]},
      {stage2_4[112]}
   );
   gpc1_1 gpc2937 (
      {stage1_4[239]},
      {stage2_4[113]}
   );
   gpc1_1 gpc2938 (
      {stage1_4[240]},
      {stage2_4[114]}
   );
   gpc1_1 gpc2939 (
      {stage1_4[241]},
      {stage2_4[115]}
   );
   gpc1_1 gpc2940 (
      {stage1_4[242]},
      {stage2_4[116]}
   );
   gpc1_1 gpc2941 (
      {stage1_4[243]},
      {stage2_4[117]}
   );
   gpc1_1 gpc2942 (
      {stage1_4[244]},
      {stage2_4[118]}
   );
   gpc1_1 gpc2943 (
      {stage1_7[166]},
      {stage2_7[89]}
   );
   gpc1_1 gpc2944 (
      {stage1_7[167]},
      {stage2_7[90]}
   );
   gpc1_1 gpc2945 (
      {stage1_7[168]},
      {stage2_7[91]}
   );
   gpc1_1 gpc2946 (
      {stage1_7[169]},
      {stage2_7[92]}
   );
   gpc1_1 gpc2947 (
      {stage1_7[170]},
      {stage2_7[93]}
   );
   gpc1_1 gpc2948 (
      {stage1_7[171]},
      {stage2_7[94]}
   );
   gpc1_1 gpc2949 (
      {stage1_7[172]},
      {stage2_7[95]}
   );
   gpc1_1 gpc2950 (
      {stage1_7[173]},
      {stage2_7[96]}
   );
   gpc1_1 gpc2951 (
      {stage1_7[174]},
      {stage2_7[97]}
   );
   gpc1_1 gpc2952 (
      {stage1_7[175]},
      {stage2_7[98]}
   );
   gpc1_1 gpc2953 (
      {stage1_7[176]},
      {stage2_7[99]}
   );
   gpc1_1 gpc2954 (
      {stage1_7[177]},
      {stage2_7[100]}
   );
   gpc1_1 gpc2955 (
      {stage1_7[178]},
      {stage2_7[101]}
   );
   gpc1_1 gpc2956 (
      {stage1_7[179]},
      {stage2_7[102]}
   );
   gpc1_1 gpc2957 (
      {stage1_7[180]},
      {stage2_7[103]}
   );
   gpc1_1 gpc2958 (
      {stage1_7[181]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2959 (
      {stage1_7[182]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2960 (
      {stage1_7[183]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2961 (
      {stage1_7[184]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2962 (
      {stage1_7[185]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2963 (
      {stage1_9[210]},
      {stage2_9[106]}
   );
   gpc1_1 gpc2964 (
      {stage1_9[211]},
      {stage2_9[107]}
   );
   gpc1_1 gpc2965 (
      {stage1_11[161]},
      {stage2_11[71]}
   );
   gpc1_1 gpc2966 (
      {stage1_11[162]},
      {stage2_11[72]}
   );
   gpc1_1 gpc2967 (
      {stage1_11[163]},
      {stage2_11[73]}
   );
   gpc1_1 gpc2968 (
      {stage1_11[164]},
      {stage2_11[74]}
   );
   gpc1_1 gpc2969 (
      {stage1_11[165]},
      {stage2_11[75]}
   );
   gpc1_1 gpc2970 (
      {stage1_11[166]},
      {stage2_11[76]}
   );
   gpc1_1 gpc2971 (
      {stage1_11[167]},
      {stage2_11[77]}
   );
   gpc1_1 gpc2972 (
      {stage1_11[168]},
      {stage2_11[78]}
   );
   gpc1_1 gpc2973 (
      {stage1_11[169]},
      {stage2_11[79]}
   );
   gpc1_1 gpc2974 (
      {stage1_11[170]},
      {stage2_11[80]}
   );
   gpc1_1 gpc2975 (
      {stage1_11[171]},
      {stage2_11[81]}
   );
   gpc1_1 gpc2976 (
      {stage1_11[172]},
      {stage2_11[82]}
   );
   gpc1_1 gpc2977 (
      {stage1_11[173]},
      {stage2_11[83]}
   );
   gpc1_1 gpc2978 (
      {stage1_11[174]},
      {stage2_11[84]}
   );
   gpc1_1 gpc2979 (
      {stage1_11[175]},
      {stage2_11[85]}
   );
   gpc1_1 gpc2980 (
      {stage1_11[176]},
      {stage2_11[86]}
   );
   gpc1_1 gpc2981 (
      {stage1_11[177]},
      {stage2_11[87]}
   );
   gpc1_1 gpc2982 (
      {stage1_11[178]},
      {stage2_11[88]}
   );
   gpc1_1 gpc2983 (
      {stage1_11[179]},
      {stage2_11[89]}
   );
   gpc1_1 gpc2984 (
      {stage1_11[180]},
      {stage2_11[90]}
   );
   gpc1_1 gpc2985 (
      {stage1_11[181]},
      {stage2_11[91]}
   );
   gpc1_1 gpc2986 (
      {stage1_11[182]},
      {stage2_11[92]}
   );
   gpc1_1 gpc2987 (
      {stage1_11[183]},
      {stage2_11[93]}
   );
   gpc1_1 gpc2988 (
      {stage1_11[184]},
      {stage2_11[94]}
   );
   gpc1_1 gpc2989 (
      {stage1_11[185]},
      {stage2_11[95]}
   );
   gpc1_1 gpc2990 (
      {stage1_11[186]},
      {stage2_11[96]}
   );
   gpc1_1 gpc2991 (
      {stage1_11[187]},
      {stage2_11[97]}
   );
   gpc1_1 gpc2992 (
      {stage1_11[188]},
      {stage2_11[98]}
   );
   gpc1_1 gpc2993 (
      {stage1_11[189]},
      {stage2_11[99]}
   );
   gpc1_1 gpc2994 (
      {stage1_11[190]},
      {stage2_11[100]}
   );
   gpc1_1 gpc2995 (
      {stage1_11[191]},
      {stage2_11[101]}
   );
   gpc1_1 gpc2996 (
      {stage1_11[192]},
      {stage2_11[102]}
   );
   gpc1_1 gpc2997 (
      {stage1_11[193]},
      {stage2_11[103]}
   );
   gpc1_1 gpc2998 (
      {stage1_11[194]},
      {stage2_11[104]}
   );
   gpc1_1 gpc2999 (
      {stage1_11[195]},
      {stage2_11[105]}
   );
   gpc1_1 gpc3000 (
      {stage1_11[196]},
      {stage2_11[106]}
   );
   gpc1_1 gpc3001 (
      {stage1_11[197]},
      {stage2_11[107]}
   );
   gpc1_1 gpc3002 (
      {stage1_11[198]},
      {stage2_11[108]}
   );
   gpc1_1 gpc3003 (
      {stage1_11[199]},
      {stage2_11[109]}
   );
   gpc1_1 gpc3004 (
      {stage1_11[200]},
      {stage2_11[110]}
   );
   gpc1_1 gpc3005 (
      {stage1_11[201]},
      {stage2_11[111]}
   );
   gpc1_1 gpc3006 (
      {stage1_11[202]},
      {stage2_11[112]}
   );
   gpc1_1 gpc3007 (
      {stage1_11[203]},
      {stage2_11[113]}
   );
   gpc1_1 gpc3008 (
      {stage1_11[204]},
      {stage2_11[114]}
   );
   gpc1_1 gpc3009 (
      {stage1_11[205]},
      {stage2_11[115]}
   );
   gpc1_1 gpc3010 (
      {stage1_12[215]},
      {stage2_12[95]}
   );
   gpc1_1 gpc3011 (
      {stage1_12[216]},
      {stage2_12[96]}
   );
   gpc1_1 gpc3012 (
      {stage1_12[217]},
      {stage2_12[97]}
   );
   gpc1_1 gpc3013 (
      {stage1_12[218]},
      {stage2_12[98]}
   );
   gpc1_1 gpc3014 (
      {stage1_12[219]},
      {stage2_12[99]}
   );
   gpc1_1 gpc3015 (
      {stage1_12[220]},
      {stage2_12[100]}
   );
   gpc1_1 gpc3016 (
      {stage1_12[221]},
      {stage2_12[101]}
   );
   gpc1_1 gpc3017 (
      {stage1_13[198]},
      {stage2_13[90]}
   );
   gpc1_1 gpc3018 (
      {stage1_13[199]},
      {stage2_13[91]}
   );
   gpc1_1 gpc3019 (
      {stage1_13[200]},
      {stage2_13[92]}
   );
   gpc1_1 gpc3020 (
      {stage1_13[201]},
      {stage2_13[93]}
   );
   gpc1_1 gpc3021 (
      {stage1_13[202]},
      {stage2_13[94]}
   );
   gpc1_1 gpc3022 (
      {stage1_13[203]},
      {stage2_13[95]}
   );
   gpc1_1 gpc3023 (
      {stage1_13[204]},
      {stage2_13[96]}
   );
   gpc1_1 gpc3024 (
      {stage1_13[205]},
      {stage2_13[97]}
   );
   gpc1_1 gpc3025 (
      {stage1_13[206]},
      {stage2_13[98]}
   );
   gpc1_1 gpc3026 (
      {stage1_13[207]},
      {stage2_13[99]}
   );
   gpc1_1 gpc3027 (
      {stage1_13[208]},
      {stage2_13[100]}
   );
   gpc1_1 gpc3028 (
      {stage1_13[209]},
      {stage2_13[101]}
   );
   gpc1_1 gpc3029 (
      {stage1_13[210]},
      {stage2_13[102]}
   );
   gpc1_1 gpc3030 (
      {stage1_13[211]},
      {stage2_13[103]}
   );
   gpc1_1 gpc3031 (
      {stage1_13[212]},
      {stage2_13[104]}
   );
   gpc1_1 gpc3032 (
      {stage1_13[213]},
      {stage2_13[105]}
   );
   gpc1_1 gpc3033 (
      {stage1_13[214]},
      {stage2_13[106]}
   );
   gpc1_1 gpc3034 (
      {stage1_13[215]},
      {stage2_13[107]}
   );
   gpc1_1 gpc3035 (
      {stage1_13[216]},
      {stage2_13[108]}
   );
   gpc1_1 gpc3036 (
      {stage1_13[217]},
      {stage2_13[109]}
   );
   gpc1_1 gpc3037 (
      {stage1_13[218]},
      {stage2_13[110]}
   );
   gpc1_1 gpc3038 (
      {stage1_13[219]},
      {stage2_13[111]}
   );
   gpc1_1 gpc3039 (
      {stage1_13[220]},
      {stage2_13[112]}
   );
   gpc1_1 gpc3040 (
      {stage1_13[221]},
      {stage2_13[113]}
   );
   gpc1_1 gpc3041 (
      {stage1_13[222]},
      {stage2_13[114]}
   );
   gpc1_1 gpc3042 (
      {stage1_13[223]},
      {stage2_13[115]}
   );
   gpc1_1 gpc3043 (
      {stage1_13[224]},
      {stage2_13[116]}
   );
   gpc1_1 gpc3044 (
      {stage1_13[225]},
      {stage2_13[117]}
   );
   gpc1_1 gpc3045 (
      {stage1_13[226]},
      {stage2_13[118]}
   );
   gpc1_1 gpc3046 (
      {stage1_13[227]},
      {stage2_13[119]}
   );
   gpc1_1 gpc3047 (
      {stage1_13[228]},
      {stage2_13[120]}
   );
   gpc1_1 gpc3048 (
      {stage1_13[229]},
      {stage2_13[121]}
   );
   gpc1_1 gpc3049 (
      {stage1_13[230]},
      {stage2_13[122]}
   );
   gpc1_1 gpc3050 (
      {stage1_13[231]},
      {stage2_13[123]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[222]},
      {stage2_15[83]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[223]},
      {stage2_15[84]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[224]},
      {stage2_15[85]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[225]},
      {stage2_15[86]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[226]},
      {stage2_15[87]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[227]},
      {stage2_15[88]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[228]},
      {stage2_15[89]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[229]},
      {stage2_15[90]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[230]},
      {stage2_15[91]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[231]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[232]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[233]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[234]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[235]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[236]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[196]},
      {stage2_16[107]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[197]},
      {stage2_16[108]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[198]},
      {stage2_16[109]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[199]},
      {stage2_16[110]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[200]},
      {stage2_16[111]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[201]},
      {stage2_16[112]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[202]},
      {stage2_16[113]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[203]},
      {stage2_16[114]}
   );
   gpc1_1 gpc3074 (
      {stage1_16[204]},
      {stage2_16[115]}
   );
   gpc1_1 gpc3075 (
      {stage1_16[205]},
      {stage2_16[116]}
   );
   gpc1_1 gpc3076 (
      {stage1_16[206]},
      {stage2_16[117]}
   );
   gpc1_1 gpc3077 (
      {stage1_16[207]},
      {stage2_16[118]}
   );
   gpc1_1 gpc3078 (
      {stage1_16[208]},
      {stage2_16[119]}
   );
   gpc1_1 gpc3079 (
      {stage1_16[209]},
      {stage2_16[120]}
   );
   gpc1_1 gpc3080 (
      {stage1_16[210]},
      {stage2_16[121]}
   );
   gpc1_1 gpc3081 (
      {stage1_16[211]},
      {stage2_16[122]}
   );
   gpc1_1 gpc3082 (
      {stage1_16[212]},
      {stage2_16[123]}
   );
   gpc1_1 gpc3083 (
      {stage1_16[213]},
      {stage2_16[124]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[178]},
      {stage2_17[82]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[179]},
      {stage2_17[83]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[180]},
      {stage2_17[84]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[181]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[182]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[183]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[184]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[185]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[186]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[187]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[188]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[189]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[190]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[191]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[192]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[193]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[194]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[195]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[196]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[197]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[198]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[199]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[200]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[201]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[202]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[203]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[204]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3111 (
      {stage1_17[205]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3112 (
      {stage1_17[206]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3113 (
      {stage1_17[207]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3114 (
      {stage1_17[208]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3115 (
      {stage1_17[209]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3116 (
      {stage1_17[210]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3117 (
      {stage1_17[211]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3118 (
      {stage1_17[212]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3119 (
      {stage1_17[213]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3120 (
      {stage1_17[214]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3121 (
      {stage1_17[215]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3122 (
      {stage1_17[216]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3123 (
      {stage1_17[217]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3124 (
      {stage1_17[218]},
      {stage2_17[122]}
   );
   gpc1_1 gpc3125 (
      {stage1_17[219]},
      {stage2_17[123]}
   );
   gpc1_1 gpc3126 (
      {stage1_17[220]},
      {stage2_17[124]}
   );
   gpc1_1 gpc3127 (
      {stage1_17[221]},
      {stage2_17[125]}
   );
   gpc1_1 gpc3128 (
      {stage1_17[222]},
      {stage2_17[126]}
   );
   gpc1_1 gpc3129 (
      {stage1_17[223]},
      {stage2_17[127]}
   );
   gpc1_1 gpc3130 (
      {stage1_18[194]},
      {stage2_18[64]}
   );
   gpc1_1 gpc3131 (
      {stage1_18[195]},
      {stage2_18[65]}
   );
   gpc1_1 gpc3132 (
      {stage1_18[196]},
      {stage2_18[66]}
   );
   gpc1_1 gpc3133 (
      {stage1_18[197]},
      {stage2_18[67]}
   );
   gpc1_1 gpc3134 (
      {stage1_18[198]},
      {stage2_18[68]}
   );
   gpc1_1 gpc3135 (
      {stage1_18[199]},
      {stage2_18[69]}
   );
   gpc1_1 gpc3136 (
      {stage1_18[200]},
      {stage2_18[70]}
   );
   gpc1_1 gpc3137 (
      {stage1_18[201]},
      {stage2_18[71]}
   );
   gpc1_1 gpc3138 (
      {stage1_18[202]},
      {stage2_18[72]}
   );
   gpc1_1 gpc3139 (
      {stage1_19[261]},
      {stage2_19[96]}
   );
   gpc1_1 gpc3140 (
      {stage1_19[262]},
      {stage2_19[97]}
   );
   gpc1_1 gpc3141 (
      {stage1_20[211]},
      {stage2_20[107]}
   );
   gpc1_1 gpc3142 (
      {stage1_20[212]},
      {stage2_20[108]}
   );
   gpc1_1 gpc3143 (
      {stage1_20[213]},
      {stage2_20[109]}
   );
   gpc1_1 gpc3144 (
      {stage1_21[227]},
      {stage2_21[82]}
   );
   gpc1_1 gpc3145 (
      {stage1_21[228]},
      {stage2_21[83]}
   );
   gpc1_1 gpc3146 (
      {stage1_21[229]},
      {stage2_21[84]}
   );
   gpc1_1 gpc3147 (
      {stage1_21[230]},
      {stage2_21[85]}
   );
   gpc1_1 gpc3148 (
      {stage1_21[231]},
      {stage2_21[86]}
   );
   gpc1_1 gpc3149 (
      {stage1_21[232]},
      {stage2_21[87]}
   );
   gpc1_1 gpc3150 (
      {stage1_21[233]},
      {stage2_21[88]}
   );
   gpc1_1 gpc3151 (
      {stage1_21[234]},
      {stage2_21[89]}
   );
   gpc1_1 gpc3152 (
      {stage1_21[235]},
      {stage2_21[90]}
   );
   gpc1_1 gpc3153 (
      {stage1_21[236]},
      {stage2_21[91]}
   );
   gpc1_1 gpc3154 (
      {stage1_21[237]},
      {stage2_21[92]}
   );
   gpc1_1 gpc3155 (
      {stage1_21[238]},
      {stage2_21[93]}
   );
   gpc1_1 gpc3156 (
      {stage1_21[239]},
      {stage2_21[94]}
   );
   gpc1_1 gpc3157 (
      {stage1_21[240]},
      {stage2_21[95]}
   );
   gpc1_1 gpc3158 (
      {stage1_21[241]},
      {stage2_21[96]}
   );
   gpc1_1 gpc3159 (
      {stage1_21[242]},
      {stage2_21[97]}
   );
   gpc1_1 gpc3160 (
      {stage1_21[243]},
      {stage2_21[98]}
   );
   gpc1_1 gpc3161 (
      {stage1_21[244]},
      {stage2_21[99]}
   );
   gpc1_1 gpc3162 (
      {stage1_21[245]},
      {stage2_21[100]}
   );
   gpc1_1 gpc3163 (
      {stage1_21[246]},
      {stage2_21[101]}
   );
   gpc1_1 gpc3164 (
      {stage1_21[247]},
      {stage2_21[102]}
   );
   gpc1_1 gpc3165 (
      {stage1_21[248]},
      {stage2_21[103]}
   );
   gpc1_1 gpc3166 (
      {stage1_21[249]},
      {stage2_21[104]}
   );
   gpc1_1 gpc3167 (
      {stage1_21[250]},
      {stage2_21[105]}
   );
   gpc1_1 gpc3168 (
      {stage1_21[251]},
      {stage2_21[106]}
   );
   gpc1_1 gpc3169 (
      {stage1_21[252]},
      {stage2_21[107]}
   );
   gpc1_1 gpc3170 (
      {stage1_21[253]},
      {stage2_21[108]}
   );
   gpc1_1 gpc3171 (
      {stage1_21[254]},
      {stage2_21[109]}
   );
   gpc1_1 gpc3172 (
      {stage1_21[255]},
      {stage2_21[110]}
   );
   gpc1_1 gpc3173 (
      {stage1_21[256]},
      {stage2_21[111]}
   );
   gpc1_1 gpc3174 (
      {stage1_21[257]},
      {stage2_21[112]}
   );
   gpc1_1 gpc3175 (
      {stage1_21[258]},
      {stage2_21[113]}
   );
   gpc1_1 gpc3176 (
      {stage1_21[259]},
      {stage2_21[114]}
   );
   gpc1_1 gpc3177 (
      {stage1_21[260]},
      {stage2_21[115]}
   );
   gpc1_1 gpc3178 (
      {stage1_21[261]},
      {stage2_21[116]}
   );
   gpc1_1 gpc3179 (
      {stage1_21[262]},
      {stage2_21[117]}
   );
   gpc1_1 gpc3180 (
      {stage1_21[263]},
      {stage2_21[118]}
   );
   gpc1_1 gpc3181 (
      {stage1_21[264]},
      {stage2_21[119]}
   );
   gpc1_1 gpc3182 (
      {stage1_21[265]},
      {stage2_21[120]}
   );
   gpc1_1 gpc3183 (
      {stage1_21[266]},
      {stage2_21[121]}
   );
   gpc1_1 gpc3184 (
      {stage1_21[267]},
      {stage2_21[122]}
   );
   gpc1_1 gpc3185 (
      {stage1_21[268]},
      {stage2_21[123]}
   );
   gpc1_1 gpc3186 (
      {stage1_21[269]},
      {stage2_21[124]}
   );
   gpc1_1 gpc3187 (
      {stage1_22[268]},
      {stage2_22[89]}
   );
   gpc1_1 gpc3188 (
      {stage1_22[269]},
      {stage2_22[90]}
   );
   gpc1_1 gpc3189 (
      {stage1_22[270]},
      {stage2_22[91]}
   );
   gpc1_1 gpc3190 (
      {stage1_22[271]},
      {stage2_22[92]}
   );
   gpc1_1 gpc3191 (
      {stage1_22[272]},
      {stage2_22[93]}
   );
   gpc1_1 gpc3192 (
      {stage1_22[273]},
      {stage2_22[94]}
   );
   gpc1_1 gpc3193 (
      {stage1_23[146]},
      {stage2_23[103]}
   );
   gpc1_1 gpc3194 (
      {stage1_23[147]},
      {stage2_23[104]}
   );
   gpc1_1 gpc3195 (
      {stage1_23[148]},
      {stage2_23[105]}
   );
   gpc1_1 gpc3196 (
      {stage1_23[149]},
      {stage2_23[106]}
   );
   gpc1_1 gpc3197 (
      {stage1_23[150]},
      {stage2_23[107]}
   );
   gpc1_1 gpc3198 (
      {stage1_23[151]},
      {stage2_23[108]}
   );
   gpc1_1 gpc3199 (
      {stage1_23[152]},
      {stage2_23[109]}
   );
   gpc1_1 gpc3200 (
      {stage1_23[153]},
      {stage2_23[110]}
   );
   gpc1_1 gpc3201 (
      {stage1_23[154]},
      {stage2_23[111]}
   );
   gpc1_1 gpc3202 (
      {stage1_23[155]},
      {stage2_23[112]}
   );
   gpc1_1 gpc3203 (
      {stage1_23[156]},
      {stage2_23[113]}
   );
   gpc1_1 gpc3204 (
      {stage1_23[157]},
      {stage2_23[114]}
   );
   gpc1_1 gpc3205 (
      {stage1_23[158]},
      {stage2_23[115]}
   );
   gpc1_1 gpc3206 (
      {stage1_23[159]},
      {stage2_23[116]}
   );
   gpc1_1 gpc3207 (
      {stage1_23[160]},
      {stage2_23[117]}
   );
   gpc1_1 gpc3208 (
      {stage1_23[161]},
      {stage2_23[118]}
   );
   gpc1_1 gpc3209 (
      {stage1_23[162]},
      {stage2_23[119]}
   );
   gpc1_1 gpc3210 (
      {stage1_23[163]},
      {stage2_23[120]}
   );
   gpc1_1 gpc3211 (
      {stage1_23[164]},
      {stage2_23[121]}
   );
   gpc1_1 gpc3212 (
      {stage1_23[165]},
      {stage2_23[122]}
   );
   gpc1_1 gpc3213 (
      {stage1_24[217]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3214 (
      {stage1_24[218]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3215 (
      {stage1_24[219]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3216 (
      {stage1_24[220]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3217 (
      {stage1_25[255]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3218 (
      {stage1_25[256]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3219 (
      {stage1_25[257]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3220 (
      {stage1_25[258]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3221 (
      {stage1_25[259]},
      {stage2_25[88]}
   );
   gpc1_1 gpc3222 (
      {stage1_25[260]},
      {stage2_25[89]}
   );
   gpc1_1 gpc3223 (
      {stage1_25[261]},
      {stage2_25[90]}
   );
   gpc1_1 gpc3224 (
      {stage1_25[262]},
      {stage2_25[91]}
   );
   gpc1_1 gpc3225 (
      {stage1_25[263]},
      {stage2_25[92]}
   );
   gpc1_1 gpc3226 (
      {stage1_25[264]},
      {stage2_25[93]}
   );
   gpc1_1 gpc3227 (
      {stage1_25[265]},
      {stage2_25[94]}
   );
   gpc1_1 gpc3228 (
      {stage1_25[266]},
      {stage2_25[95]}
   );
   gpc1_1 gpc3229 (
      {stage1_25[267]},
      {stage2_25[96]}
   );
   gpc1_1 gpc3230 (
      {stage1_25[268]},
      {stage2_25[97]}
   );
   gpc1_1 gpc3231 (
      {stage1_25[269]},
      {stage2_25[98]}
   );
   gpc1_1 gpc3232 (
      {stage1_25[270]},
      {stage2_25[99]}
   );
   gpc1_1 gpc3233 (
      {stage1_25[271]},
      {stage2_25[100]}
   );
   gpc1_1 gpc3234 (
      {stage1_25[272]},
      {stage2_25[101]}
   );
   gpc1_1 gpc3235 (
      {stage1_25[273]},
      {stage2_25[102]}
   );
   gpc1_1 gpc3236 (
      {stage1_26[186]},
      {stage2_26[95]}
   );
   gpc1_1 gpc3237 (
      {stage1_26[187]},
      {stage2_26[96]}
   );
   gpc1_1 gpc3238 (
      {stage1_26[188]},
      {stage2_26[97]}
   );
   gpc1_1 gpc3239 (
      {stage1_26[189]},
      {stage2_26[98]}
   );
   gpc1_1 gpc3240 (
      {stage1_26[190]},
      {stage2_26[99]}
   );
   gpc1_1 gpc3241 (
      {stage1_27[196]},
      {stage2_27[81]}
   );
   gpc1_1 gpc3242 (
      {stage1_27[197]},
      {stage2_27[82]}
   );
   gpc1_1 gpc3243 (
      {stage1_27[198]},
      {stage2_27[83]}
   );
   gpc1_1 gpc3244 (
      {stage1_27[199]},
      {stage2_27[84]}
   );
   gpc1_1 gpc3245 (
      {stage1_28[149]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3246 (
      {stage1_28[150]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3247 (
      {stage1_28[151]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3248 (
      {stage1_28[152]},
      {stage2_28[75]}
   );
   gpc1_1 gpc3249 (
      {stage1_28[153]},
      {stage2_28[76]}
   );
   gpc1_1 gpc3250 (
      {stage1_28[154]},
      {stage2_28[77]}
   );
   gpc1_1 gpc3251 (
      {stage1_28[155]},
      {stage2_28[78]}
   );
   gpc1_1 gpc3252 (
      {stage1_28[156]},
      {stage2_28[79]}
   );
   gpc1_1 gpc3253 (
      {stage1_28[157]},
      {stage2_28[80]}
   );
   gpc1_1 gpc3254 (
      {stage1_28[158]},
      {stage2_28[81]}
   );
   gpc1_1 gpc3255 (
      {stage1_28[159]},
      {stage2_28[82]}
   );
   gpc1_1 gpc3256 (
      {stage1_28[160]},
      {stage2_28[83]}
   );
   gpc1_1 gpc3257 (
      {stage1_28[161]},
      {stage2_28[84]}
   );
   gpc1_1 gpc3258 (
      {stage1_28[162]},
      {stage2_28[85]}
   );
   gpc1_1 gpc3259 (
      {stage1_28[163]},
      {stage2_28[86]}
   );
   gpc1_1 gpc3260 (
      {stage1_28[164]},
      {stage2_28[87]}
   );
   gpc1_1 gpc3261 (
      {stage1_28[165]},
      {stage2_28[88]}
   );
   gpc1_1 gpc3262 (
      {stage1_28[166]},
      {stage2_28[89]}
   );
   gpc1_1 gpc3263 (
      {stage1_28[167]},
      {stage2_28[90]}
   );
   gpc1_1 gpc3264 (
      {stage1_28[168]},
      {stage2_28[91]}
   );
   gpc1_1 gpc3265 (
      {stage1_28[169]},
      {stage2_28[92]}
   );
   gpc1_1 gpc3266 (
      {stage1_28[170]},
      {stage2_28[93]}
   );
   gpc1_1 gpc3267 (
      {stage1_28[171]},
      {stage2_28[94]}
   );
   gpc1_1 gpc3268 (
      {stage1_28[172]},
      {stage2_28[95]}
   );
   gpc1_1 gpc3269 (
      {stage1_28[173]},
      {stage2_28[96]}
   );
   gpc1_1 gpc3270 (
      {stage1_28[174]},
      {stage2_28[97]}
   );
   gpc1_1 gpc3271 (
      {stage1_28[175]},
      {stage2_28[98]}
   );
   gpc1_1 gpc3272 (
      {stage1_28[176]},
      {stage2_28[99]}
   );
   gpc1_1 gpc3273 (
      {stage1_28[177]},
      {stage2_28[100]}
   );
   gpc1_1 gpc3274 (
      {stage1_28[178]},
      {stage2_28[101]}
   );
   gpc1_1 gpc3275 (
      {stage1_28[179]},
      {stage2_28[102]}
   );
   gpc1_1 gpc3276 (
      {stage1_28[180]},
      {stage2_28[103]}
   );
   gpc1_1 gpc3277 (
      {stage1_28[181]},
      {stage2_28[104]}
   );
   gpc1_1 gpc3278 (
      {stage1_28[182]},
      {stage2_28[105]}
   );
   gpc1_1 gpc3279 (
      {stage1_28[183]},
      {stage2_28[106]}
   );
   gpc1_1 gpc3280 (
      {stage1_28[184]},
      {stage2_28[107]}
   );
   gpc1_1 gpc3281 (
      {stage1_28[185]},
      {stage2_28[108]}
   );
   gpc1_1 gpc3282 (
      {stage1_28[186]},
      {stage2_28[109]}
   );
   gpc1_1 gpc3283 (
      {stage1_28[187]},
      {stage2_28[110]}
   );
   gpc1_1 gpc3284 (
      {stage1_28[188]},
      {stage2_28[111]}
   );
   gpc1_1 gpc3285 (
      {stage1_28[189]},
      {stage2_28[112]}
   );
   gpc1_1 gpc3286 (
      {stage1_28[190]},
      {stage2_28[113]}
   );
   gpc1_1 gpc3287 (
      {stage1_28[191]},
      {stage2_28[114]}
   );
   gpc1_1 gpc3288 (
      {stage1_28[192]},
      {stage2_28[115]}
   );
   gpc1_1 gpc3289 (
      {stage1_28[193]},
      {stage2_28[116]}
   );
   gpc1_1 gpc3290 (
      {stage1_28[194]},
      {stage2_28[117]}
   );
   gpc1_1 gpc3291 (
      {stage1_28[195]},
      {stage2_28[118]}
   );
   gpc1_1 gpc3292 (
      {stage1_28[196]},
      {stage2_28[119]}
   );
   gpc1_1 gpc3293 (
      {stage1_28[197]},
      {stage2_28[120]}
   );
   gpc1_1 gpc3294 (
      {stage1_28[198]},
      {stage2_28[121]}
   );
   gpc1_1 gpc3295 (
      {stage1_28[199]},
      {stage2_28[122]}
   );
   gpc1_1 gpc3296 (
      {stage1_28[200]},
      {stage2_28[123]}
   );
   gpc1_1 gpc3297 (
      {stage1_28[201]},
      {stage2_28[124]}
   );
   gpc1_1 gpc3298 (
      {stage1_28[202]},
      {stage2_28[125]}
   );
   gpc1_1 gpc3299 (
      {stage1_28[203]},
      {stage2_28[126]}
   );
   gpc1_1 gpc3300 (
      {stage1_28[204]},
      {stage2_28[127]}
   );
   gpc1_1 gpc3301 (
      {stage1_28[205]},
      {stage2_28[128]}
   );
   gpc1_1 gpc3302 (
      {stage1_28[206]},
      {stage2_28[129]}
   );
   gpc1_1 gpc3303 (
      {stage1_28[207]},
      {stage2_28[130]}
   );
   gpc1_1 gpc3304 (
      {stage1_28[208]},
      {stage2_28[131]}
   );
   gpc1_1 gpc3305 (
      {stage1_28[209]},
      {stage2_28[132]}
   );
   gpc1_1 gpc3306 (
      {stage1_28[210]},
      {stage2_28[133]}
   );
   gpc1_1 gpc3307 (
      {stage1_28[211]},
      {stage2_28[134]}
   );
   gpc1_1 gpc3308 (
      {stage1_28[212]},
      {stage2_28[135]}
   );
   gpc1_1 gpc3309 (
      {stage1_28[213]},
      {stage2_28[136]}
   );
   gpc1_1 gpc3310 (
      {stage1_28[214]},
      {stage2_28[137]}
   );
   gpc1_1 gpc3311 (
      {stage1_28[215]},
      {stage2_28[138]}
   );
   gpc1_1 gpc3312 (
      {stage1_28[216]},
      {stage2_28[139]}
   );
   gpc1_1 gpc3313 (
      {stage1_28[217]},
      {stage2_28[140]}
   );
   gpc1_1 gpc3314 (
      {stage1_28[218]},
      {stage2_28[141]}
   );
   gpc1_1 gpc3315 (
      {stage1_28[219]},
      {stage2_28[142]}
   );
   gpc1_1 gpc3316 (
      {stage1_28[220]},
      {stage2_28[143]}
   );
   gpc1_1 gpc3317 (
      {stage1_28[221]},
      {stage2_28[144]}
   );
   gpc1_1 gpc3318 (
      {stage1_28[222]},
      {stage2_28[145]}
   );
   gpc1_1 gpc3319 (
      {stage1_28[223]},
      {stage2_28[146]}
   );
   gpc1_1 gpc3320 (
      {stage1_28[224]},
      {stage2_28[147]}
   );
   gpc1_1 gpc3321 (
      {stage1_28[225]},
      {stage2_28[148]}
   );
   gpc1_1 gpc3322 (
      {stage1_28[226]},
      {stage2_28[149]}
   );
   gpc1_1 gpc3323 (
      {stage1_28[227]},
      {stage2_28[150]}
   );
   gpc1_1 gpc3324 (
      {stage1_28[228]},
      {stage2_28[151]}
   );
   gpc1_1 gpc3325 (
      {stage1_28[229]},
      {stage2_28[152]}
   );
   gpc1_1 gpc3326 (
      {stage1_28[230]},
      {stage2_28[153]}
   );
   gpc1_1 gpc3327 (
      {stage1_28[231]},
      {stage2_28[154]}
   );
   gpc1_1 gpc3328 (
      {stage1_28[232]},
      {stage2_28[155]}
   );
   gpc1_1 gpc3329 (
      {stage1_28[233]},
      {stage2_28[156]}
   );
   gpc1_1 gpc3330 (
      {stage1_28[234]},
      {stage2_28[157]}
   );
   gpc1_1 gpc3331 (
      {stage1_28[235]},
      {stage2_28[158]}
   );
   gpc1_1 gpc3332 (
      {stage1_28[236]},
      {stage2_28[159]}
   );
   gpc1_1 gpc3333 (
      {stage1_28[237]},
      {stage2_28[160]}
   );
   gpc1_1 gpc3334 (
      {stage1_28[238]},
      {stage2_28[161]}
   );
   gpc1_1 gpc3335 (
      {stage1_28[239]},
      {stage2_28[162]}
   );
   gpc1_1 gpc3336 (
      {stage1_28[240]},
      {stage2_28[163]}
   );
   gpc1_1 gpc3337 (
      {stage1_28[241]},
      {stage2_28[164]}
   );
   gpc1_1 gpc3338 (
      {stage1_28[242]},
      {stage2_28[165]}
   );
   gpc1_1 gpc3339 (
      {stage1_28[243]},
      {stage2_28[166]}
   );
   gpc1_1 gpc3340 (
      {stage1_28[244]},
      {stage2_28[167]}
   );
   gpc1_1 gpc3341 (
      {stage1_28[245]},
      {stage2_28[168]}
   );
   gpc1_1 gpc3342 (
      {stage1_28[246]},
      {stage2_28[169]}
   );
   gpc1_1 gpc3343 (
      {stage1_28[247]},
      {stage2_28[170]}
   );
   gpc1_1 gpc3344 (
      {stage1_29[180]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3345 (
      {stage1_29[181]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3346 (
      {stage1_29[182]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3347 (
      {stage1_29[183]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3348 (
      {stage1_29[184]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3349 (
      {stage1_29[185]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3350 (
      {stage1_29[186]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3351 (
      {stage1_29[187]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3352 (
      {stage1_29[188]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3353 (
      {stage1_29[189]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3354 (
      {stage1_29[190]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3355 (
      {stage1_29[191]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3356 (
      {stage1_29[192]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3357 (
      {stage1_29[193]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3358 (
      {stage1_29[194]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3359 (
      {stage1_29[195]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3360 (
      {stage1_29[196]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3361 (
      {stage1_29[197]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3362 (
      {stage1_29[198]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3363 (
      {stage1_29[199]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3364 (
      {stage1_29[200]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3365 (
      {stage1_29[201]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3366 (
      {stage1_29[202]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3367 (
      {stage1_29[203]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3368 (
      {stage1_29[204]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3369 (
      {stage1_29[205]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3370 (
      {stage1_29[206]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3371 (
      {stage1_29[207]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3372 (
      {stage1_29[208]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3373 (
      {stage1_29[209]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3374 (
      {stage1_29[210]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3375 (
      {stage1_29[211]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3376 (
      {stage1_29[212]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3377 (
      {stage1_29[213]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3378 (
      {stage1_29[214]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3379 (
      {stage1_29[215]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3380 (
      {stage1_29[216]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3381 (
      {stage1_29[217]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3382 (
      {stage1_29[218]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3383 (
      {stage1_29[219]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3384 (
      {stage1_29[220]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3385 (
      {stage1_29[221]},
      {stage2_29[121]}
   );
   gpc1_1 gpc3386 (
      {stage1_29[222]},
      {stage2_29[122]}
   );
   gpc1_1 gpc3387 (
      {stage1_29[223]},
      {stage2_29[123]}
   );
   gpc1_1 gpc3388 (
      {stage1_29[224]},
      {stage2_29[124]}
   );
   gpc1_1 gpc3389 (
      {stage1_29[225]},
      {stage2_29[125]}
   );
   gpc1_1 gpc3390 (
      {stage1_29[226]},
      {stage2_29[126]}
   );
   gpc1_1 gpc3391 (
      {stage1_29[227]},
      {stage2_29[127]}
   );
   gpc1_1 gpc3392 (
      {stage1_29[228]},
      {stage2_29[128]}
   );
   gpc1_1 gpc3393 (
      {stage1_29[229]},
      {stage2_29[129]}
   );
   gpc1_1 gpc3394 (
      {stage1_29[230]},
      {stage2_29[130]}
   );
   gpc1_1 gpc3395 (
      {stage1_29[231]},
      {stage2_29[131]}
   );
   gpc1_1 gpc3396 (
      {stage1_29[232]},
      {stage2_29[132]}
   );
   gpc1_1 gpc3397 (
      {stage1_29[233]},
      {stage2_29[133]}
   );
   gpc1_1 gpc3398 (
      {stage1_29[234]},
      {stage2_29[134]}
   );
   gpc1_1 gpc3399 (
      {stage1_29[235]},
      {stage2_29[135]}
   );
   gpc1_1 gpc3400 (
      {stage1_29[236]},
      {stage2_29[136]}
   );
   gpc1_1 gpc3401 (
      {stage1_29[237]},
      {stage2_29[137]}
   );
   gpc1_1 gpc3402 (
      {stage1_29[238]},
      {stage2_29[138]}
   );
   gpc1_1 gpc3403 (
      {stage1_29[239]},
      {stage2_29[139]}
   );
   gpc1_1 gpc3404 (
      {stage1_29[240]},
      {stage2_29[140]}
   );
   gpc1_1 gpc3405 (
      {stage1_29[241]},
      {stage2_29[141]}
   );
   gpc1_1 gpc3406 (
      {stage1_29[242]},
      {stage2_29[142]}
   );
   gpc1_1 gpc3407 (
      {stage1_30[192]},
      {stage2_30[77]}
   );
   gpc1_1 gpc3408 (
      {stage1_30[193]},
      {stage2_30[78]}
   );
   gpc1_1 gpc3409 (
      {stage1_30[194]},
      {stage2_30[79]}
   );
   gpc1_1 gpc3410 (
      {stage1_30[195]},
      {stage2_30[80]}
   );
   gpc1_1 gpc3411 (
      {stage1_30[196]},
      {stage2_30[81]}
   );
   gpc1_1 gpc3412 (
      {stage1_30[197]},
      {stage2_30[82]}
   );
   gpc1_1 gpc3413 (
      {stage1_30[198]},
      {stage2_30[83]}
   );
   gpc1_1 gpc3414 (
      {stage1_30[199]},
      {stage2_30[84]}
   );
   gpc1_1 gpc3415 (
      {stage1_30[200]},
      {stage2_30[85]}
   );
   gpc1_1 gpc3416 (
      {stage1_30[201]},
      {stage2_30[86]}
   );
   gpc1_1 gpc3417 (
      {stage1_30[202]},
      {stage2_30[87]}
   );
   gpc1_1 gpc3418 (
      {stage1_30[203]},
      {stage2_30[88]}
   );
   gpc1_1 gpc3419 (
      {stage1_30[204]},
      {stage2_30[89]}
   );
   gpc1_1 gpc3420 (
      {stage1_30[205]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3421 (
      {stage1_30[206]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3422 (
      {stage1_31[215]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3423 (
      {stage1_31[216]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3424 (
      {stage1_31[217]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3425 (
      {stage1_31[218]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3426 (
      {stage1_31[219]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3427 (
      {stage1_31[220]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3428 (
      {stage1_31[221]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3429 (
      {stage1_31[222]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3430 (
      {stage1_31[223]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3431 (
      {stage1_31[224]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3432 (
      {stage1_31[225]},
      {stage2_31[84]}
   );
   gpc1_1 gpc3433 (
      {stage1_31[226]},
      {stage2_31[85]}
   );
   gpc1_1 gpc3434 (
      {stage1_31[227]},
      {stage2_31[86]}
   );
   gpc1_1 gpc3435 (
      {stage1_31[228]},
      {stage2_31[87]}
   );
   gpc1_1 gpc3436 (
      {stage1_31[229]},
      {stage2_31[88]}
   );
   gpc1_1 gpc3437 (
      {stage1_31[230]},
      {stage2_31[89]}
   );
   gpc1_1 gpc3438 (
      {stage1_31[231]},
      {stage2_31[90]}
   );
   gpc1_1 gpc3439 (
      {stage1_31[232]},
      {stage2_31[91]}
   );
   gpc1_1 gpc3440 (
      {stage1_31[233]},
      {stage2_31[92]}
   );
   gpc1_1 gpc3441 (
      {stage1_31[234]},
      {stage2_31[93]}
   );
   gpc1_1 gpc3442 (
      {stage1_31[235]},
      {stage2_31[94]}
   );
   gpc1_1 gpc3443 (
      {stage1_31[236]},
      {stage2_31[95]}
   );
   gpc1_1 gpc3444 (
      {stage1_31[237]},
      {stage2_31[96]}
   );
   gpc1_1 gpc3445 (
      {stage1_31[238]},
      {stage2_31[97]}
   );
   gpc1_1 gpc3446 (
      {stage1_31[239]},
      {stage2_31[98]}
   );
   gpc1_1 gpc3447 (
      {stage1_31[240]},
      {stage2_31[99]}
   );
   gpc1_1 gpc3448 (
      {stage1_31[241]},
      {stage2_31[100]}
   );
   gpc1_1 gpc3449 (
      {stage1_31[242]},
      {stage2_31[101]}
   );
   gpc1_1 gpc3450 (
      {stage1_32[145]},
      {stage2_32[69]}
   );
   gpc1_1 gpc3451 (
      {stage1_32[146]},
      {stage2_32[70]}
   );
   gpc1_1 gpc3452 (
      {stage1_32[147]},
      {stage2_32[71]}
   );
   gpc1_1 gpc3453 (
      {stage1_32[148]},
      {stage2_32[72]}
   );
   gpc1_1 gpc3454 (
      {stage1_32[149]},
      {stage2_32[73]}
   );
   gpc1163_5 gpc3455 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3456 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc3457 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc3458 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc3459 (
      {stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24], stage2_0[25], stage2_0[26]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc3460 (
      {stage2_0[27], stage2_0[28], stage2_0[29], stage2_0[30], stage2_0[31], stage2_0[32]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc3461 (
      {stage2_0[33], stage2_0[34], stage2_0[35], stage2_0[36], stage2_0[37], stage2_0[38]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3462 (
      {stage2_0[39], stage2_0[40], stage2_0[41], stage2_0[42], stage2_0[43], stage2_0[44]},
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7],stage3_0[7]}
   );
   gpc606_5 gpc3463 (
      {stage2_0[45], stage2_0[46], stage2_0[47], stage2_0[48], stage2_0[49], stage2_0[50]},
      {stage2_2[43], stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8],stage3_0[8]}
   );
   gpc606_5 gpc3464 (
      {stage2_0[51], stage2_0[52], stage2_0[53], stage2_0[54], stage2_0[55], stage2_0[56]},
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9],stage3_0[9]}
   );
   gpc606_5 gpc3465 (
      {stage2_0[57], stage2_0[58], stage2_0[59], stage2_0[60], stage2_0[61], stage2_0[62]},
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60]},
      {stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10],stage3_0[10]}
   );
   gpc606_5 gpc3466 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3467 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3468 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3469 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3470 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3471 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3472 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[6],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc615_5 gpc3473 (
      {stage2_2[61], stage2_2[62], stage2_2[63], stage2_2[64], stage2_2[65]},
      {stage2_3[43]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[7],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc3474 (
      {stage2_2[66], stage2_2[67], stage2_2[68], stage2_2[69], stage2_2[70]},
      {stage2_3[44]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[8],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc615_5 gpc3475 (
      {stage2_2[71], stage2_2[72], stage2_2[73], stage2_2[74], stage2_2[75]},
      {stage2_3[45]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[9],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc615_5 gpc3476 (
      {stage2_2[76], stage2_2[77], stage2_2[78], stage2_2[79], stage2_2[80]},
      {stage2_3[46]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[10],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc615_5 gpc3477 (
      {stage2_3[47], stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[11],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc3478 (
      {stage2_3[52], stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[12],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc3479 (
      {stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[13],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3480 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage2_4[27]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[7],stage3_5[14],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3481 (
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71]},
      {stage2_4[28]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[8],stage3_5[15],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc3482 (
      {stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76]},
      {stage2_4[29]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[9],stage3_5[16],stage3_4[27],stage3_3[27]}
   );
   gpc606_5 gpc3483 (
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[6],stage3_6[10],stage3_5[17],stage3_4[28]}
   );
   gpc606_5 gpc3484 (
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[7],stage3_6[11],stage3_5[18],stage3_4[29]}
   );
   gpc606_5 gpc3485 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46], stage2_4[47]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[8],stage3_6[12],stage3_5[19],stage3_4[30]}
   );
   gpc606_5 gpc3486 (
      {stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[9],stage3_6[13],stage3_5[20],stage3_4[31]}
   );
   gpc606_5 gpc3487 (
      {stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[10],stage3_6[14],stage3_5[21],stage3_4[32]}
   );
   gpc606_5 gpc3488 (
      {stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[11],stage3_6[15],stage3_5[22],stage3_4[33]}
   );
   gpc606_5 gpc3489 (
      {stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[12],stage3_6[16],stage3_5[23],stage3_4[34]}
   );
   gpc606_5 gpc3490 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[13],stage3_6[17],stage3_5[24],stage3_4[35]}
   );
   gpc606_5 gpc3491 (
      {stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[14],stage3_6[18],stage3_5[25],stage3_4[36]}
   );
   gpc606_5 gpc3492 (
      {stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88], stage2_4[89]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[15],stage3_6[19],stage3_5[26],stage3_4[37]}
   );
   gpc606_5 gpc3493 (
      {stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94], stage2_4[95]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[16],stage3_6[20],stage3_5[27],stage3_4[38]}
   );
   gpc606_5 gpc3494 (
      {stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100], stage2_4[101]},
      {stage2_6[66], stage2_6[67], stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71]},
      {stage3_8[11],stage3_7[17],stage3_6[21],stage3_5[28],stage3_4[39]}
   );
   gpc606_5 gpc3495 (
      {stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106], stage2_4[107]},
      {stage2_6[72], stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage3_8[12],stage3_7[18],stage3_6[22],stage3_5[29],stage3_4[40]}
   );
   gpc606_5 gpc3496 (
      {stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111], stage2_4[112], stage2_4[113]},
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage3_8[13],stage3_7[19],stage3_6[23],stage3_5[30],stage3_4[41]}
   );
   gpc606_5 gpc3497 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[14],stage3_7[20],stage3_6[24],stage3_5[31]}
   );
   gpc606_5 gpc3498 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[15],stage3_7[21],stage3_6[25],stage3_5[32]}
   );
   gpc606_5 gpc3499 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[16],stage3_7[22],stage3_6[26],stage3_5[33]}
   );
   gpc606_5 gpc3500 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[17],stage3_7[23],stage3_6[27],stage3_5[34]}
   );
   gpc606_5 gpc3501 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[18],stage3_7[24],stage3_6[28],stage3_5[35]}
   );
   gpc606_5 gpc3502 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[19],stage3_7[25],stage3_6[29],stage3_5[36]}
   );
   gpc615_5 gpc3503 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[36]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[6],stage3_8[20],stage3_7[26],stage3_6[30]}
   );
   gpc615_5 gpc3504 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[7],stage3_8[21],stage3_7[27]}
   );
   gpc615_5 gpc3505 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[8],stage3_8[22],stage3_7[28]}
   );
   gpc615_5 gpc3506 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[9],stage3_8[23],stage3_7[29]}
   );
   gpc615_5 gpc3507 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[10],stage3_8[24],stage3_7[30]}
   );
   gpc615_5 gpc3508 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[10]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[5],stage3_9[11],stage3_8[25],stage3_7[31]}
   );
   gpc615_5 gpc3509 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[11]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[6],stage3_9[12],stage3_8[26],stage3_7[32]}
   );
   gpc615_5 gpc3510 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[12]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[7],stage3_9[13],stage3_8[27],stage3_7[33]}
   );
   gpc615_5 gpc3511 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[13]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[8],stage3_9[14],stage3_8[28],stage3_7[34]}
   );
   gpc615_5 gpc3512 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[14]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[9],stage3_9[15],stage3_8[29],stage3_7[35]}
   );
   gpc615_5 gpc3513 (
      {stage2_7[82], stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86]},
      {stage2_8[15]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[10],stage3_9[16],stage3_8[30],stage3_7[36]}
   );
   gpc615_5 gpc3514 (
      {stage2_7[87], stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91]},
      {stage2_8[16]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[11],stage3_9[17],stage3_8[31],stage3_7[37]}
   );
   gpc615_5 gpc3515 (
      {stage2_7[92], stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96]},
      {stage2_8[17]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[12],stage3_9[18],stage3_8[32],stage3_7[38]}
   );
   gpc615_5 gpc3516 (
      {stage2_7[97], stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101]},
      {stage2_8[18]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[13],stage3_9[19],stage3_8[33],stage3_7[39]}
   );
   gpc606_5 gpc3517 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[13],stage3_10[14],stage3_9[20],stage3_8[34]}
   );
   gpc606_5 gpc3518 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[14],stage3_10[15],stage3_9[21],stage3_8[35]}
   );
   gpc606_5 gpc3519 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[15],stage3_10[16],stage3_9[22],stage3_8[36]}
   );
   gpc606_5 gpc3520 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[16],stage3_10[17],stage3_9[23],stage3_8[37]}
   );
   gpc615_5 gpc3521 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82]},
      {stage2_10[24]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[4],stage3_11[17],stage3_10[18],stage3_9[24]}
   );
   gpc606_5 gpc3522 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[5],stage3_11[18],stage3_10[19]}
   );
   gpc606_5 gpc3523 (
      {stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[6],stage3_11[19],stage3_10[20]}
   );
   gpc606_5 gpc3524 (
      {stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[7],stage3_11[20],stage3_10[21]}
   );
   gpc606_5 gpc3525 (
      {stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[8],stage3_11[21],stage3_10[22]}
   );
   gpc606_5 gpc3526 (
      {stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[9],stage3_11[22],stage3_10[23]}
   );
   gpc606_5 gpc3527 (
      {stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[6],stage3_12[10],stage3_11[23],stage3_10[24]}
   );
   gpc606_5 gpc3528 (
      {stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[7],stage3_12[11],stage3_11[24],stage3_10[25]}
   );
   gpc615_5 gpc3529 (
      {stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_11[6]},
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage3_14[7],stage3_13[8],stage3_12[12],stage3_11[25],stage3_10[26]}
   );
   gpc615_5 gpc3530 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[7]},
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage3_14[8],stage3_13[9],stage3_12[13],stage3_11[26],stage3_10[27]}
   );
   gpc615_5 gpc3531 (
      {stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81]},
      {stage2_11[8]},
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage3_14[9],stage3_13[10],stage3_12[14],stage3_11[27],stage3_10[28]}
   );
   gpc615_5 gpc3532 (
      {stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_11[9]},
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage3_14[10],stage3_13[11],stage3_12[15],stage3_11[28],stage3_10[29]}
   );
   gpc615_5 gpc3533 (
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[66]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[12],stage3_12[16],stage3_11[29]}
   );
   gpc615_5 gpc3534 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[67]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[13],stage3_12[17],stage3_11[30]}
   );
   gpc615_5 gpc3535 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[68]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[14],stage3_12[18],stage3_11[31]}
   );
   gpc615_5 gpc3536 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_12[69]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[15],stage3_12[19],stage3_11[32]}
   );
   gpc615_5 gpc3537 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34]},
      {stage2_12[70]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[16],stage3_12[20],stage3_11[33]}
   );
   gpc615_5 gpc3538 (
      {stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_12[71]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[17],stage3_12[21],stage3_11[34]}
   );
   gpc615_5 gpc3539 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_12[72]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[18],stage3_12[22],stage3_11[35]}
   );
   gpc615_5 gpc3540 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_12[73]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[18],stage3_13[19],stage3_12[23],stage3_11[36]}
   );
   gpc615_5 gpc3541 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54]},
      {stage2_12[74]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[19],stage3_13[20],stage3_12[24],stage3_11[37]}
   );
   gpc615_5 gpc3542 (
      {stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage2_12[75]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[20],stage3_13[21],stage3_12[25],stage3_11[38]}
   );
   gpc615_5 gpc3543 (
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64]},
      {stage2_12[76]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[21],stage3_13[22],stage3_12[26],stage3_11[39]}
   );
   gpc615_5 gpc3544 (
      {stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69]},
      {stage2_12[77]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[22],stage3_13[23],stage3_12[27],stage3_11[40]}
   );
   gpc615_5 gpc3545 (
      {stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_12[78]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[23],stage3_13[24],stage3_12[28],stage3_11[41]}
   );
   gpc615_5 gpc3546 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_12[79]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[24],stage3_13[25],stage3_12[29],stage3_11[42]}
   );
   gpc615_5 gpc3547 (
      {stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84]},
      {stage2_12[80]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[25],stage3_13[26],stage3_12[30],stage3_11[43]}
   );
   gpc615_5 gpc3548 (
      {stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage2_12[81]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[26],stage3_13[27],stage3_12[31],stage3_11[44]}
   );
   gpc615_5 gpc3549 (
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94]},
      {stage2_12[82]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[27],stage3_13[28],stage3_12[32],stage3_11[45]}
   );
   gpc615_5 gpc3550 (
      {stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99]},
      {stage2_12[83]},
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage3_15[17],stage3_14[28],stage3_13[29],stage3_12[33],stage3_11[46]}
   );
   gpc615_5 gpc3551 (
      {stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_12[84]},
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage3_15[18],stage3_14[29],stage3_13[30],stage3_12[34],stage3_11[47]}
   );
   gpc615_5 gpc3552 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109]},
      {stage2_12[85]},
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage3_15[19],stage3_14[30],stage3_13[31],stage3_12[35],stage3_11[48]}
   );
   gpc606_5 gpc3553 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[20],stage3_14[31],stage3_13[32],stage3_12[36]}
   );
   gpc615_5 gpc3554 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[21],stage3_14[32]}
   );
   gpc615_5 gpc3555 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[22],stage3_14[33]}
   );
   gpc615_5 gpc3556 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[23],stage3_14[34]}
   );
   gpc615_5 gpc3557 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[4],stage3_15[24],stage3_14[35]}
   );
   gpc615_5 gpc3558 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[5],stage3_15[25],stage3_14[36]}
   );
   gpc615_5 gpc3559 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[5]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[5],stage3_16[6],stage3_15[26],stage3_14[37]}
   );
   gpc615_5 gpc3560 (
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40]},
      {stage2_15[6]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[6],stage3_16[7],stage3_15[27],stage3_14[38]}
   );
   gpc615_5 gpc3561 (
      {stage2_14[41], stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45]},
      {stage2_15[7]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[7],stage3_16[8],stage3_15[28],stage3_14[39]}
   );
   gpc615_5 gpc3562 (
      {stage2_14[46], stage2_14[47], stage2_14[48], stage2_14[49], stage2_14[50]},
      {stage2_15[8]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[8],stage3_16[9],stage3_15[29],stage3_14[40]}
   );
   gpc615_5 gpc3563 (
      {stage2_14[51], stage2_14[52], stage2_14[53], stage2_14[54], stage2_14[55]},
      {stage2_15[9]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[9],stage3_16[10],stage3_15[30],stage3_14[41]}
   );
   gpc615_5 gpc3564 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[10],stage3_16[11],stage3_15[31]}
   );
   gpc615_5 gpc3565 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[11],stage3_16[12],stage3_15[32]}
   );
   gpc615_5 gpc3566 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[12],stage3_16[13],stage3_15[33]}
   );
   gpc615_5 gpc3567 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[13],stage3_16[14],stage3_15[34]}
   );
   gpc615_5 gpc3568 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[14],stage3_16[15],stage3_15[35]}
   );
   gpc615_5 gpc3569 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[15],stage3_16[16],stage3_15[36]}
   );
   gpc615_5 gpc3570 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[16],stage3_16[17],stage3_15[37]}
   );
   gpc615_5 gpc3571 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[17],stage3_16[18],stage3_15[38]}
   );
   gpc615_5 gpc3572 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[68]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[18],stage3_17[18],stage3_16[19],stage3_15[39]}
   );
   gpc615_5 gpc3573 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[69]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[19],stage3_17[19],stage3_16[20],stage3_15[40]}
   );
   gpc615_5 gpc3574 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[70]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[20],stage3_17[20],stage3_16[21],stage3_15[41]}
   );
   gpc615_5 gpc3575 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[71]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[21],stage3_17[21],stage3_16[22],stage3_15[42]}
   );
   gpc135_4 gpc3576 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76]},
      {stage2_17[72], stage2_17[73], stage2_17[74]},
      {stage2_18[0]},
      {stage3_19[12],stage3_18[22],stage3_17[22],stage3_16[23]}
   );
   gpc606_5 gpc3577 (
      {stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[13],stage3_18[23],stage3_17[23],stage3_16[24]}
   );
   gpc606_5 gpc3578 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[14],stage3_18[24]}
   );
   gpc606_5 gpc3579 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[15],stage3_18[25]}
   );
   gpc606_5 gpc3580 (
      {stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[16],stage3_18[26]}
   );
   gpc606_5 gpc3581 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[17],stage3_18[27]}
   );
   gpc606_5 gpc3582 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35], stage2_18[36]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[18],stage3_18[28]}
   );
   gpc606_5 gpc3583 (
      {stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41], stage2_18[42]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[19],stage3_18[29]}
   );
   gpc606_5 gpc3584 (
      {stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[20],stage3_18[30]}
   );
   gpc606_5 gpc3585 (
      {stage2_18[49], stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[21],stage3_18[31]}
   );
   gpc606_5 gpc3586 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[22],stage3_18[32]}
   );
   gpc606_5 gpc3587 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[23],stage3_18[33]}
   );
   gpc606_5 gpc3588 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71], stage2_18[72]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[24],stage3_18[34]}
   );
   gpc606_5 gpc3589 (
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[25]}
   );
   gpc606_5 gpc3590 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[26]}
   );
   gpc606_5 gpc3591 (
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[27]}
   );
   gpc606_5 gpc3592 (
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[28]}
   );
   gpc606_5 gpc3593 (
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[29]}
   );
   gpc606_5 gpc3594 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[5],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[30]}
   );
   gpc606_5 gpc3595 (
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[6],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[31]}
   );
   gpc606_5 gpc3596 (
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[7],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[32]}
   );
   gpc606_5 gpc3597 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[8],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[33]}
   );
   gpc615_5 gpc3598 (
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58]},
      {stage2_20[66]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[9],stage3_22[20],stage3_21[20],stage3_20[21],stage3_19[34]}
   );
   gpc615_5 gpc3599 (
      {stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[67]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[10],stage3_22[21],stage3_21[21],stage3_20[22],stage3_19[35]}
   );
   gpc606_5 gpc3600 (
      {stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71], stage2_20[72], stage2_20[73]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[11],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc606_5 gpc3601 (
      {stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77], stage2_20[78], stage2_20[79]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[12],stage3_22[23],stage3_21[23],stage3_20[24]}
   );
   gpc606_5 gpc3602 (
      {stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83], stage2_20[84], stage2_20[85]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[13],stage3_22[24],stage3_21[24],stage3_20[25]}
   );
   gpc606_5 gpc3603 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[14],stage3_22[25],stage3_21[25],stage3_20[26]}
   );
   gpc606_5 gpc3604 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[15],stage3_22[26],stage3_21[26],stage3_20[27]}
   );
   gpc606_5 gpc3605 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[16],stage3_22[27],stage3_21[27],stage3_20[28]}
   );
   gpc606_5 gpc3606 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[17],stage3_22[28],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3607 (
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[7],stage3_23[18],stage3_22[29],stage3_21[29]}
   );
   gpc606_5 gpc3608 (
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[8],stage3_23[19],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc3609 (
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[9],stage3_23[20],stage3_22[31],stage3_21[31]}
   );
   gpc606_5 gpc3610 (
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[10],stage3_23[21],stage3_22[32],stage3_21[32]}
   );
   gpc606_5 gpc3611 (
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[11],stage3_23[22],stage3_22[33],stage3_21[33]}
   );
   gpc615_5 gpc3612 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[30]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[5],stage3_24[12],stage3_23[23],stage3_22[34]}
   );
   gpc615_5 gpc3613 (
      {stage2_22[47], stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51]},
      {stage2_23[31]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[6],stage3_24[13],stage3_23[24],stage3_22[35]}
   );
   gpc615_5 gpc3614 (
      {stage2_22[52], stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56]},
      {stage2_23[32]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[7],stage3_24[14],stage3_23[25],stage3_22[36]}
   );
   gpc615_5 gpc3615 (
      {stage2_22[57], stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61]},
      {stage2_23[33]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[8],stage3_24[15],stage3_23[26],stage3_22[37]}
   );
   gpc615_5 gpc3616 (
      {stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66]},
      {stage2_23[34]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[9],stage3_24[16],stage3_23[27],stage3_22[38]}
   );
   gpc615_5 gpc3617 (
      {stage2_22[67], stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71]},
      {stage2_23[35]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[10],stage3_24[17],stage3_23[28],stage3_22[39]}
   );
   gpc615_5 gpc3618 (
      {stage2_22[72], stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76]},
      {stage2_23[36]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[11],stage3_24[18],stage3_23[29],stage3_22[40]}
   );
   gpc615_5 gpc3619 (
      {stage2_22[77], stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81]},
      {stage2_23[37]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[12],stage3_24[19],stage3_23[30],stage3_22[41]}
   );
   gpc615_5 gpc3620 (
      {stage2_22[82], stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86]},
      {stage2_23[38]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[13],stage3_24[20],stage3_23[31],stage3_22[42]}
   );
   gpc606_5 gpc3621 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[9],stage3_25[14],stage3_24[21],stage3_23[32]}
   );
   gpc606_5 gpc3622 (
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[10],stage3_25[15],stage3_24[22],stage3_23[33]}
   );
   gpc606_5 gpc3623 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[11],stage3_25[16],stage3_24[23],stage3_23[34]}
   );
   gpc606_5 gpc3624 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[12],stage3_25[17],stage3_24[24],stage3_23[35]}
   );
   gpc606_5 gpc3625 (
      {stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[13],stage3_25[18],stage3_24[25],stage3_23[36]}
   );
   gpc606_5 gpc3626 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[14],stage3_25[19],stage3_24[26],stage3_23[37]}
   );
   gpc606_5 gpc3627 (
      {stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[15],stage3_25[20],stage3_24[27],stage3_23[38]}
   );
   gpc606_5 gpc3628 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85], stage2_23[86]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[16],stage3_25[21],stage3_24[28],stage3_23[39]}
   );
   gpc606_5 gpc3629 (
      {stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90], stage2_23[91], stage2_23[92]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[17],stage3_25[22],stage3_24[29],stage3_23[40]}
   );
   gpc606_5 gpc3630 (
      {stage2_23[93], stage2_23[94], stage2_23[95], stage2_23[96], stage2_23[97], stage2_23[98]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[18],stage3_25[23],stage3_24[30],stage3_23[41]}
   );
   gpc606_5 gpc3631 (
      {stage2_23[99], stage2_23[100], stage2_23[101], stage2_23[102], stage2_23[103], stage2_23[104]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[19],stage3_25[24],stage3_24[31],stage3_23[42]}
   );
   gpc606_5 gpc3632 (
      {stage2_23[105], stage2_23[106], stage2_23[107], stage2_23[108], stage2_23[109], stage2_23[110]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[20],stage3_25[25],stage3_24[32],stage3_23[43]}
   );
   gpc606_5 gpc3633 (
      {stage2_23[111], stage2_23[112], stage2_23[113], stage2_23[114], stage2_23[115], stage2_23[116]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[21],stage3_25[26],stage3_24[33],stage3_23[44]}
   );
   gpc606_5 gpc3634 (
      {stage2_23[117], stage2_23[118], stage2_23[119], stage2_23[120], stage2_23[121], stage2_23[122]},
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage3_27[13],stage3_26[22],stage3_25[27],stage3_24[34],stage3_23[45]}
   );
   gpc606_5 gpc3635 (
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[14],stage3_26[23],stage3_25[28],stage3_24[35]}
   );
   gpc606_5 gpc3636 (
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[15],stage3_26[24],stage3_25[29],stage3_24[36]}
   );
   gpc1163_5 gpc3637 (
      {stage2_26[12], stage2_26[13], stage2_26[14]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage2_28[0]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[0],stage3_28[2],stage3_27[16],stage3_26[25]}
   );
   gpc606_5 gpc3638 (
      {stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6]},
      {stage3_30[1],stage3_29[1],stage3_28[3],stage3_27[17],stage3_26[26]}
   );
   gpc606_5 gpc3639 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26]},
      {stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12]},
      {stage3_30[2],stage3_29[2],stage3_28[4],stage3_27[18],stage3_26[27]}
   );
   gpc606_5 gpc3640 (
      {stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18]},
      {stage3_30[3],stage3_29[3],stage3_28[5],stage3_27[19],stage3_26[28]}
   );
   gpc606_5 gpc3641 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23], stage2_28[24]},
      {stage3_30[4],stage3_29[4],stage3_28[6],stage3_27[20],stage3_26[29]}
   );
   gpc606_5 gpc3642 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44]},
      {stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28], stage2_28[29], stage2_28[30]},
      {stage3_30[5],stage3_29[5],stage3_28[7],stage3_27[21],stage3_26[30]}
   );
   gpc606_5 gpc3643 (
      {stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50]},
      {stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35], stage2_28[36]},
      {stage3_30[6],stage3_29[6],stage3_28[8],stage3_27[22],stage3_26[31]}
   );
   gpc606_5 gpc3644 (
      {stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56]},
      {stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42]},
      {stage3_30[7],stage3_29[7],stage3_28[9],stage3_27[23],stage3_26[32]}
   );
   gpc606_5 gpc3645 (
      {stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage3_30[8],stage3_29[8],stage3_28[10],stage3_27[24],stage3_26[33]}
   );
   gpc606_5 gpc3646 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68]},
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53], stage2_28[54]},
      {stage3_30[9],stage3_29[9],stage3_28[11],stage3_27[25],stage3_26[34]}
   );
   gpc606_5 gpc3647 (
      {stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74]},
      {stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58], stage2_28[59], stage2_28[60]},
      {stage3_30[10],stage3_29[10],stage3_28[12],stage3_27[26],stage3_26[35]}
   );
   gpc606_5 gpc3648 (
      {stage2_26[75], stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80]},
      {stage2_28[61], stage2_28[62], stage2_28[63], stage2_28[64], stage2_28[65], stage2_28[66]},
      {stage3_30[11],stage3_29[11],stage3_28[13],stage3_27[27],stage3_26[36]}
   );
   gpc606_5 gpc3649 (
      {stage2_26[81], stage2_26[82], stage2_26[83], stage2_26[84], stage2_26[85], stage2_26[86]},
      {stage2_28[67], stage2_28[68], stage2_28[69], stage2_28[70], stage2_28[71], stage2_28[72]},
      {stage3_30[12],stage3_29[12],stage3_28[14],stage3_27[28],stage3_26[37]}
   );
   gpc606_5 gpc3650 (
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[13],stage3_29[13],stage3_28[15],stage3_27[29]}
   );
   gpc615_5 gpc3651 (
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16]},
      {stage2_28[73]},
      {stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11], stage2_29[12]},
      {stage3_31[1],stage3_30[14],stage3_29[14],stage3_28[16],stage3_27[30]}
   );
   gpc615_5 gpc3652 (
      {stage2_27[17], stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21]},
      {stage2_28[74]},
      {stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage3_31[2],stage3_30[15],stage3_29[15],stage3_28[17],stage3_27[31]}
   );
   gpc615_5 gpc3653 (
      {stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26]},
      {stage2_28[75]},
      {stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage3_31[3],stage3_30[16],stage3_29[16],stage3_28[18],stage3_27[32]}
   );
   gpc615_5 gpc3654 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31]},
      {stage2_28[76]},
      {stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage3_31[4],stage3_30[17],stage3_29[17],stage3_28[19],stage3_27[33]}
   );
   gpc615_5 gpc3655 (
      {stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36]},
      {stage2_28[77]},
      {stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35], stage2_29[36]},
      {stage3_31[5],stage3_30[18],stage3_29[18],stage3_28[20],stage3_27[34]}
   );
   gpc615_5 gpc3656 (
      {stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[78]},
      {stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41], stage2_29[42]},
      {stage3_31[6],stage3_30[19],stage3_29[19],stage3_28[21],stage3_27[35]}
   );
   gpc615_5 gpc3657 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[79]},
      {stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47], stage2_29[48]},
      {stage3_31[7],stage3_30[20],stage3_29[20],stage3_28[22],stage3_27[36]}
   );
   gpc615_5 gpc3658 (
      {stage2_27[47], stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51]},
      {stage2_28[80]},
      {stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53], stage2_29[54]},
      {stage3_31[8],stage3_30[21],stage3_29[21],stage3_28[23],stage3_27[37]}
   );
   gpc615_5 gpc3659 (
      {stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[81]},
      {stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59], stage2_29[60]},
      {stage3_31[9],stage3_30[22],stage3_29[22],stage3_28[24],stage3_27[38]}
   );
   gpc615_5 gpc3660 (
      {stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61]},
      {stage2_28[82]},
      {stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65], stage2_29[66]},
      {stage3_31[10],stage3_30[23],stage3_29[23],stage3_28[25],stage3_27[39]}
   );
   gpc615_5 gpc3661 (
      {stage2_27[62], stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66]},
      {stage2_28[83]},
      {stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71], stage2_29[72]},
      {stage3_31[11],stage3_30[24],stage3_29[24],stage3_28[26],stage3_27[40]}
   );
   gpc615_5 gpc3662 (
      {stage2_27[67], stage2_27[68], stage2_27[69], stage2_27[70], stage2_27[71]},
      {stage2_28[84]},
      {stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77], stage2_29[78]},
      {stage3_31[12],stage3_30[25],stage3_29[25],stage3_28[27],stage3_27[41]}
   );
   gpc606_5 gpc3663 (
      {stage2_28[85], stage2_28[86], stage2_28[87], stage2_28[88], stage2_28[89], stage2_28[90]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[13],stage3_30[26],stage3_29[26],stage3_28[28]}
   );
   gpc606_5 gpc3664 (
      {stage2_28[91], stage2_28[92], stage2_28[93], stage2_28[94], stage2_28[95], stage2_28[96]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[14],stage3_30[27],stage3_29[27],stage3_28[29]}
   );
   gpc606_5 gpc3665 (
      {stage2_28[97], stage2_28[98], stage2_28[99], stage2_28[100], stage2_28[101], stage2_28[102]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[15],stage3_30[28],stage3_29[28],stage3_28[30]}
   );
   gpc606_5 gpc3666 (
      {stage2_28[103], stage2_28[104], stage2_28[105], stage2_28[106], stage2_28[107], stage2_28[108]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[16],stage3_30[29],stage3_29[29],stage3_28[31]}
   );
   gpc606_5 gpc3667 (
      {stage2_28[109], stage2_28[110], stage2_28[111], stage2_28[112], stage2_28[113], stage2_28[114]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[17],stage3_30[30],stage3_29[30],stage3_28[32]}
   );
   gpc606_5 gpc3668 (
      {stage2_28[115], stage2_28[116], stage2_28[117], stage2_28[118], stage2_28[119], stage2_28[120]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[18],stage3_30[31],stage3_29[31],stage3_28[33]}
   );
   gpc606_5 gpc3669 (
      {stage2_28[121], stage2_28[122], stage2_28[123], stage2_28[124], stage2_28[125], stage2_28[126]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[19],stage3_30[32],stage3_29[32],stage3_28[34]}
   );
   gpc606_5 gpc3670 (
      {stage2_28[127], stage2_28[128], stage2_28[129], stage2_28[130], stage2_28[131], stage2_28[132]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[20],stage3_30[33],stage3_29[33],stage3_28[35]}
   );
   gpc606_5 gpc3671 (
      {stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83], stage2_29[84]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[8],stage3_31[21],stage3_30[34],stage3_29[34]}
   );
   gpc606_5 gpc3672 (
      {stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89], stage2_29[90]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[9],stage3_31[22],stage3_30[35],stage3_29[35]}
   );
   gpc606_5 gpc3673 (
      {stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95], stage2_29[96]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[10],stage3_31[23],stage3_30[36],stage3_29[36]}
   );
   gpc606_5 gpc3674 (
      {stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101], stage2_29[102]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[11],stage3_31[24],stage3_30[37],stage3_29[37]}
   );
   gpc606_5 gpc3675 (
      {stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106], stage2_29[107], stage2_29[108]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[12],stage3_31[25],stage3_30[38],stage3_29[38]}
   );
   gpc606_5 gpc3676 (
      {stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112], stage2_29[113], stage2_29[114]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[5],stage3_32[13],stage3_31[26],stage3_30[39],stage3_29[39]}
   );
   gpc606_5 gpc3677 (
      {stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118], stage2_29[119], stage2_29[120]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[6],stage3_32[14],stage3_31[27],stage3_30[40],stage3_29[40]}
   );
   gpc606_5 gpc3678 (
      {stage2_29[121], stage2_29[122], stage2_29[123], stage2_29[124], stage2_29[125], stage2_29[126]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[7],stage3_32[15],stage3_31[28],stage3_30[41],stage3_29[41]}
   );
   gpc606_5 gpc3679 (
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[8],stage3_32[16],stage3_31[29],stage3_30[42]}
   );
   gpc606_5 gpc3680 (
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[9],stage3_32[17],stage3_31[30],stage3_30[43]}
   );
   gpc606_5 gpc3681 (
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[10],stage3_32[18],stage3_31[31],stage3_30[44]}
   );
   gpc615_5 gpc3682 (
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[11],stage3_32[19],stage3_31[32]}
   );
   gpc615_5 gpc3683 (
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[12],stage3_32[20],stage3_31[33]}
   );
   gpc615_5 gpc3684 (
      {stage2_31[58], stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[13],stage3_32[21],stage3_31[34]}
   );
   gpc615_5 gpc3685 (
      {stage2_31[63], stage2_31[64], stage2_31[65], stage2_31[66], stage2_31[67]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[14],stage3_32[22],stage3_31[35]}
   );
   gpc615_5 gpc3686 (
      {stage2_31[68], stage2_31[69], stage2_31[70], stage2_31[71], stage2_31[72]},
      {stage2_32[22]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[7],stage3_33[15],stage3_32[23],stage3_31[36]}
   );
   gpc615_5 gpc3687 (
      {stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76], stage2_31[77]},
      {stage2_32[23]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[8],stage3_33[16],stage3_32[24],stage3_31[37]}
   );
   gpc615_5 gpc3688 (
      {stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_32[24]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[9],stage3_33[17],stage3_32[25],stage3_31[38]}
   );
   gpc606_5 gpc3689 (
      {stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[10],stage3_33[18],stage3_32[26]}
   );
   gpc615_5 gpc3690 (
      {stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_33[42]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[11],stage3_33[19],stage3_32[27]}
   );
   gpc615_5 gpc3691 (
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_33[43]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[12],stage3_33[20],stage3_32[28]}
   );
   gpc615_5 gpc3692 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[44]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[13],stage3_33[21],stage3_32[29]}
   );
   gpc606_5 gpc3693 (
      {stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48], stage2_33[49], stage2_33[50]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[4],stage3_35[11],stage3_34[14],stage3_33[22]}
   );
   gpc606_5 gpc3694 (
      {stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54], stage2_33[55], stage2_33[56]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[5],stage3_35[12],stage3_34[15],stage3_33[23]}
   );
   gpc1_1 gpc3695 (
      {stage2_1[48]},
      {stage3_1[18]}
   );
   gpc1_1 gpc3696 (
      {stage2_1[49]},
      {stage3_1[19]}
   );
   gpc1_1 gpc3697 (
      {stage2_1[50]},
      {stage3_1[20]}
   );
   gpc1_1 gpc3698 (
      {stage2_1[51]},
      {stage3_1[21]}
   );
   gpc1_1 gpc3699 (
      {stage2_1[52]},
      {stage3_1[22]}
   );
   gpc1_1 gpc3700 (
      {stage2_1[53]},
      {stage3_1[23]}
   );
   gpc1_1 gpc3701 (
      {stage2_1[54]},
      {stage3_1[24]}
   );
   gpc1_1 gpc3702 (
      {stage2_1[55]},
      {stage3_1[25]}
   );
   gpc1_1 gpc3703 (
      {stage2_2[81]},
      {stage3_2[22]}
   );
   gpc1_1 gpc3704 (
      {stage2_2[82]},
      {stage3_2[23]}
   );
   gpc1_1 gpc3705 (
      {stage2_2[83]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3706 (
      {stage2_2[84]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3707 (
      {stage2_2[85]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3708 (
      {stage2_2[86]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3709 (
      {stage2_2[87]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3710 (
      {stage2_2[88]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3711 (
      {stage2_2[89]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3712 (
      {stage2_2[90]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3713 (
      {stage2_2[91]},
      {stage3_2[32]}
   );
   gpc1_1 gpc3714 (
      {stage2_2[92]},
      {stage3_2[33]}
   );
   gpc1_1 gpc3715 (
      {stage2_2[93]},
      {stage3_2[34]}
   );
   gpc1_1 gpc3716 (
      {stage2_2[94]},
      {stage3_2[35]}
   );
   gpc1_1 gpc3717 (
      {stage2_4[114]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3718 (
      {stage2_4[115]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3719 (
      {stage2_4[116]},
      {stage3_4[44]}
   );
   gpc1_1 gpc3720 (
      {stage2_4[117]},
      {stage3_4[45]}
   );
   gpc1_1 gpc3721 (
      {stage2_4[118]},
      {stage3_4[46]}
   );
   gpc1_1 gpc3722 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3723 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3724 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3725 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3726 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3727 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3728 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3729 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3730 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3731 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3732 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3733 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3734 (
      {stage2_5[84]},
      {stage3_5[49]}
   );
   gpc1_1 gpc3735 (
      {stage2_5[85]},
      {stage3_5[50]}
   );
   gpc1_1 gpc3736 (
      {stage2_5[86]},
      {stage3_5[51]}
   );
   gpc1_1 gpc3737 (
      {stage2_5[87]},
      {stage3_5[52]}
   );
   gpc1_1 gpc3738 (
      {stage2_5[88]},
      {stage3_5[53]}
   );
   gpc1_1 gpc3739 (
      {stage2_5[89]},
      {stage3_5[54]}
   );
   gpc1_1 gpc3740 (
      {stage2_5[90]},
      {stage3_5[55]}
   );
   gpc1_1 gpc3741 (
      {stage2_5[91]},
      {stage3_5[56]}
   );
   gpc1_1 gpc3742 (
      {stage2_5[92]},
      {stage3_5[57]}
   );
   gpc1_1 gpc3743 (
      {stage2_5[93]},
      {stage3_5[58]}
   );
   gpc1_1 gpc3744 (
      {stage2_6[89]},
      {stage3_6[31]}
   );
   gpc1_1 gpc3745 (
      {stage2_6[90]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3746 (
      {stage2_6[91]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3747 (
      {stage2_6[92]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3748 (
      {stage2_6[93]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3749 (
      {stage2_6[94]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3750 (
      {stage2_6[95]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3751 (
      {stage2_7[102]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3752 (
      {stage2_7[103]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3753 (
      {stage2_7[104]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3754 (
      {stage2_7[105]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3755 (
      {stage2_7[106]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3756 (
      {stage2_7[107]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3757 (
      {stage2_7[108]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3758 (
      {stage2_8[43]},
      {stage3_8[38]}
   );
   gpc1_1 gpc3759 (
      {stage2_8[44]},
      {stage3_8[39]}
   );
   gpc1_1 gpc3760 (
      {stage2_8[45]},
      {stage3_8[40]}
   );
   gpc1_1 gpc3761 (
      {stage2_8[46]},
      {stage3_8[41]}
   );
   gpc1_1 gpc3762 (
      {stage2_8[47]},
      {stage3_8[42]}
   );
   gpc1_1 gpc3763 (
      {stage2_8[48]},
      {stage3_8[43]}
   );
   gpc1_1 gpc3764 (
      {stage2_8[49]},
      {stage3_8[44]}
   );
   gpc1_1 gpc3765 (
      {stage2_8[50]},
      {stage3_8[45]}
   );
   gpc1_1 gpc3766 (
      {stage2_8[51]},
      {stage3_8[46]}
   );
   gpc1_1 gpc3767 (
      {stage2_8[52]},
      {stage3_8[47]}
   );
   gpc1_1 gpc3768 (
      {stage2_8[53]},
      {stage3_8[48]}
   );
   gpc1_1 gpc3769 (
      {stage2_8[54]},
      {stage3_8[49]}
   );
   gpc1_1 gpc3770 (
      {stage2_8[55]},
      {stage3_8[50]}
   );
   gpc1_1 gpc3771 (
      {stage2_8[56]},
      {stage3_8[51]}
   );
   gpc1_1 gpc3772 (
      {stage2_8[57]},
      {stage3_8[52]}
   );
   gpc1_1 gpc3773 (
      {stage2_8[58]},
      {stage3_8[53]}
   );
   gpc1_1 gpc3774 (
      {stage2_8[59]},
      {stage3_8[54]}
   );
   gpc1_1 gpc3775 (
      {stage2_8[60]},
      {stage3_8[55]}
   );
   gpc1_1 gpc3776 (
      {stage2_8[61]},
      {stage3_8[56]}
   );
   gpc1_1 gpc3777 (
      {stage2_8[62]},
      {stage3_8[57]}
   );
   gpc1_1 gpc3778 (
      {stage2_8[63]},
      {stage3_8[58]}
   );
   gpc1_1 gpc3779 (
      {stage2_8[64]},
      {stage3_8[59]}
   );
   gpc1_1 gpc3780 (
      {stage2_8[65]},
      {stage3_8[60]}
   );
   gpc1_1 gpc3781 (
      {stage2_8[66]},
      {stage3_8[61]}
   );
   gpc1_1 gpc3782 (
      {stage2_8[67]},
      {stage3_8[62]}
   );
   gpc1_1 gpc3783 (
      {stage2_8[68]},
      {stage3_8[63]}
   );
   gpc1_1 gpc3784 (
      {stage2_8[69]},
      {stage3_8[64]}
   );
   gpc1_1 gpc3785 (
      {stage2_8[70]},
      {stage3_8[65]}
   );
   gpc1_1 gpc3786 (
      {stage2_8[71]},
      {stage3_8[66]}
   );
   gpc1_1 gpc3787 (
      {stage2_8[72]},
      {stage3_8[67]}
   );
   gpc1_1 gpc3788 (
      {stage2_8[73]},
      {stage3_8[68]}
   );
   gpc1_1 gpc3789 (
      {stage2_8[74]},
      {stage3_8[69]}
   );
   gpc1_1 gpc3790 (
      {stage2_8[75]},
      {stage3_8[70]}
   );
   gpc1_1 gpc3791 (
      {stage2_8[76]},
      {stage3_8[71]}
   );
   gpc1_1 gpc3792 (
      {stage2_8[77]},
      {stage3_8[72]}
   );
   gpc1_1 gpc3793 (
      {stage2_8[78]},
      {stage3_8[73]}
   );
   gpc1_1 gpc3794 (
      {stage2_8[79]},
      {stage3_8[74]}
   );
   gpc1_1 gpc3795 (
      {stage2_8[80]},
      {stage3_8[75]}
   );
   gpc1_1 gpc3796 (
      {stage2_8[81]},
      {stage3_8[76]}
   );
   gpc1_1 gpc3797 (
      {stage2_8[82]},
      {stage3_8[77]}
   );
   gpc1_1 gpc3798 (
      {stage2_8[83]},
      {stage3_8[78]}
   );
   gpc1_1 gpc3799 (
      {stage2_8[84]},
      {stage3_8[79]}
   );
   gpc1_1 gpc3800 (
      {stage2_8[85]},
      {stage3_8[80]}
   );
   gpc1_1 gpc3801 (
      {stage2_8[86]},
      {stage3_8[81]}
   );
   gpc1_1 gpc3802 (
      {stage2_8[87]},
      {stage3_8[82]}
   );
   gpc1_1 gpc3803 (
      {stage2_8[88]},
      {stage3_8[83]}
   );
   gpc1_1 gpc3804 (
      {stage2_8[89]},
      {stage3_8[84]}
   );
   gpc1_1 gpc3805 (
      {stage2_8[90]},
      {stage3_8[85]}
   );
   gpc1_1 gpc3806 (
      {stage2_8[91]},
      {stage3_8[86]}
   );
   gpc1_1 gpc3807 (
      {stage2_8[92]},
      {stage3_8[87]}
   );
   gpc1_1 gpc3808 (
      {stage2_8[93]},
      {stage3_8[88]}
   );
   gpc1_1 gpc3809 (
      {stage2_8[94]},
      {stage3_8[89]}
   );
   gpc1_1 gpc3810 (
      {stage2_8[95]},
      {stage3_8[90]}
   );
   gpc1_1 gpc3811 (
      {stage2_8[96]},
      {stage3_8[91]}
   );
   gpc1_1 gpc3812 (
      {stage2_8[97]},
      {stage3_8[92]}
   );
   gpc1_1 gpc3813 (
      {stage2_9[83]},
      {stage3_9[25]}
   );
   gpc1_1 gpc3814 (
      {stage2_9[84]},
      {stage3_9[26]}
   );
   gpc1_1 gpc3815 (
      {stage2_9[85]},
      {stage3_9[27]}
   );
   gpc1_1 gpc3816 (
      {stage2_9[86]},
      {stage3_9[28]}
   );
   gpc1_1 gpc3817 (
      {stage2_9[87]},
      {stage3_9[29]}
   );
   gpc1_1 gpc3818 (
      {stage2_9[88]},
      {stage3_9[30]}
   );
   gpc1_1 gpc3819 (
      {stage2_9[89]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3820 (
      {stage2_9[90]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3821 (
      {stage2_9[91]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3822 (
      {stage2_9[92]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3823 (
      {stage2_9[93]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3824 (
      {stage2_9[94]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3825 (
      {stage2_9[95]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3826 (
      {stage2_9[96]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3827 (
      {stage2_9[97]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3828 (
      {stage2_9[98]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3829 (
      {stage2_9[99]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3830 (
      {stage2_9[100]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3831 (
      {stage2_9[101]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3832 (
      {stage2_9[102]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3833 (
      {stage2_9[103]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3834 (
      {stage2_9[104]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3835 (
      {stage2_9[105]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3836 (
      {stage2_9[106]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3837 (
      {stage2_9[107]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3838 (
      {stage2_10[87]},
      {stage3_10[30]}
   );
   gpc1_1 gpc3839 (
      {stage2_10[88]},
      {stage3_10[31]}
   );
   gpc1_1 gpc3840 (
      {stage2_10[89]},
      {stage3_10[32]}
   );
   gpc1_1 gpc3841 (
      {stage2_10[90]},
      {stage3_10[33]}
   );
   gpc1_1 gpc3842 (
      {stage2_10[91]},
      {stage3_10[34]}
   );
   gpc1_1 gpc3843 (
      {stage2_10[92]},
      {stage3_10[35]}
   );
   gpc1_1 gpc3844 (
      {stage2_10[93]},
      {stage3_10[36]}
   );
   gpc1_1 gpc3845 (
      {stage2_10[94]},
      {stage3_10[37]}
   );
   gpc1_1 gpc3846 (
      {stage2_11[110]},
      {stage3_11[49]}
   );
   gpc1_1 gpc3847 (
      {stage2_11[111]},
      {stage3_11[50]}
   );
   gpc1_1 gpc3848 (
      {stage2_11[112]},
      {stage3_11[51]}
   );
   gpc1_1 gpc3849 (
      {stage2_11[113]},
      {stage3_11[52]}
   );
   gpc1_1 gpc3850 (
      {stage2_11[114]},
      {stage3_11[53]}
   );
   gpc1_1 gpc3851 (
      {stage2_11[115]},
      {stage3_11[54]}
   );
   gpc1_1 gpc3852 (
      {stage2_12[92]},
      {stage3_12[37]}
   );
   gpc1_1 gpc3853 (
      {stage2_12[93]},
      {stage3_12[38]}
   );
   gpc1_1 gpc3854 (
      {stage2_12[94]},
      {stage3_12[39]}
   );
   gpc1_1 gpc3855 (
      {stage2_12[95]},
      {stage3_12[40]}
   );
   gpc1_1 gpc3856 (
      {stage2_12[96]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3857 (
      {stage2_12[97]},
      {stage3_12[42]}
   );
   gpc1_1 gpc3858 (
      {stage2_12[98]},
      {stage3_12[43]}
   );
   gpc1_1 gpc3859 (
      {stage2_12[99]},
      {stage3_12[44]}
   );
   gpc1_1 gpc3860 (
      {stage2_12[100]},
      {stage3_12[45]}
   );
   gpc1_1 gpc3861 (
      {stage2_12[101]},
      {stage3_12[46]}
   );
   gpc1_1 gpc3862 (
      {stage2_13[120]},
      {stage3_13[33]}
   );
   gpc1_1 gpc3863 (
      {stage2_13[121]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3864 (
      {stage2_13[122]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3865 (
      {stage2_13[123]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3866 (
      {stage2_14[56]},
      {stage3_14[42]}
   );
   gpc1_1 gpc3867 (
      {stage2_14[57]},
      {stage3_14[43]}
   );
   gpc1_1 gpc3868 (
      {stage2_14[58]},
      {stage3_14[44]}
   );
   gpc1_1 gpc3869 (
      {stage2_14[59]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3870 (
      {stage2_14[60]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3871 (
      {stage2_14[61]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3872 (
      {stage2_14[62]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3873 (
      {stage2_14[63]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3874 (
      {stage2_14[64]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3875 (
      {stage2_14[65]},
      {stage3_14[51]}
   );
   gpc1_1 gpc3876 (
      {stage2_14[66]},
      {stage3_14[52]}
   );
   gpc1_1 gpc3877 (
      {stage2_14[67]},
      {stage3_14[53]}
   );
   gpc1_1 gpc3878 (
      {stage2_14[68]},
      {stage3_14[54]}
   );
   gpc1_1 gpc3879 (
      {stage2_14[69]},
      {stage3_14[55]}
   );
   gpc1_1 gpc3880 (
      {stage2_15[70]},
      {stage3_15[43]}
   );
   gpc1_1 gpc3881 (
      {stage2_15[71]},
      {stage3_15[44]}
   );
   gpc1_1 gpc3882 (
      {stage2_15[72]},
      {stage3_15[45]}
   );
   gpc1_1 gpc3883 (
      {stage2_15[73]},
      {stage3_15[46]}
   );
   gpc1_1 gpc3884 (
      {stage2_15[74]},
      {stage3_15[47]}
   );
   gpc1_1 gpc3885 (
      {stage2_15[75]},
      {stage3_15[48]}
   );
   gpc1_1 gpc3886 (
      {stage2_15[76]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3887 (
      {stage2_15[77]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3888 (
      {stage2_15[78]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3889 (
      {stage2_15[79]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3890 (
      {stage2_15[80]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3891 (
      {stage2_15[81]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3892 (
      {stage2_15[82]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3893 (
      {stage2_15[83]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3894 (
      {stage2_15[84]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3895 (
      {stage2_15[85]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3896 (
      {stage2_15[86]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3897 (
      {stage2_15[87]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3898 (
      {stage2_15[88]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3899 (
      {stage2_15[89]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3900 (
      {stage2_15[90]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3901 (
      {stage2_15[91]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3902 (
      {stage2_15[92]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3903 (
      {stage2_15[93]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3904 (
      {stage2_15[94]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3905 (
      {stage2_15[95]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3906 (
      {stage2_15[96]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3907 (
      {stage2_15[97]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3908 (
      {stage2_16[83]},
      {stage3_16[25]}
   );
   gpc1_1 gpc3909 (
      {stage2_16[84]},
      {stage3_16[26]}
   );
   gpc1_1 gpc3910 (
      {stage2_16[85]},
      {stage3_16[27]}
   );
   gpc1_1 gpc3911 (
      {stage2_16[86]},
      {stage3_16[28]}
   );
   gpc1_1 gpc3912 (
      {stage2_16[87]},
      {stage3_16[29]}
   );
   gpc1_1 gpc3913 (
      {stage2_16[88]},
      {stage3_16[30]}
   );
   gpc1_1 gpc3914 (
      {stage2_16[89]},
      {stage3_16[31]}
   );
   gpc1_1 gpc3915 (
      {stage2_16[90]},
      {stage3_16[32]}
   );
   gpc1_1 gpc3916 (
      {stage2_16[91]},
      {stage3_16[33]}
   );
   gpc1_1 gpc3917 (
      {stage2_16[92]},
      {stage3_16[34]}
   );
   gpc1_1 gpc3918 (
      {stage2_16[93]},
      {stage3_16[35]}
   );
   gpc1_1 gpc3919 (
      {stage2_16[94]},
      {stage3_16[36]}
   );
   gpc1_1 gpc3920 (
      {stage2_16[95]},
      {stage3_16[37]}
   );
   gpc1_1 gpc3921 (
      {stage2_16[96]},
      {stage3_16[38]}
   );
   gpc1_1 gpc3922 (
      {stage2_16[97]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3923 (
      {stage2_16[98]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3924 (
      {stage2_16[99]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3925 (
      {stage2_16[100]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3926 (
      {stage2_16[101]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3927 (
      {stage2_16[102]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3928 (
      {stage2_16[103]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3929 (
      {stage2_16[104]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3930 (
      {stage2_16[105]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3931 (
      {stage2_16[106]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3932 (
      {stage2_16[107]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3933 (
      {stage2_16[108]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3934 (
      {stage2_16[109]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3935 (
      {stage2_16[110]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3936 (
      {stage2_16[111]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3937 (
      {stage2_16[112]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3938 (
      {stage2_16[113]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3939 (
      {stage2_16[114]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3940 (
      {stage2_16[115]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3941 (
      {stage2_16[116]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3942 (
      {stage2_16[117]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3943 (
      {stage2_16[118]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3944 (
      {stage2_16[119]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3945 (
      {stage2_16[120]},
      {stage3_16[62]}
   );
   gpc1_1 gpc3946 (
      {stage2_16[121]},
      {stage3_16[63]}
   );
   gpc1_1 gpc3947 (
      {stage2_16[122]},
      {stage3_16[64]}
   );
   gpc1_1 gpc3948 (
      {stage2_16[123]},
      {stage3_16[65]}
   );
   gpc1_1 gpc3949 (
      {stage2_16[124]},
      {stage3_16[66]}
   );
   gpc1_1 gpc3950 (
      {stage2_17[75]},
      {stage3_17[24]}
   );
   gpc1_1 gpc3951 (
      {stage2_17[76]},
      {stage3_17[25]}
   );
   gpc1_1 gpc3952 (
      {stage2_17[77]},
      {stage3_17[26]}
   );
   gpc1_1 gpc3953 (
      {stage2_17[78]},
      {stage3_17[27]}
   );
   gpc1_1 gpc3954 (
      {stage2_17[79]},
      {stage3_17[28]}
   );
   gpc1_1 gpc3955 (
      {stage2_17[80]},
      {stage3_17[29]}
   );
   gpc1_1 gpc3956 (
      {stage2_17[81]},
      {stage3_17[30]}
   );
   gpc1_1 gpc3957 (
      {stage2_17[82]},
      {stage3_17[31]}
   );
   gpc1_1 gpc3958 (
      {stage2_17[83]},
      {stage3_17[32]}
   );
   gpc1_1 gpc3959 (
      {stage2_17[84]},
      {stage3_17[33]}
   );
   gpc1_1 gpc3960 (
      {stage2_17[85]},
      {stage3_17[34]}
   );
   gpc1_1 gpc3961 (
      {stage2_17[86]},
      {stage3_17[35]}
   );
   gpc1_1 gpc3962 (
      {stage2_17[87]},
      {stage3_17[36]}
   );
   gpc1_1 gpc3963 (
      {stage2_17[88]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3964 (
      {stage2_17[89]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3965 (
      {stage2_17[90]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3966 (
      {stage2_17[91]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3967 (
      {stage2_17[92]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3968 (
      {stage2_17[93]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3969 (
      {stage2_17[94]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3970 (
      {stage2_17[95]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3971 (
      {stage2_17[96]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3972 (
      {stage2_17[97]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3973 (
      {stage2_17[98]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3974 (
      {stage2_17[99]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3975 (
      {stage2_17[100]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3976 (
      {stage2_17[101]},
      {stage3_17[50]}
   );
   gpc1_1 gpc3977 (
      {stage2_17[102]},
      {stage3_17[51]}
   );
   gpc1_1 gpc3978 (
      {stage2_17[103]},
      {stage3_17[52]}
   );
   gpc1_1 gpc3979 (
      {stage2_17[104]},
      {stage3_17[53]}
   );
   gpc1_1 gpc3980 (
      {stage2_17[105]},
      {stage3_17[54]}
   );
   gpc1_1 gpc3981 (
      {stage2_17[106]},
      {stage3_17[55]}
   );
   gpc1_1 gpc3982 (
      {stage2_17[107]},
      {stage3_17[56]}
   );
   gpc1_1 gpc3983 (
      {stage2_17[108]},
      {stage3_17[57]}
   );
   gpc1_1 gpc3984 (
      {stage2_17[109]},
      {stage3_17[58]}
   );
   gpc1_1 gpc3985 (
      {stage2_17[110]},
      {stage3_17[59]}
   );
   gpc1_1 gpc3986 (
      {stage2_17[111]},
      {stage3_17[60]}
   );
   gpc1_1 gpc3987 (
      {stage2_17[112]},
      {stage3_17[61]}
   );
   gpc1_1 gpc3988 (
      {stage2_17[113]},
      {stage3_17[62]}
   );
   gpc1_1 gpc3989 (
      {stage2_17[114]},
      {stage3_17[63]}
   );
   gpc1_1 gpc3990 (
      {stage2_17[115]},
      {stage3_17[64]}
   );
   gpc1_1 gpc3991 (
      {stage2_17[116]},
      {stage3_17[65]}
   );
   gpc1_1 gpc3992 (
      {stage2_17[117]},
      {stage3_17[66]}
   );
   gpc1_1 gpc3993 (
      {stage2_17[118]},
      {stage3_17[67]}
   );
   gpc1_1 gpc3994 (
      {stage2_17[119]},
      {stage3_17[68]}
   );
   gpc1_1 gpc3995 (
      {stage2_17[120]},
      {stage3_17[69]}
   );
   gpc1_1 gpc3996 (
      {stage2_17[121]},
      {stage3_17[70]}
   );
   gpc1_1 gpc3997 (
      {stage2_17[122]},
      {stage3_17[71]}
   );
   gpc1_1 gpc3998 (
      {stage2_17[123]},
      {stage3_17[72]}
   );
   gpc1_1 gpc3999 (
      {stage2_17[124]},
      {stage3_17[73]}
   );
   gpc1_1 gpc4000 (
      {stage2_17[125]},
      {stage3_17[74]}
   );
   gpc1_1 gpc4001 (
      {stage2_17[126]},
      {stage3_17[75]}
   );
   gpc1_1 gpc4002 (
      {stage2_17[127]},
      {stage3_17[76]}
   );
   gpc1_1 gpc4003 (
      {stage2_19[64]},
      {stage3_19[36]}
   );
   gpc1_1 gpc4004 (
      {stage2_19[65]},
      {stage3_19[37]}
   );
   gpc1_1 gpc4005 (
      {stage2_19[66]},
      {stage3_19[38]}
   );
   gpc1_1 gpc4006 (
      {stage2_19[67]},
      {stage3_19[39]}
   );
   gpc1_1 gpc4007 (
      {stage2_19[68]},
      {stage3_19[40]}
   );
   gpc1_1 gpc4008 (
      {stage2_19[69]},
      {stage3_19[41]}
   );
   gpc1_1 gpc4009 (
      {stage2_19[70]},
      {stage3_19[42]}
   );
   gpc1_1 gpc4010 (
      {stage2_19[71]},
      {stage3_19[43]}
   );
   gpc1_1 gpc4011 (
      {stage2_19[72]},
      {stage3_19[44]}
   );
   gpc1_1 gpc4012 (
      {stage2_19[73]},
      {stage3_19[45]}
   );
   gpc1_1 gpc4013 (
      {stage2_19[74]},
      {stage3_19[46]}
   );
   gpc1_1 gpc4014 (
      {stage2_19[75]},
      {stage3_19[47]}
   );
   gpc1_1 gpc4015 (
      {stage2_19[76]},
      {stage3_19[48]}
   );
   gpc1_1 gpc4016 (
      {stage2_19[77]},
      {stage3_19[49]}
   );
   gpc1_1 gpc4017 (
      {stage2_19[78]},
      {stage3_19[50]}
   );
   gpc1_1 gpc4018 (
      {stage2_19[79]},
      {stage3_19[51]}
   );
   gpc1_1 gpc4019 (
      {stage2_19[80]},
      {stage3_19[52]}
   );
   gpc1_1 gpc4020 (
      {stage2_19[81]},
      {stage3_19[53]}
   );
   gpc1_1 gpc4021 (
      {stage2_19[82]},
      {stage3_19[54]}
   );
   gpc1_1 gpc4022 (
      {stage2_19[83]},
      {stage3_19[55]}
   );
   gpc1_1 gpc4023 (
      {stage2_19[84]},
      {stage3_19[56]}
   );
   gpc1_1 gpc4024 (
      {stage2_19[85]},
      {stage3_19[57]}
   );
   gpc1_1 gpc4025 (
      {stage2_19[86]},
      {stage3_19[58]}
   );
   gpc1_1 gpc4026 (
      {stage2_19[87]},
      {stage3_19[59]}
   );
   gpc1_1 gpc4027 (
      {stage2_19[88]},
      {stage3_19[60]}
   );
   gpc1_1 gpc4028 (
      {stage2_19[89]},
      {stage3_19[61]}
   );
   gpc1_1 gpc4029 (
      {stage2_19[90]},
      {stage3_19[62]}
   );
   gpc1_1 gpc4030 (
      {stage2_19[91]},
      {stage3_19[63]}
   );
   gpc1_1 gpc4031 (
      {stage2_19[92]},
      {stage3_19[64]}
   );
   gpc1_1 gpc4032 (
      {stage2_19[93]},
      {stage3_19[65]}
   );
   gpc1_1 gpc4033 (
      {stage2_19[94]},
      {stage3_19[66]}
   );
   gpc1_1 gpc4034 (
      {stage2_19[95]},
      {stage3_19[67]}
   );
   gpc1_1 gpc4035 (
      {stage2_19[96]},
      {stage3_19[68]}
   );
   gpc1_1 gpc4036 (
      {stage2_19[97]},
      {stage3_19[69]}
   );
   gpc1_1 gpc4037 (
      {stage2_21[96]},
      {stage3_21[34]}
   );
   gpc1_1 gpc4038 (
      {stage2_21[97]},
      {stage3_21[35]}
   );
   gpc1_1 gpc4039 (
      {stage2_21[98]},
      {stage3_21[36]}
   );
   gpc1_1 gpc4040 (
      {stage2_21[99]},
      {stage3_21[37]}
   );
   gpc1_1 gpc4041 (
      {stage2_21[100]},
      {stage3_21[38]}
   );
   gpc1_1 gpc4042 (
      {stage2_21[101]},
      {stage3_21[39]}
   );
   gpc1_1 gpc4043 (
      {stage2_21[102]},
      {stage3_21[40]}
   );
   gpc1_1 gpc4044 (
      {stage2_21[103]},
      {stage3_21[41]}
   );
   gpc1_1 gpc4045 (
      {stage2_21[104]},
      {stage3_21[42]}
   );
   gpc1_1 gpc4046 (
      {stage2_21[105]},
      {stage3_21[43]}
   );
   gpc1_1 gpc4047 (
      {stage2_21[106]},
      {stage3_21[44]}
   );
   gpc1_1 gpc4048 (
      {stage2_21[107]},
      {stage3_21[45]}
   );
   gpc1_1 gpc4049 (
      {stage2_21[108]},
      {stage3_21[46]}
   );
   gpc1_1 gpc4050 (
      {stage2_21[109]},
      {stage3_21[47]}
   );
   gpc1_1 gpc4051 (
      {stage2_21[110]},
      {stage3_21[48]}
   );
   gpc1_1 gpc4052 (
      {stage2_21[111]},
      {stage3_21[49]}
   );
   gpc1_1 gpc4053 (
      {stage2_21[112]},
      {stage3_21[50]}
   );
   gpc1_1 gpc4054 (
      {stage2_21[113]},
      {stage3_21[51]}
   );
   gpc1_1 gpc4055 (
      {stage2_21[114]},
      {stage3_21[52]}
   );
   gpc1_1 gpc4056 (
      {stage2_21[115]},
      {stage3_21[53]}
   );
   gpc1_1 gpc4057 (
      {stage2_21[116]},
      {stage3_21[54]}
   );
   gpc1_1 gpc4058 (
      {stage2_21[117]},
      {stage3_21[55]}
   );
   gpc1_1 gpc4059 (
      {stage2_21[118]},
      {stage3_21[56]}
   );
   gpc1_1 gpc4060 (
      {stage2_21[119]},
      {stage3_21[57]}
   );
   gpc1_1 gpc4061 (
      {stage2_21[120]},
      {stage3_21[58]}
   );
   gpc1_1 gpc4062 (
      {stage2_21[121]},
      {stage3_21[59]}
   );
   gpc1_1 gpc4063 (
      {stage2_21[122]},
      {stage3_21[60]}
   );
   gpc1_1 gpc4064 (
      {stage2_21[123]},
      {stage3_21[61]}
   );
   gpc1_1 gpc4065 (
      {stage2_21[124]},
      {stage3_21[62]}
   );
   gpc1_1 gpc4066 (
      {stage2_22[87]},
      {stage3_22[43]}
   );
   gpc1_1 gpc4067 (
      {stage2_22[88]},
      {stage3_22[44]}
   );
   gpc1_1 gpc4068 (
      {stage2_22[89]},
      {stage3_22[45]}
   );
   gpc1_1 gpc4069 (
      {stage2_22[90]},
      {stage3_22[46]}
   );
   gpc1_1 gpc4070 (
      {stage2_22[91]},
      {stage3_22[47]}
   );
   gpc1_1 gpc4071 (
      {stage2_22[92]},
      {stage3_22[48]}
   );
   gpc1_1 gpc4072 (
      {stage2_22[93]},
      {stage3_22[49]}
   );
   gpc1_1 gpc4073 (
      {stage2_22[94]},
      {stage3_22[50]}
   );
   gpc1_1 gpc4074 (
      {stage2_24[66]},
      {stage3_24[37]}
   );
   gpc1_1 gpc4075 (
      {stage2_24[67]},
      {stage3_24[38]}
   );
   gpc1_1 gpc4076 (
      {stage2_24[68]},
      {stage3_24[39]}
   );
   gpc1_1 gpc4077 (
      {stage2_24[69]},
      {stage3_24[40]}
   );
   gpc1_1 gpc4078 (
      {stage2_24[70]},
      {stage3_24[41]}
   );
   gpc1_1 gpc4079 (
      {stage2_24[71]},
      {stage3_24[42]}
   );
   gpc1_1 gpc4080 (
      {stage2_24[72]},
      {stage3_24[43]}
   );
   gpc1_1 gpc4081 (
      {stage2_24[73]},
      {stage3_24[44]}
   );
   gpc1_1 gpc4082 (
      {stage2_24[74]},
      {stage3_24[45]}
   );
   gpc1_1 gpc4083 (
      {stage2_24[75]},
      {stage3_24[46]}
   );
   gpc1_1 gpc4084 (
      {stage2_24[76]},
      {stage3_24[47]}
   );
   gpc1_1 gpc4085 (
      {stage2_24[77]},
      {stage3_24[48]}
   );
   gpc1_1 gpc4086 (
      {stage2_24[78]},
      {stage3_24[49]}
   );
   gpc1_1 gpc4087 (
      {stage2_24[79]},
      {stage3_24[50]}
   );
   gpc1_1 gpc4088 (
      {stage2_24[80]},
      {stage3_24[51]}
   );
   gpc1_1 gpc4089 (
      {stage2_24[81]},
      {stage3_24[52]}
   );
   gpc1_1 gpc4090 (
      {stage2_24[82]},
      {stage3_24[53]}
   );
   gpc1_1 gpc4091 (
      {stage2_24[83]},
      {stage3_24[54]}
   );
   gpc1_1 gpc4092 (
      {stage2_24[84]},
      {stage3_24[55]}
   );
   gpc1_1 gpc4093 (
      {stage2_24[85]},
      {stage3_24[56]}
   );
   gpc1_1 gpc4094 (
      {stage2_24[86]},
      {stage3_24[57]}
   );
   gpc1_1 gpc4095 (
      {stage2_24[87]},
      {stage3_24[58]}
   );
   gpc1_1 gpc4096 (
      {stage2_24[88]},
      {stage3_24[59]}
   );
   gpc1_1 gpc4097 (
      {stage2_24[89]},
      {stage3_24[60]}
   );
   gpc1_1 gpc4098 (
      {stage2_25[84]},
      {stage3_25[30]}
   );
   gpc1_1 gpc4099 (
      {stage2_25[85]},
      {stage3_25[31]}
   );
   gpc1_1 gpc4100 (
      {stage2_25[86]},
      {stage3_25[32]}
   );
   gpc1_1 gpc4101 (
      {stage2_25[87]},
      {stage3_25[33]}
   );
   gpc1_1 gpc4102 (
      {stage2_25[88]},
      {stage3_25[34]}
   );
   gpc1_1 gpc4103 (
      {stage2_25[89]},
      {stage3_25[35]}
   );
   gpc1_1 gpc4104 (
      {stage2_25[90]},
      {stage3_25[36]}
   );
   gpc1_1 gpc4105 (
      {stage2_25[91]},
      {stage3_25[37]}
   );
   gpc1_1 gpc4106 (
      {stage2_25[92]},
      {stage3_25[38]}
   );
   gpc1_1 gpc4107 (
      {stage2_25[93]},
      {stage3_25[39]}
   );
   gpc1_1 gpc4108 (
      {stage2_25[94]},
      {stage3_25[40]}
   );
   gpc1_1 gpc4109 (
      {stage2_25[95]},
      {stage3_25[41]}
   );
   gpc1_1 gpc4110 (
      {stage2_25[96]},
      {stage3_25[42]}
   );
   gpc1_1 gpc4111 (
      {stage2_25[97]},
      {stage3_25[43]}
   );
   gpc1_1 gpc4112 (
      {stage2_25[98]},
      {stage3_25[44]}
   );
   gpc1_1 gpc4113 (
      {stage2_25[99]},
      {stage3_25[45]}
   );
   gpc1_1 gpc4114 (
      {stage2_25[100]},
      {stage3_25[46]}
   );
   gpc1_1 gpc4115 (
      {stage2_25[101]},
      {stage3_25[47]}
   );
   gpc1_1 gpc4116 (
      {stage2_25[102]},
      {stage3_25[48]}
   );
   gpc1_1 gpc4117 (
      {stage2_26[87]},
      {stage3_26[38]}
   );
   gpc1_1 gpc4118 (
      {stage2_26[88]},
      {stage3_26[39]}
   );
   gpc1_1 gpc4119 (
      {stage2_26[89]},
      {stage3_26[40]}
   );
   gpc1_1 gpc4120 (
      {stage2_26[90]},
      {stage3_26[41]}
   );
   gpc1_1 gpc4121 (
      {stage2_26[91]},
      {stage3_26[42]}
   );
   gpc1_1 gpc4122 (
      {stage2_26[92]},
      {stage3_26[43]}
   );
   gpc1_1 gpc4123 (
      {stage2_26[93]},
      {stage3_26[44]}
   );
   gpc1_1 gpc4124 (
      {stage2_26[94]},
      {stage3_26[45]}
   );
   gpc1_1 gpc4125 (
      {stage2_26[95]},
      {stage3_26[46]}
   );
   gpc1_1 gpc4126 (
      {stage2_26[96]},
      {stage3_26[47]}
   );
   gpc1_1 gpc4127 (
      {stage2_26[97]},
      {stage3_26[48]}
   );
   gpc1_1 gpc4128 (
      {stage2_26[98]},
      {stage3_26[49]}
   );
   gpc1_1 gpc4129 (
      {stage2_26[99]},
      {stage3_26[50]}
   );
   gpc1_1 gpc4130 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc4131 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc4132 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc4133 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc4134 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc4135 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc4136 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc4137 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc4138 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc4139 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc4140 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc4141 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc4142 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc4143 (
      {stage2_28[133]},
      {stage3_28[36]}
   );
   gpc1_1 gpc4144 (
      {stage2_28[134]},
      {stage3_28[37]}
   );
   gpc1_1 gpc4145 (
      {stage2_28[135]},
      {stage3_28[38]}
   );
   gpc1_1 gpc4146 (
      {stage2_28[136]},
      {stage3_28[39]}
   );
   gpc1_1 gpc4147 (
      {stage2_28[137]},
      {stage3_28[40]}
   );
   gpc1_1 gpc4148 (
      {stage2_28[138]},
      {stage3_28[41]}
   );
   gpc1_1 gpc4149 (
      {stage2_28[139]},
      {stage3_28[42]}
   );
   gpc1_1 gpc4150 (
      {stage2_28[140]},
      {stage3_28[43]}
   );
   gpc1_1 gpc4151 (
      {stage2_28[141]},
      {stage3_28[44]}
   );
   gpc1_1 gpc4152 (
      {stage2_28[142]},
      {stage3_28[45]}
   );
   gpc1_1 gpc4153 (
      {stage2_28[143]},
      {stage3_28[46]}
   );
   gpc1_1 gpc4154 (
      {stage2_28[144]},
      {stage3_28[47]}
   );
   gpc1_1 gpc4155 (
      {stage2_28[145]},
      {stage3_28[48]}
   );
   gpc1_1 gpc4156 (
      {stage2_28[146]},
      {stage3_28[49]}
   );
   gpc1_1 gpc4157 (
      {stage2_28[147]},
      {stage3_28[50]}
   );
   gpc1_1 gpc4158 (
      {stage2_28[148]},
      {stage3_28[51]}
   );
   gpc1_1 gpc4159 (
      {stage2_28[149]},
      {stage3_28[52]}
   );
   gpc1_1 gpc4160 (
      {stage2_28[150]},
      {stage3_28[53]}
   );
   gpc1_1 gpc4161 (
      {stage2_28[151]},
      {stage3_28[54]}
   );
   gpc1_1 gpc4162 (
      {stage2_28[152]},
      {stage3_28[55]}
   );
   gpc1_1 gpc4163 (
      {stage2_28[153]},
      {stage3_28[56]}
   );
   gpc1_1 gpc4164 (
      {stage2_28[154]},
      {stage3_28[57]}
   );
   gpc1_1 gpc4165 (
      {stage2_28[155]},
      {stage3_28[58]}
   );
   gpc1_1 gpc4166 (
      {stage2_28[156]},
      {stage3_28[59]}
   );
   gpc1_1 gpc4167 (
      {stage2_28[157]},
      {stage3_28[60]}
   );
   gpc1_1 gpc4168 (
      {stage2_28[158]},
      {stage3_28[61]}
   );
   gpc1_1 gpc4169 (
      {stage2_28[159]},
      {stage3_28[62]}
   );
   gpc1_1 gpc4170 (
      {stage2_28[160]},
      {stage3_28[63]}
   );
   gpc1_1 gpc4171 (
      {stage2_28[161]},
      {stage3_28[64]}
   );
   gpc1_1 gpc4172 (
      {stage2_28[162]},
      {stage3_28[65]}
   );
   gpc1_1 gpc4173 (
      {stage2_28[163]},
      {stage3_28[66]}
   );
   gpc1_1 gpc4174 (
      {stage2_28[164]},
      {stage3_28[67]}
   );
   gpc1_1 gpc4175 (
      {stage2_28[165]},
      {stage3_28[68]}
   );
   gpc1_1 gpc4176 (
      {stage2_28[166]},
      {stage3_28[69]}
   );
   gpc1_1 gpc4177 (
      {stage2_28[167]},
      {stage3_28[70]}
   );
   gpc1_1 gpc4178 (
      {stage2_28[168]},
      {stage3_28[71]}
   );
   gpc1_1 gpc4179 (
      {stage2_28[169]},
      {stage3_28[72]}
   );
   gpc1_1 gpc4180 (
      {stage2_28[170]},
      {stage3_28[73]}
   );
   gpc1_1 gpc4181 (
      {stage2_29[127]},
      {stage3_29[42]}
   );
   gpc1_1 gpc4182 (
      {stage2_29[128]},
      {stage3_29[43]}
   );
   gpc1_1 gpc4183 (
      {stage2_29[129]},
      {stage3_29[44]}
   );
   gpc1_1 gpc4184 (
      {stage2_29[130]},
      {stage3_29[45]}
   );
   gpc1_1 gpc4185 (
      {stage2_29[131]},
      {stage3_29[46]}
   );
   gpc1_1 gpc4186 (
      {stage2_29[132]},
      {stage3_29[47]}
   );
   gpc1_1 gpc4187 (
      {stage2_29[133]},
      {stage3_29[48]}
   );
   gpc1_1 gpc4188 (
      {stage2_29[134]},
      {stage3_29[49]}
   );
   gpc1_1 gpc4189 (
      {stage2_29[135]},
      {stage3_29[50]}
   );
   gpc1_1 gpc4190 (
      {stage2_29[136]},
      {stage3_29[51]}
   );
   gpc1_1 gpc4191 (
      {stage2_29[137]},
      {stage3_29[52]}
   );
   gpc1_1 gpc4192 (
      {stage2_29[138]},
      {stage3_29[53]}
   );
   gpc1_1 gpc4193 (
      {stage2_29[139]},
      {stage3_29[54]}
   );
   gpc1_1 gpc4194 (
      {stage2_29[140]},
      {stage3_29[55]}
   );
   gpc1_1 gpc4195 (
      {stage2_29[141]},
      {stage3_29[56]}
   );
   gpc1_1 gpc4196 (
      {stage2_29[142]},
      {stage3_29[57]}
   );
   gpc1_1 gpc4197 (
      {stage2_30[66]},
      {stage3_30[45]}
   );
   gpc1_1 gpc4198 (
      {stage2_30[67]},
      {stage3_30[46]}
   );
   gpc1_1 gpc4199 (
      {stage2_30[68]},
      {stage3_30[47]}
   );
   gpc1_1 gpc4200 (
      {stage2_30[69]},
      {stage3_30[48]}
   );
   gpc1_1 gpc4201 (
      {stage2_30[70]},
      {stage3_30[49]}
   );
   gpc1_1 gpc4202 (
      {stage2_30[71]},
      {stage3_30[50]}
   );
   gpc1_1 gpc4203 (
      {stage2_30[72]},
      {stage3_30[51]}
   );
   gpc1_1 gpc4204 (
      {stage2_30[73]},
      {stage3_30[52]}
   );
   gpc1_1 gpc4205 (
      {stage2_30[74]},
      {stage3_30[53]}
   );
   gpc1_1 gpc4206 (
      {stage2_30[75]},
      {stage3_30[54]}
   );
   gpc1_1 gpc4207 (
      {stage2_30[76]},
      {stage3_30[55]}
   );
   gpc1_1 gpc4208 (
      {stage2_30[77]},
      {stage3_30[56]}
   );
   gpc1_1 gpc4209 (
      {stage2_30[78]},
      {stage3_30[57]}
   );
   gpc1_1 gpc4210 (
      {stage2_30[79]},
      {stage3_30[58]}
   );
   gpc1_1 gpc4211 (
      {stage2_30[80]},
      {stage3_30[59]}
   );
   gpc1_1 gpc4212 (
      {stage2_30[81]},
      {stage3_30[60]}
   );
   gpc1_1 gpc4213 (
      {stage2_30[82]},
      {stage3_30[61]}
   );
   gpc1_1 gpc4214 (
      {stage2_30[83]},
      {stage3_30[62]}
   );
   gpc1_1 gpc4215 (
      {stage2_30[84]},
      {stage3_30[63]}
   );
   gpc1_1 gpc4216 (
      {stage2_30[85]},
      {stage3_30[64]}
   );
   gpc1_1 gpc4217 (
      {stage2_30[86]},
      {stage3_30[65]}
   );
   gpc1_1 gpc4218 (
      {stage2_30[87]},
      {stage3_30[66]}
   );
   gpc1_1 gpc4219 (
      {stage2_30[88]},
      {stage3_30[67]}
   );
   gpc1_1 gpc4220 (
      {stage2_30[89]},
      {stage3_30[68]}
   );
   gpc1_1 gpc4221 (
      {stage2_30[90]},
      {stage3_30[69]}
   );
   gpc1_1 gpc4222 (
      {stage2_30[91]},
      {stage3_30[70]}
   );
   gpc1_1 gpc4223 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc4224 (
      {stage2_31[84]},
      {stage3_31[40]}
   );
   gpc1_1 gpc4225 (
      {stage2_31[85]},
      {stage3_31[41]}
   );
   gpc1_1 gpc4226 (
      {stage2_31[86]},
      {stage3_31[42]}
   );
   gpc1_1 gpc4227 (
      {stage2_31[87]},
      {stage3_31[43]}
   );
   gpc1_1 gpc4228 (
      {stage2_31[88]},
      {stage3_31[44]}
   );
   gpc1_1 gpc4229 (
      {stage2_31[89]},
      {stage3_31[45]}
   );
   gpc1_1 gpc4230 (
      {stage2_31[90]},
      {stage3_31[46]}
   );
   gpc1_1 gpc4231 (
      {stage2_31[91]},
      {stage3_31[47]}
   );
   gpc1_1 gpc4232 (
      {stage2_31[92]},
      {stage3_31[48]}
   );
   gpc1_1 gpc4233 (
      {stage2_31[93]},
      {stage3_31[49]}
   );
   gpc1_1 gpc4234 (
      {stage2_31[94]},
      {stage3_31[50]}
   );
   gpc1_1 gpc4235 (
      {stage2_31[95]},
      {stage3_31[51]}
   );
   gpc1_1 gpc4236 (
      {stage2_31[96]},
      {stage3_31[52]}
   );
   gpc1_1 gpc4237 (
      {stage2_31[97]},
      {stage3_31[53]}
   );
   gpc1_1 gpc4238 (
      {stage2_31[98]},
      {stage3_31[54]}
   );
   gpc1_1 gpc4239 (
      {stage2_31[99]},
      {stage3_31[55]}
   );
   gpc1_1 gpc4240 (
      {stage2_31[100]},
      {stage3_31[56]}
   );
   gpc1_1 gpc4241 (
      {stage2_31[101]},
      {stage3_31[57]}
   );
   gpc1_1 gpc4242 (
      {stage2_32[46]},
      {stage3_32[30]}
   );
   gpc1_1 gpc4243 (
      {stage2_32[47]},
      {stage3_32[31]}
   );
   gpc1_1 gpc4244 (
      {stage2_32[48]},
      {stage3_32[32]}
   );
   gpc1_1 gpc4245 (
      {stage2_32[49]},
      {stage3_32[33]}
   );
   gpc1_1 gpc4246 (
      {stage2_32[50]},
      {stage3_32[34]}
   );
   gpc1_1 gpc4247 (
      {stage2_32[51]},
      {stage3_32[35]}
   );
   gpc1_1 gpc4248 (
      {stage2_32[52]},
      {stage3_32[36]}
   );
   gpc1_1 gpc4249 (
      {stage2_32[53]},
      {stage3_32[37]}
   );
   gpc1_1 gpc4250 (
      {stage2_32[54]},
      {stage3_32[38]}
   );
   gpc1_1 gpc4251 (
      {stage2_32[55]},
      {stage3_32[39]}
   );
   gpc1_1 gpc4252 (
      {stage2_32[56]},
      {stage3_32[40]}
   );
   gpc1_1 gpc4253 (
      {stage2_32[57]},
      {stage3_32[41]}
   );
   gpc1_1 gpc4254 (
      {stage2_32[58]},
      {stage3_32[42]}
   );
   gpc1_1 gpc4255 (
      {stage2_32[59]},
      {stage3_32[43]}
   );
   gpc1_1 gpc4256 (
      {stage2_32[60]},
      {stage3_32[44]}
   );
   gpc1_1 gpc4257 (
      {stage2_32[61]},
      {stage3_32[45]}
   );
   gpc1_1 gpc4258 (
      {stage2_32[62]},
      {stage3_32[46]}
   );
   gpc1_1 gpc4259 (
      {stage2_32[63]},
      {stage3_32[47]}
   );
   gpc1_1 gpc4260 (
      {stage2_32[64]},
      {stage3_32[48]}
   );
   gpc1_1 gpc4261 (
      {stage2_32[65]},
      {stage3_32[49]}
   );
   gpc1_1 gpc4262 (
      {stage2_32[66]},
      {stage3_32[50]}
   );
   gpc1_1 gpc4263 (
      {stage2_32[67]},
      {stage3_32[51]}
   );
   gpc1_1 gpc4264 (
      {stage2_32[68]},
      {stage3_32[52]}
   );
   gpc1_1 gpc4265 (
      {stage2_32[69]},
      {stage3_32[53]}
   );
   gpc1_1 gpc4266 (
      {stage2_32[70]},
      {stage3_32[54]}
   );
   gpc1_1 gpc4267 (
      {stage2_32[71]},
      {stage3_32[55]}
   );
   gpc1_1 gpc4268 (
      {stage2_32[72]},
      {stage3_32[56]}
   );
   gpc1_1 gpc4269 (
      {stage2_32[73]},
      {stage3_32[57]}
   );
   gpc1_1 gpc4270 (
      {stage2_33[57]},
      {stage3_33[24]}
   );
   gpc1_1 gpc4271 (
      {stage2_33[58]},
      {stage3_33[25]}
   );
   gpc1_1 gpc4272 (
      {stage2_33[59]},
      {stage3_33[26]}
   );
   gpc1_1 gpc4273 (
      {stage2_34[24]},
      {stage3_34[16]}
   );
   gpc1_1 gpc4274 (
      {stage2_34[25]},
      {stage3_34[17]}
   );
   gpc1_1 gpc4275 (
      {stage2_34[26]},
      {stage3_34[18]}
   );
   gpc1_1 gpc4276 (
      {stage2_34[27]},
      {stage3_34[19]}
   );
   gpc1_1 gpc4277 (
      {stage2_34[28]},
      {stage3_34[20]}
   );
   gpc1_1 gpc4278 (
      {stage2_34[29]},
      {stage3_34[21]}
   );
   gpc1_1 gpc4279 (
      {stage2_34[30]},
      {stage3_34[22]}
   );
   gpc1_1 gpc4280 (
      {stage2_34[31]},
      {stage3_34[23]}
   );
   gpc1_1 gpc4281 (
      {stage2_34[32]},
      {stage3_34[24]}
   );
   gpc1_1 gpc4282 (
      {stage2_34[33]},
      {stage3_34[25]}
   );
   gpc1_1 gpc4283 (
      {stage2_34[34]},
      {stage3_34[26]}
   );
   gpc606_5 gpc4284 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc4285 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc4286 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4287 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc4288 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc4289 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc4290 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage4_6[4],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc4291 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[5],stage4_5[7]}
   );
   gpc606_5 gpc4292 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[1],stage4_7[1],stage4_6[6],stage4_5[8]}
   );
   gpc606_5 gpc4293 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[2],stage4_7[2],stage4_6[7],stage4_5[9]}
   );
   gpc606_5 gpc4294 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[3],stage4_7[3],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc4295 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[24]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[4],stage4_7[4],stage4_6[9]}
   );
   gpc615_5 gpc4296 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[25]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[5],stage4_7[5],stage4_6[10]}
   );
   gpc615_5 gpc4297 (
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14]},
      {stage3_7[26]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[6],stage4_7[6],stage4_6[11]}
   );
   gpc615_5 gpc4298 (
      {stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19]},
      {stage3_7[27]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[7],stage4_7[7],stage4_6[12]}
   );
   gpc615_5 gpc4299 (
      {stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_7[28]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[8],stage4_7[8],stage4_6[13]}
   );
   gpc615_5 gpc4300 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage3_7[29]},
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], stage3_8[35]},
      {stage4_10[5],stage4_9[9],stage4_8[9],stage4_7[9],stage4_6[14]}
   );
   gpc615_5 gpc4301 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[36]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[6],stage4_9[10],stage4_8[10],stage4_7[10]}
   );
   gpc615_5 gpc4302 (
      {stage3_7[35], stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39]},
      {stage3_8[37]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[7],stage4_9[11],stage4_8[11],stage4_7[11]}
   );
   gpc615_5 gpc4303 (
      {stage3_7[40], stage3_7[41], stage3_7[42], stage3_7[43], stage3_7[44]},
      {stage3_8[38]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[8],stage4_9[12],stage4_8[12],stage4_7[12]}
   );
   gpc117_4 gpc4304 (
      {stage3_8[39], stage3_8[40], stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45]},
      {stage3_9[18]},
      {stage3_10[0]},
      {stage4_11[3],stage4_10[9],stage4_9[13],stage4_8[13]}
   );
   gpc117_4 gpc4305 (
      {stage3_8[46], stage3_8[47], stage3_8[48], stage3_8[49], stage3_8[50], stage3_8[51], stage3_8[52]},
      {stage3_9[19]},
      {stage3_10[1]},
      {stage4_11[4],stage4_10[10],stage4_9[14],stage4_8[14]}
   );
   gpc606_5 gpc4306 (
      {stage3_8[53], stage3_8[54], stage3_8[55], stage3_8[56], stage3_8[57], stage3_8[58]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[5],stage4_10[11],stage4_9[15],stage4_8[15]}
   );
   gpc606_5 gpc4307 (
      {stage3_8[59], stage3_8[60], stage3_8[61], stage3_8[62], stage3_8[63], stage3_8[64]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[6],stage4_10[12],stage4_9[16],stage4_8[16]}
   );
   gpc615_5 gpc4308 (
      {stage3_8[65], stage3_8[66], stage3_8[67], stage3_8[68], stage3_8[69]},
      {stage3_9[20]},
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage4_12[2],stage4_11[7],stage4_10[13],stage4_9[17],stage4_8[17]}
   );
   gpc615_5 gpc4309 (
      {stage3_8[70], stage3_8[71], stage3_8[72], stage3_8[73], stage3_8[74]},
      {stage3_9[21]},
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage4_12[3],stage4_11[8],stage4_10[14],stage4_9[18],stage4_8[18]}
   );
   gpc615_5 gpc4310 (
      {stage3_8[75], stage3_8[76], stage3_8[77], stage3_8[78], stage3_8[79]},
      {stage3_9[22]},
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage4_12[4],stage4_11[9],stage4_10[15],stage4_9[19],stage4_8[19]}
   );
   gpc615_5 gpc4311 (
      {stage3_8[80], stage3_8[81], stage3_8[82], stage3_8[83], stage3_8[84]},
      {stage3_9[23]},
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage4_12[5],stage4_11[10],stage4_10[16],stage4_9[20],stage4_8[20]}
   );
   gpc606_5 gpc4312 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[6],stage4_11[11],stage4_10[17],stage4_9[21]}
   );
   gpc1163_5 gpc4313 (
      {stage3_11[6], stage3_11[7], stage3_11[8]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[7],stage4_11[12]}
   );
   gpc1163_5 gpc4314 (
      {stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_13[1]},
      {stage3_14[1]},
      {stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[8],stage4_11[13]}
   );
   gpc1163_5 gpc4315 (
      {stage3_11[12], stage3_11[13], stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_13[2]},
      {stage3_14[2]},
      {stage4_15[2],stage4_14[2],stage4_13[3],stage4_12[9],stage4_11[14]}
   );
   gpc1163_5 gpc4316 (
      {stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[3]},
      {stage3_14[3]},
      {stage4_15[3],stage4_14[3],stage4_13[4],stage4_12[10],stage4_11[15]}
   );
   gpc1163_5 gpc4317 (
      {stage3_11[18], stage3_11[19], stage3_11[20]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_13[4]},
      {stage3_14[4]},
      {stage4_15[4],stage4_14[4],stage4_13[5],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc4318 (
      {stage3_11[21], stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25]},
      {stage3_12[30]},
      {stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage4_15[5],stage4_14[5],stage4_13[6],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc4319 (
      {stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29], stage3_11[30]},
      {stage3_12[31]},
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16]},
      {stage4_15[6],stage4_14[6],stage4_13[7],stage4_12[13],stage4_11[18]}
   );
   gpc606_5 gpc4320 (
      {stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37]},
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage4_16[0],stage4_15[7],stage4_14[7],stage4_13[8],stage4_12[14]}
   );
   gpc606_5 gpc4321 (
      {stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[8],stage4_14[8],stage4_13[9]}
   );
   gpc606_5 gpc4322 (
      {stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[9],stage4_14[9],stage4_13[10]}
   );
   gpc615_5 gpc4323 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[10],stage4_14[10]}
   );
   gpc615_5 gpc4324 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[13]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[11],stage4_14[11]}
   );
   gpc615_5 gpc4325 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[14]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[12],stage4_14[12]}
   );
   gpc615_5 gpc4326 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[15]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[13],stage4_14[13]}
   );
   gpc615_5 gpc4327 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[16]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[14],stage4_14[14]}
   );
   gpc1163_5 gpc4328 (
      {stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[15]}
   );
   gpc615_5 gpc4329 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[36]},
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage4_19[1],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[16]}
   );
   gpc615_5 gpc4330 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[37]},
      {stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11], stage3_17[12]},
      {stage4_19[2],stage4_18[7],stage4_17[9],stage4_16[10],stage4_15[17]}
   );
   gpc615_5 gpc4331 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[38]},
      {stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage4_19[3],stage4_18[8],stage4_17[10],stage4_16[11],stage4_15[18]}
   );
   gpc615_5 gpc4332 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[39]},
      {stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23], stage3_17[24]},
      {stage4_19[4],stage4_18[9],stage4_17[11],stage4_16[12],stage4_15[19]}
   );
   gpc615_5 gpc4333 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[40]},
      {stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29], stage3_17[30]},
      {stage4_19[5],stage4_18[10],stage4_17[12],stage4_16[13],stage4_15[20]}
   );
   gpc615_5 gpc4334 (
      {stage3_15[45], stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49]},
      {stage3_16[41]},
      {stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35], stage3_17[36]},
      {stage4_19[6],stage4_18[11],stage4_17[13],stage4_16[14],stage4_15[21]}
   );
   gpc615_5 gpc4335 (
      {stage3_15[50], stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54]},
      {stage3_16[42]},
      {stage3_17[37], stage3_17[38], stage3_17[39], stage3_17[40], stage3_17[41], stage3_17[42]},
      {stage4_19[7],stage4_18[12],stage4_17[14],stage4_16[15],stage4_15[22]}
   );
   gpc606_5 gpc4336 (
      {stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46], stage3_16[47], stage3_16[48]},
      {stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage4_20[0],stage4_19[8],stage4_18[13],stage4_17[15],stage4_16[16]}
   );
   gpc606_5 gpc4337 (
      {stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52], stage3_16[53], stage3_16[54]},
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage4_20[1],stage4_19[9],stage4_18[14],stage4_17[16],stage4_16[17]}
   );
   gpc606_5 gpc4338 (
      {stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58], stage3_16[59], stage3_16[60]},
      {stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18]},
      {stage4_20[2],stage4_19[10],stage4_18[15],stage4_17[17],stage4_16[18]}
   );
   gpc606_5 gpc4339 (
      {stage3_16[61], stage3_16[62], stage3_16[63], stage3_16[64], stage3_16[65], stage3_16[66]},
      {stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24]},
      {stage4_20[3],stage4_19[11],stage4_18[16],stage4_17[18],stage4_16[19]}
   );
   gpc606_5 gpc4340 (
      {stage3_17[43], stage3_17[44], stage3_17[45], stage3_17[46], stage3_17[47], stage3_17[48]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[12],stage4_18[17],stage4_17[19]}
   );
   gpc606_5 gpc4341 (
      {stage3_17[49], stage3_17[50], stage3_17[51], stage3_17[52], stage3_17[53], stage3_17[54]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[13],stage4_18[18],stage4_17[20]}
   );
   gpc615_5 gpc4342 (
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[6],stage4_19[14]}
   );
   gpc615_5 gpc4343 (
      {stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21]},
      {stage3_20[1]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[3],stage4_20[7],stage4_19[15]}
   );
   gpc615_5 gpc4344 (
      {stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25], stage3_19[26]},
      {stage3_20[2]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[4],stage4_20[8],stage4_19[16]}
   );
   gpc615_5 gpc4345 (
      {stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30], stage3_19[31]},
      {stage3_20[3]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[5],stage4_20[9],stage4_19[17]}
   );
   gpc615_5 gpc4346 (
      {stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35], stage3_19[36]},
      {stage3_20[4]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[4],stage4_21[6],stage4_20[10],stage4_19[18]}
   );
   gpc615_5 gpc4347 (
      {stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40], stage3_19[41]},
      {stage3_20[5]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[5],stage4_21[7],stage4_20[11],stage4_19[19]}
   );
   gpc615_5 gpc4348 (
      {stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45], stage3_19[46]},
      {stage3_20[6]},
      {stage3_21[36], stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41]},
      {stage4_23[6],stage4_22[6],stage4_21[8],stage4_20[12],stage4_19[20]}
   );
   gpc615_5 gpc4349 (
      {stage3_19[47], stage3_19[48], stage3_19[49], stage3_19[50], stage3_19[51]},
      {stage3_20[7]},
      {stage3_21[42], stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47]},
      {stage4_23[7],stage4_22[7],stage4_21[9],stage4_20[13],stage4_19[21]}
   );
   gpc1325_5 gpc4350 (
      {stage3_19[52], stage3_19[53], stage3_19[54], stage3_19[55], stage3_19[56]},
      {stage3_20[8], stage3_20[9]},
      {stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_22[0]},
      {stage4_23[8],stage4_22[8],stage4_21[10],stage4_20[14],stage4_19[22]}
   );
   gpc1325_5 gpc4351 (
      {stage3_19[57], stage3_19[58], stage3_19[59], stage3_19[60], stage3_19[61]},
      {stage3_20[10], stage3_20[11]},
      {stage3_21[51], stage3_21[52], stage3_21[53]},
      {stage3_22[1]},
      {stage4_23[9],stage4_22[9],stage4_21[11],stage4_20[15],stage4_19[23]}
   );
   gpc606_5 gpc4352 (
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6], stage3_22[7]},
      {stage4_24[0],stage4_23[10],stage4_22[10],stage4_21[12],stage4_20[16]}
   );
   gpc606_5 gpc4353 (
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12], stage3_22[13]},
      {stage4_24[1],stage4_23[11],stage4_22[11],stage4_21[13],stage4_20[17]}
   );
   gpc606_5 gpc4354 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage4_24[2],stage4_23[12],stage4_22[12],stage4_21[14],stage4_20[18]}
   );
   gpc606_5 gpc4355 (
      {stage3_21[54], stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[3],stage4_23[13],stage4_22[13],stage4_21[15]}
   );
   gpc207_4 gpc4356 (
      {stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[1],stage4_24[4],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc4357 (
      {stage3_22[27], stage3_22[28], stage3_22[29], stage3_22[30], stage3_22[31]},
      {stage3_23[6]},
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7]},
      {stage4_26[0],stage4_25[2],stage4_24[5],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc4358 (
      {stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35], stage3_22[36]},
      {stage3_23[7]},
      {stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11], stage3_24[12], stage3_24[13]},
      {stage4_26[1],stage4_25[3],stage4_24[6],stage4_23[16],stage4_22[16]}
   );
   gpc606_5 gpc4359 (
      {stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12], stage3_23[13]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[4],stage4_24[7],stage4_23[17]}
   );
   gpc615_5 gpc4360 (
      {stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage3_24[14]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[5],stage4_24[8],stage4_23[18]}
   );
   gpc615_5 gpc4361 (
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage3_24[15]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[6],stage4_24[9],stage4_23[19]}
   );
   gpc615_5 gpc4362 (
      {stage3_23[24], stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28]},
      {stage3_24[16]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[5],stage4_25[7],stage4_24[10],stage4_23[20]}
   );
   gpc606_5 gpc4363 (
      {stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[4],stage4_26[6],stage4_25[8],stage4_24[11]}
   );
   gpc606_5 gpc4364 (
      {stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26], stage3_24[27], stage3_24[28]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[5],stage4_26[7],stage4_25[9],stage4_24[12]}
   );
   gpc606_5 gpc4365 (
      {stage3_24[29], stage3_24[30], stage3_24[31], stage3_24[32], stage3_24[33], stage3_24[34]},
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage4_28[2],stage4_27[6],stage4_26[8],stage4_25[10],stage4_24[13]}
   );
   gpc606_5 gpc4366 (
      {stage3_24[35], stage3_24[36], stage3_24[37], stage3_24[38], stage3_24[39], stage3_24[40]},
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage4_28[3],stage4_27[7],stage4_26[9],stage4_25[11],stage4_24[14]}
   );
   gpc606_5 gpc4367 (
      {stage3_24[41], stage3_24[42], stage3_24[43], stage3_24[44], stage3_24[45], stage3_24[46]},
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage4_28[4],stage4_27[8],stage4_26[10],stage4_25[12],stage4_24[15]}
   );
   gpc606_5 gpc4368 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[5],stage4_27[9],stage4_26[11],stage4_25[13]}
   );
   gpc606_5 gpc4369 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[6],stage4_27[10],stage4_26[12],stage4_25[14]}
   );
   gpc606_5 gpc4370 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[7],stage4_27[11],stage4_26[13],stage4_25[15]}
   );
   gpc615_5 gpc4371 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46]},
      {stage3_26[30]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[8],stage4_27[12],stage4_26[14],stage4_25[16]}
   );
   gpc615_5 gpc4372 (
      {stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[9],stage4_27[13],stage4_26[15]}
   );
   gpc615_5 gpc4373 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40]},
      {stage3_27[25]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[5],stage4_28[10],stage4_27[14],stage4_26[16]}
   );
   gpc615_5 gpc4374 (
      {stage3_26[41], stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45]},
      {stage3_27[26]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[6],stage4_28[11],stage4_27[15],stage4_26[17]}
   );
   gpc606_5 gpc4375 (
      {stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30], stage3_27[31], stage3_27[32]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[3],stage4_29[7],stage4_28[12],stage4_27[16]}
   );
   gpc615_5 gpc4376 (
      {stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_28[18]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[4],stage4_29[8],stage4_28[13],stage4_27[17]}
   );
   gpc615_5 gpc4377 (
      {stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_28[19]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[5],stage4_29[9],stage4_28[14],stage4_27[18]}
   );
   gpc615_5 gpc4378 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47]},
      {stage3_28[20]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[6],stage4_29[10],stage4_28[15],stage4_27[19]}
   );
   gpc606_5 gpc4379 (
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[4],stage4_30[7],stage4_29[11],stage4_28[16]}
   );
   gpc606_5 gpc4380 (
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[5],stage4_30[8],stage4_29[12],stage4_28[17]}
   );
   gpc606_5 gpc4381 (
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[6],stage4_30[9],stage4_29[13],stage4_28[18]}
   );
   gpc606_5 gpc4382 (
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[7],stage4_30[10],stage4_29[14],stage4_28[19]}
   );
   gpc606_5 gpc4383 (
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[8],stage4_30[11],stage4_29[15],stage4_28[20]}
   );
   gpc606_5 gpc4384 (
      {stage3_28[51], stage3_28[52], stage3_28[53], stage3_28[54], stage3_28[55], stage3_28[56]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[9],stage4_30[12],stage4_29[16],stage4_28[21]}
   );
   gpc606_5 gpc4385 (
      {stage3_28[57], stage3_28[58], stage3_28[59], stage3_28[60], stage3_28[61], stage3_28[62]},
      {stage3_30[36], stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41]},
      {stage4_32[6],stage4_31[10],stage4_30[13],stage4_29[17],stage4_28[22]}
   );
   gpc606_5 gpc4386 (
      {stage3_28[63], stage3_28[64], stage3_28[65], stage3_28[66], stage3_28[67], stage3_28[68]},
      {stage3_30[42], stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage4_32[7],stage4_31[11],stage4_30[14],stage4_29[18],stage4_28[23]}
   );
   gpc606_5 gpc4387 (
      {stage3_28[69], stage3_28[70], stage3_28[71], stage3_28[72], stage3_28[73], 1'b0},
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52], stage3_30[53]},
      {stage4_32[8],stage4_31[12],stage4_30[15],stage4_29[19],stage4_28[24]}
   );
   gpc606_5 gpc4388 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[9],stage4_31[13],stage4_30[16],stage4_29[20]}
   );
   gpc606_5 gpc4389 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[10],stage4_31[14],stage4_30[17],stage4_29[21]}
   );
   gpc606_5 gpc4390 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[11],stage4_31[15],stage4_30[18],stage4_29[22]}
   );
   gpc606_5 gpc4391 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23]},
      {stage4_33[3],stage4_32[12],stage4_31[16],stage4_30[19],stage4_29[23]}
   );
   gpc615_5 gpc4392 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52]},
      {stage3_30[54]},
      {stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage4_33[4],stage4_32[13],stage4_31[17],stage4_30[20],stage4_29[24]}
   );
   gpc615_5 gpc4393 (
      {stage3_29[53], stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57]},
      {stage3_30[55]},
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34], stage3_31[35]},
      {stage4_33[5],stage4_32[14],stage4_31[18],stage4_30[21],stage4_29[25]}
   );
   gpc606_5 gpc4394 (
      {stage3_30[56], stage3_30[57], stage3_30[58], stage3_30[59], stage3_30[60], stage3_30[61]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[6],stage4_32[15],stage4_31[19],stage4_30[22]}
   );
   gpc606_5 gpc4395 (
      {stage3_30[62], stage3_30[63], stage3_30[64], stage3_30[65], stage3_30[66], stage3_30[67]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[7],stage4_32[16],stage4_31[20],stage4_30[23]}
   );
   gpc615_5 gpc4396 (
      {stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39], stage3_31[40]},
      {stage3_32[12]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[8],stage4_32[17],stage4_31[21]}
   );
   gpc615_5 gpc4397 (
      {stage3_31[41], stage3_31[42], stage3_31[43], stage3_31[44], stage3_31[45]},
      {stage3_32[13]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[9],stage4_32[18],stage4_31[22]}
   );
   gpc615_5 gpc4398 (
      {stage3_31[46], stage3_31[47], stage3_31[48], stage3_31[49], stage3_31[50]},
      {stage3_32[14]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[10],stage4_32[19],stage4_31[23]}
   );
   gpc606_5 gpc4399 (
      {stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[11],stage4_32[20]}
   );
   gpc606_5 gpc4400 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[12],stage4_32[21]}
   );
   gpc606_5 gpc4401 (
      {stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[13],stage4_32[22]}
   );
   gpc606_5 gpc4402 (
      {stage3_32[33], stage3_32[34], stage3_32[35], stage3_32[36], stage3_32[37], stage3_32[38]},
      {stage3_34[18], stage3_34[19], stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[14],stage4_32[23]}
   );
   gpc606_5 gpc4403 (
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[15]}
   );
   gpc1_1 gpc4404 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc4405 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4406 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4407 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4408 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc4409 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc4410 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc4411 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc4412 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc4413 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc4414 (
      {stage3_0[10]},
      {stage4_0[10]}
   );
   gpc1_1 gpc4415 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4416 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4417 (
      {stage3_1[14]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4418 (
      {stage3_1[15]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4419 (
      {stage3_1[16]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4420 (
      {stage3_1[17]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4421 (
      {stage3_1[18]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4422 (
      {stage3_1[19]},
      {stage4_1[9]}
   );
   gpc1_1 gpc4423 (
      {stage3_1[20]},
      {stage4_1[10]}
   );
   gpc1_1 gpc4424 (
      {stage3_1[21]},
      {stage4_1[11]}
   );
   gpc1_1 gpc4425 (
      {stage3_1[22]},
      {stage4_1[12]}
   );
   gpc1_1 gpc4426 (
      {stage3_1[23]},
      {stage4_1[13]}
   );
   gpc1_1 gpc4427 (
      {stage3_1[24]},
      {stage4_1[14]}
   );
   gpc1_1 gpc4428 (
      {stage3_1[25]},
      {stage4_1[15]}
   );
   gpc1_1 gpc4429 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4430 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4431 (
      {stage3_2[32]},
      {stage4_2[9]}
   );
   gpc1_1 gpc4432 (
      {stage3_2[33]},
      {stage4_2[10]}
   );
   gpc1_1 gpc4433 (
      {stage3_2[34]},
      {stage4_2[11]}
   );
   gpc1_1 gpc4434 (
      {stage3_2[35]},
      {stage4_2[12]}
   );
   gpc1_1 gpc4435 (
      {stage3_3[12]},
      {stage4_3[7]}
   );
   gpc1_1 gpc4436 (
      {stage3_3[13]},
      {stage4_3[8]}
   );
   gpc1_1 gpc4437 (
      {stage3_3[14]},
      {stage4_3[9]}
   );
   gpc1_1 gpc4438 (
      {stage3_3[15]},
      {stage4_3[10]}
   );
   gpc1_1 gpc4439 (
      {stage3_3[16]},
      {stage4_3[11]}
   );
   gpc1_1 gpc4440 (
      {stage3_3[17]},
      {stage4_3[12]}
   );
   gpc1_1 gpc4441 (
      {stage3_3[18]},
      {stage4_3[13]}
   );
   gpc1_1 gpc4442 (
      {stage3_3[19]},
      {stage4_3[14]}
   );
   gpc1_1 gpc4443 (
      {stage3_3[20]},
      {stage4_3[15]}
   );
   gpc1_1 gpc4444 (
      {stage3_3[21]},
      {stage4_3[16]}
   );
   gpc1_1 gpc4445 (
      {stage3_3[22]},
      {stage4_3[17]}
   );
   gpc1_1 gpc4446 (
      {stage3_3[23]},
      {stage4_3[18]}
   );
   gpc1_1 gpc4447 (
      {stage3_3[24]},
      {stage4_3[19]}
   );
   gpc1_1 gpc4448 (
      {stage3_3[25]},
      {stage4_3[20]}
   );
   gpc1_1 gpc4449 (
      {stage3_3[26]},
      {stage4_3[21]}
   );
   gpc1_1 gpc4450 (
      {stage3_3[27]},
      {stage4_3[22]}
   );
   gpc1_1 gpc4451 (
      {stage3_4[30]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4452 (
      {stage3_4[31]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4453 (
      {stage3_4[32]},
      {stage4_4[9]}
   );
   gpc1_1 gpc4454 (
      {stage3_4[33]},
      {stage4_4[10]}
   );
   gpc1_1 gpc4455 (
      {stage3_4[34]},
      {stage4_4[11]}
   );
   gpc1_1 gpc4456 (
      {stage3_4[35]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4457 (
      {stage3_4[36]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4458 (
      {stage3_4[37]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4459 (
      {stage3_4[38]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4460 (
      {stage3_4[39]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4461 (
      {stage3_4[40]},
      {stage4_4[17]}
   );
   gpc1_1 gpc4462 (
      {stage3_4[41]},
      {stage4_4[18]}
   );
   gpc1_1 gpc4463 (
      {stage3_4[42]},
      {stage4_4[19]}
   );
   gpc1_1 gpc4464 (
      {stage3_4[43]},
      {stage4_4[20]}
   );
   gpc1_1 gpc4465 (
      {stage3_4[44]},
      {stage4_4[21]}
   );
   gpc1_1 gpc4466 (
      {stage3_4[45]},
      {stage4_4[22]}
   );
   gpc1_1 gpc4467 (
      {stage3_4[46]},
      {stage4_4[23]}
   );
   gpc1_1 gpc4468 (
      {stage3_5[24]},
      {stage4_5[11]}
   );
   gpc1_1 gpc4469 (
      {stage3_5[25]},
      {stage4_5[12]}
   );
   gpc1_1 gpc4470 (
      {stage3_5[26]},
      {stage4_5[13]}
   );
   gpc1_1 gpc4471 (
      {stage3_5[27]},
      {stage4_5[14]}
   );
   gpc1_1 gpc4472 (
      {stage3_5[28]},
      {stage4_5[15]}
   );
   gpc1_1 gpc4473 (
      {stage3_5[29]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4474 (
      {stage3_5[30]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4475 (
      {stage3_5[31]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4476 (
      {stage3_5[32]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4477 (
      {stage3_5[33]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4478 (
      {stage3_5[34]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4479 (
      {stage3_5[35]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4480 (
      {stage3_5[36]},
      {stage4_5[23]}
   );
   gpc1_1 gpc4481 (
      {stage3_5[37]},
      {stage4_5[24]}
   );
   gpc1_1 gpc4482 (
      {stage3_5[38]},
      {stage4_5[25]}
   );
   gpc1_1 gpc4483 (
      {stage3_5[39]},
      {stage4_5[26]}
   );
   gpc1_1 gpc4484 (
      {stage3_5[40]},
      {stage4_5[27]}
   );
   gpc1_1 gpc4485 (
      {stage3_5[41]},
      {stage4_5[28]}
   );
   gpc1_1 gpc4486 (
      {stage3_5[42]},
      {stage4_5[29]}
   );
   gpc1_1 gpc4487 (
      {stage3_5[43]},
      {stage4_5[30]}
   );
   gpc1_1 gpc4488 (
      {stage3_5[44]},
      {stage4_5[31]}
   );
   gpc1_1 gpc4489 (
      {stage3_5[45]},
      {stage4_5[32]}
   );
   gpc1_1 gpc4490 (
      {stage3_5[46]},
      {stage4_5[33]}
   );
   gpc1_1 gpc4491 (
      {stage3_5[47]},
      {stage4_5[34]}
   );
   gpc1_1 gpc4492 (
      {stage3_5[48]},
      {stage4_5[35]}
   );
   gpc1_1 gpc4493 (
      {stage3_5[49]},
      {stage4_5[36]}
   );
   gpc1_1 gpc4494 (
      {stage3_5[50]},
      {stage4_5[37]}
   );
   gpc1_1 gpc4495 (
      {stage3_5[51]},
      {stage4_5[38]}
   );
   gpc1_1 gpc4496 (
      {stage3_5[52]},
      {stage4_5[39]}
   );
   gpc1_1 gpc4497 (
      {stage3_5[53]},
      {stage4_5[40]}
   );
   gpc1_1 gpc4498 (
      {stage3_5[54]},
      {stage4_5[41]}
   );
   gpc1_1 gpc4499 (
      {stage3_5[55]},
      {stage4_5[42]}
   );
   gpc1_1 gpc4500 (
      {stage3_5[56]},
      {stage4_5[43]}
   );
   gpc1_1 gpc4501 (
      {stage3_5[57]},
      {stage4_5[44]}
   );
   gpc1_1 gpc4502 (
      {stage3_5[58]},
      {stage4_5[45]}
   );
   gpc1_1 gpc4503 (
      {stage3_6[30]},
      {stage4_6[15]}
   );
   gpc1_1 gpc4504 (
      {stage3_6[31]},
      {stage4_6[16]}
   );
   gpc1_1 gpc4505 (
      {stage3_6[32]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4506 (
      {stage3_6[33]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4507 (
      {stage3_6[34]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4508 (
      {stage3_6[35]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4509 (
      {stage3_6[36]},
      {stage4_6[21]}
   );
   gpc1_1 gpc4510 (
      {stage3_6[37]},
      {stage4_6[22]}
   );
   gpc1_1 gpc4511 (
      {stage3_7[45]},
      {stage4_7[13]}
   );
   gpc1_1 gpc4512 (
      {stage3_7[46]},
      {stage4_7[14]}
   );
   gpc1_1 gpc4513 (
      {stage3_8[85]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4514 (
      {stage3_8[86]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4515 (
      {stage3_8[87]},
      {stage4_8[23]}
   );
   gpc1_1 gpc4516 (
      {stage3_8[88]},
      {stage4_8[24]}
   );
   gpc1_1 gpc4517 (
      {stage3_8[89]},
      {stage4_8[25]}
   );
   gpc1_1 gpc4518 (
      {stage3_8[90]},
      {stage4_8[26]}
   );
   gpc1_1 gpc4519 (
      {stage3_8[91]},
      {stage4_8[27]}
   );
   gpc1_1 gpc4520 (
      {stage3_8[92]},
      {stage4_8[28]}
   );
   gpc1_1 gpc4521 (
      {stage3_9[30]},
      {stage4_9[22]}
   );
   gpc1_1 gpc4522 (
      {stage3_9[31]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4523 (
      {stage3_9[32]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4524 (
      {stage3_9[33]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4525 (
      {stage3_9[34]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4526 (
      {stage3_9[35]},
      {stage4_9[27]}
   );
   gpc1_1 gpc4527 (
      {stage3_9[36]},
      {stage4_9[28]}
   );
   gpc1_1 gpc4528 (
      {stage3_9[37]},
      {stage4_9[29]}
   );
   gpc1_1 gpc4529 (
      {stage3_9[38]},
      {stage4_9[30]}
   );
   gpc1_1 gpc4530 (
      {stage3_9[39]},
      {stage4_9[31]}
   );
   gpc1_1 gpc4531 (
      {stage3_9[40]},
      {stage4_9[32]}
   );
   gpc1_1 gpc4532 (
      {stage3_9[41]},
      {stage4_9[33]}
   );
   gpc1_1 gpc4533 (
      {stage3_9[42]},
      {stage4_9[34]}
   );
   gpc1_1 gpc4534 (
      {stage3_9[43]},
      {stage4_9[35]}
   );
   gpc1_1 gpc4535 (
      {stage3_9[44]},
      {stage4_9[36]}
   );
   gpc1_1 gpc4536 (
      {stage3_9[45]},
      {stage4_9[37]}
   );
   gpc1_1 gpc4537 (
      {stage3_9[46]},
      {stage4_9[38]}
   );
   gpc1_1 gpc4538 (
      {stage3_9[47]},
      {stage4_9[39]}
   );
   gpc1_1 gpc4539 (
      {stage3_9[48]},
      {stage4_9[40]}
   );
   gpc1_1 gpc4540 (
      {stage3_9[49]},
      {stage4_9[41]}
   );
   gpc1_1 gpc4541 (
      {stage3_11[31]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4542 (
      {stage3_11[32]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4543 (
      {stage3_11[33]},
      {stage4_11[21]}
   );
   gpc1_1 gpc4544 (
      {stage3_11[34]},
      {stage4_11[22]}
   );
   gpc1_1 gpc4545 (
      {stage3_11[35]},
      {stage4_11[23]}
   );
   gpc1_1 gpc4546 (
      {stage3_11[36]},
      {stage4_11[24]}
   );
   gpc1_1 gpc4547 (
      {stage3_11[37]},
      {stage4_11[25]}
   );
   gpc1_1 gpc4548 (
      {stage3_11[38]},
      {stage4_11[26]}
   );
   gpc1_1 gpc4549 (
      {stage3_11[39]},
      {stage4_11[27]}
   );
   gpc1_1 gpc4550 (
      {stage3_11[40]},
      {stage4_11[28]}
   );
   gpc1_1 gpc4551 (
      {stage3_11[41]},
      {stage4_11[29]}
   );
   gpc1_1 gpc4552 (
      {stage3_11[42]},
      {stage4_11[30]}
   );
   gpc1_1 gpc4553 (
      {stage3_11[43]},
      {stage4_11[31]}
   );
   gpc1_1 gpc4554 (
      {stage3_11[44]},
      {stage4_11[32]}
   );
   gpc1_1 gpc4555 (
      {stage3_11[45]},
      {stage4_11[33]}
   );
   gpc1_1 gpc4556 (
      {stage3_11[46]},
      {stage4_11[34]}
   );
   gpc1_1 gpc4557 (
      {stage3_11[47]},
      {stage4_11[35]}
   );
   gpc1_1 gpc4558 (
      {stage3_11[48]},
      {stage4_11[36]}
   );
   gpc1_1 gpc4559 (
      {stage3_11[49]},
      {stage4_11[37]}
   );
   gpc1_1 gpc4560 (
      {stage3_11[50]},
      {stage4_11[38]}
   );
   gpc1_1 gpc4561 (
      {stage3_11[51]},
      {stage4_11[39]}
   );
   gpc1_1 gpc4562 (
      {stage3_11[52]},
      {stage4_11[40]}
   );
   gpc1_1 gpc4563 (
      {stage3_11[53]},
      {stage4_11[41]}
   );
   gpc1_1 gpc4564 (
      {stage3_11[54]},
      {stage4_11[42]}
   );
   gpc1_1 gpc4565 (
      {stage3_12[38]},
      {stage4_12[15]}
   );
   gpc1_1 gpc4566 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc4567 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc4568 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc4569 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc4570 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc4571 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc4572 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc4573 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc4574 (
      {stage3_13[29]},
      {stage4_13[11]}
   );
   gpc1_1 gpc4575 (
      {stage3_13[30]},
      {stage4_13[12]}
   );
   gpc1_1 gpc4576 (
      {stage3_13[31]},
      {stage4_13[13]}
   );
   gpc1_1 gpc4577 (
      {stage3_13[32]},
      {stage4_13[14]}
   );
   gpc1_1 gpc4578 (
      {stage3_13[33]},
      {stage4_13[15]}
   );
   gpc1_1 gpc4579 (
      {stage3_13[34]},
      {stage4_13[16]}
   );
   gpc1_1 gpc4580 (
      {stage3_13[35]},
      {stage4_13[17]}
   );
   gpc1_1 gpc4581 (
      {stage3_13[36]},
      {stage4_13[18]}
   );
   gpc1_1 gpc4582 (
      {stage3_14[36]},
      {stage4_14[15]}
   );
   gpc1_1 gpc4583 (
      {stage3_14[37]},
      {stage4_14[16]}
   );
   gpc1_1 gpc4584 (
      {stage3_14[38]},
      {stage4_14[17]}
   );
   gpc1_1 gpc4585 (
      {stage3_14[39]},
      {stage4_14[18]}
   );
   gpc1_1 gpc4586 (
      {stage3_14[40]},
      {stage4_14[19]}
   );
   gpc1_1 gpc4587 (
      {stage3_14[41]},
      {stage4_14[20]}
   );
   gpc1_1 gpc4588 (
      {stage3_14[42]},
      {stage4_14[21]}
   );
   gpc1_1 gpc4589 (
      {stage3_14[43]},
      {stage4_14[22]}
   );
   gpc1_1 gpc4590 (
      {stage3_14[44]},
      {stage4_14[23]}
   );
   gpc1_1 gpc4591 (
      {stage3_14[45]},
      {stage4_14[24]}
   );
   gpc1_1 gpc4592 (
      {stage3_14[46]},
      {stage4_14[25]}
   );
   gpc1_1 gpc4593 (
      {stage3_14[47]},
      {stage4_14[26]}
   );
   gpc1_1 gpc4594 (
      {stage3_14[48]},
      {stage4_14[27]}
   );
   gpc1_1 gpc4595 (
      {stage3_14[49]},
      {stage4_14[28]}
   );
   gpc1_1 gpc4596 (
      {stage3_14[50]},
      {stage4_14[29]}
   );
   gpc1_1 gpc4597 (
      {stage3_14[51]},
      {stage4_14[30]}
   );
   gpc1_1 gpc4598 (
      {stage3_14[52]},
      {stage4_14[31]}
   );
   gpc1_1 gpc4599 (
      {stage3_14[53]},
      {stage4_14[32]}
   );
   gpc1_1 gpc4600 (
      {stage3_14[54]},
      {stage4_14[33]}
   );
   gpc1_1 gpc4601 (
      {stage3_14[55]},
      {stage4_14[34]}
   );
   gpc1_1 gpc4602 (
      {stage3_15[55]},
      {stage4_15[23]}
   );
   gpc1_1 gpc4603 (
      {stage3_15[56]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4604 (
      {stage3_15[57]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4605 (
      {stage3_15[58]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4606 (
      {stage3_15[59]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4607 (
      {stage3_15[60]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4608 (
      {stage3_15[61]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4609 (
      {stage3_15[62]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4610 (
      {stage3_15[63]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4611 (
      {stage3_15[64]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4612 (
      {stage3_15[65]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4613 (
      {stage3_15[66]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4614 (
      {stage3_15[67]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4615 (
      {stage3_15[68]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4616 (
      {stage3_15[69]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4617 (
      {stage3_15[70]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4618 (
      {stage3_17[55]},
      {stage4_17[21]}
   );
   gpc1_1 gpc4619 (
      {stage3_17[56]},
      {stage4_17[22]}
   );
   gpc1_1 gpc4620 (
      {stage3_17[57]},
      {stage4_17[23]}
   );
   gpc1_1 gpc4621 (
      {stage3_17[58]},
      {stage4_17[24]}
   );
   gpc1_1 gpc4622 (
      {stage3_17[59]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4623 (
      {stage3_17[60]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4624 (
      {stage3_17[61]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4625 (
      {stage3_17[62]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4626 (
      {stage3_17[63]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4627 (
      {stage3_17[64]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4628 (
      {stage3_17[65]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4629 (
      {stage3_17[66]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4630 (
      {stage3_17[67]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4631 (
      {stage3_17[68]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4632 (
      {stage3_17[69]},
      {stage4_17[35]}
   );
   gpc1_1 gpc4633 (
      {stage3_17[70]},
      {stage4_17[36]}
   );
   gpc1_1 gpc4634 (
      {stage3_17[71]},
      {stage4_17[37]}
   );
   gpc1_1 gpc4635 (
      {stage3_17[72]},
      {stage4_17[38]}
   );
   gpc1_1 gpc4636 (
      {stage3_17[73]},
      {stage4_17[39]}
   );
   gpc1_1 gpc4637 (
      {stage3_17[74]},
      {stage4_17[40]}
   );
   gpc1_1 gpc4638 (
      {stage3_17[75]},
      {stage4_17[41]}
   );
   gpc1_1 gpc4639 (
      {stage3_17[76]},
      {stage4_17[42]}
   );
   gpc1_1 gpc4640 (
      {stage3_18[25]},
      {stage4_18[19]}
   );
   gpc1_1 gpc4641 (
      {stage3_18[26]},
      {stage4_18[20]}
   );
   gpc1_1 gpc4642 (
      {stage3_18[27]},
      {stage4_18[21]}
   );
   gpc1_1 gpc4643 (
      {stage3_18[28]},
      {stage4_18[22]}
   );
   gpc1_1 gpc4644 (
      {stage3_18[29]},
      {stage4_18[23]}
   );
   gpc1_1 gpc4645 (
      {stage3_18[30]},
      {stage4_18[24]}
   );
   gpc1_1 gpc4646 (
      {stage3_18[31]},
      {stage4_18[25]}
   );
   gpc1_1 gpc4647 (
      {stage3_18[32]},
      {stage4_18[26]}
   );
   gpc1_1 gpc4648 (
      {stage3_18[33]},
      {stage4_18[27]}
   );
   gpc1_1 gpc4649 (
      {stage3_18[34]},
      {stage4_18[28]}
   );
   gpc1_1 gpc4650 (
      {stage3_19[62]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4651 (
      {stage3_19[63]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4652 (
      {stage3_19[64]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4653 (
      {stage3_19[65]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4654 (
      {stage3_19[66]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4655 (
      {stage3_19[67]},
      {stage4_19[29]}
   );
   gpc1_1 gpc4656 (
      {stage3_19[68]},
      {stage4_19[30]}
   );
   gpc1_1 gpc4657 (
      {stage3_19[69]},
      {stage4_19[31]}
   );
   gpc1_1 gpc4658 (
      {stage3_21[60]},
      {stage4_21[16]}
   );
   gpc1_1 gpc4659 (
      {stage3_21[61]},
      {stage4_21[17]}
   );
   gpc1_1 gpc4660 (
      {stage3_21[62]},
      {stage4_21[18]}
   );
   gpc1_1 gpc4661 (
      {stage3_22[37]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4662 (
      {stage3_22[38]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4663 (
      {stage3_22[39]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4664 (
      {stage3_22[40]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4665 (
      {stage3_22[41]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4666 (
      {stage3_22[42]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4667 (
      {stage3_22[43]},
      {stage4_22[23]}
   );
   gpc1_1 gpc4668 (
      {stage3_22[44]},
      {stage4_22[24]}
   );
   gpc1_1 gpc4669 (
      {stage3_22[45]},
      {stage4_22[25]}
   );
   gpc1_1 gpc4670 (
      {stage3_22[46]},
      {stage4_22[26]}
   );
   gpc1_1 gpc4671 (
      {stage3_22[47]},
      {stage4_22[27]}
   );
   gpc1_1 gpc4672 (
      {stage3_22[48]},
      {stage4_22[28]}
   );
   gpc1_1 gpc4673 (
      {stage3_22[49]},
      {stage4_22[29]}
   );
   gpc1_1 gpc4674 (
      {stage3_22[50]},
      {stage4_22[30]}
   );
   gpc1_1 gpc4675 (
      {stage3_23[29]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4676 (
      {stage3_23[30]},
      {stage4_23[22]}
   );
   gpc1_1 gpc4677 (
      {stage3_23[31]},
      {stage4_23[23]}
   );
   gpc1_1 gpc4678 (
      {stage3_23[32]},
      {stage4_23[24]}
   );
   gpc1_1 gpc4679 (
      {stage3_23[33]},
      {stage4_23[25]}
   );
   gpc1_1 gpc4680 (
      {stage3_23[34]},
      {stage4_23[26]}
   );
   gpc1_1 gpc4681 (
      {stage3_23[35]},
      {stage4_23[27]}
   );
   gpc1_1 gpc4682 (
      {stage3_23[36]},
      {stage4_23[28]}
   );
   gpc1_1 gpc4683 (
      {stage3_23[37]},
      {stage4_23[29]}
   );
   gpc1_1 gpc4684 (
      {stage3_23[38]},
      {stage4_23[30]}
   );
   gpc1_1 gpc4685 (
      {stage3_23[39]},
      {stage4_23[31]}
   );
   gpc1_1 gpc4686 (
      {stage3_23[40]},
      {stage4_23[32]}
   );
   gpc1_1 gpc4687 (
      {stage3_23[41]},
      {stage4_23[33]}
   );
   gpc1_1 gpc4688 (
      {stage3_23[42]},
      {stage4_23[34]}
   );
   gpc1_1 gpc4689 (
      {stage3_23[43]},
      {stage4_23[35]}
   );
   gpc1_1 gpc4690 (
      {stage3_23[44]},
      {stage4_23[36]}
   );
   gpc1_1 gpc4691 (
      {stage3_23[45]},
      {stage4_23[37]}
   );
   gpc1_1 gpc4692 (
      {stage3_24[47]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4693 (
      {stage3_24[48]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4694 (
      {stage3_24[49]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4695 (
      {stage3_24[50]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4696 (
      {stage3_24[51]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4697 (
      {stage3_24[52]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4698 (
      {stage3_24[53]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4699 (
      {stage3_24[54]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4700 (
      {stage3_24[55]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4701 (
      {stage3_24[56]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4702 (
      {stage3_24[57]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4703 (
      {stage3_24[58]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4704 (
      {stage3_24[59]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4705 (
      {stage3_24[60]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4706 (
      {stage3_25[47]},
      {stage4_25[17]}
   );
   gpc1_1 gpc4707 (
      {stage3_25[48]},
      {stage4_25[18]}
   );
   gpc1_1 gpc4708 (
      {stage3_26[46]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4709 (
      {stage3_26[47]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4710 (
      {stage3_26[48]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4711 (
      {stage3_26[49]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4712 (
      {stage3_26[50]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4713 (
      {stage3_27[48]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4714 (
      {stage3_27[49]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4715 (
      {stage3_27[50]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4716 (
      {stage3_27[51]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4717 (
      {stage3_27[52]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4718 (
      {stage3_27[53]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4719 (
      {stage3_27[54]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4720 (
      {stage3_30[68]},
      {stage4_30[24]}
   );
   gpc1_1 gpc4721 (
      {stage3_30[69]},
      {stage4_30[25]}
   );
   gpc1_1 gpc4722 (
      {stage3_30[70]},
      {stage4_30[26]}
   );
   gpc1_1 gpc4723 (
      {stage3_31[51]},
      {stage4_31[24]}
   );
   gpc1_1 gpc4724 (
      {stage3_31[52]},
      {stage4_31[25]}
   );
   gpc1_1 gpc4725 (
      {stage3_31[53]},
      {stage4_31[26]}
   );
   gpc1_1 gpc4726 (
      {stage3_31[54]},
      {stage4_31[27]}
   );
   gpc1_1 gpc4727 (
      {stage3_31[55]},
      {stage4_31[28]}
   );
   gpc1_1 gpc4728 (
      {stage3_31[56]},
      {stage4_31[29]}
   );
   gpc1_1 gpc4729 (
      {stage3_31[57]},
      {stage4_31[30]}
   );
   gpc1_1 gpc4730 (
      {stage3_32[39]},
      {stage4_32[24]}
   );
   gpc1_1 gpc4731 (
      {stage3_32[40]},
      {stage4_32[25]}
   );
   gpc1_1 gpc4732 (
      {stage3_32[41]},
      {stage4_32[26]}
   );
   gpc1_1 gpc4733 (
      {stage3_32[42]},
      {stage4_32[27]}
   );
   gpc1_1 gpc4734 (
      {stage3_32[43]},
      {stage4_32[28]}
   );
   gpc1_1 gpc4735 (
      {stage3_32[44]},
      {stage4_32[29]}
   );
   gpc1_1 gpc4736 (
      {stage3_32[45]},
      {stage4_32[30]}
   );
   gpc1_1 gpc4737 (
      {stage3_32[46]},
      {stage4_32[31]}
   );
   gpc1_1 gpc4738 (
      {stage3_32[47]},
      {stage4_32[32]}
   );
   gpc1_1 gpc4739 (
      {stage3_32[48]},
      {stage4_32[33]}
   );
   gpc1_1 gpc4740 (
      {stage3_32[49]},
      {stage4_32[34]}
   );
   gpc1_1 gpc4741 (
      {stage3_32[50]},
      {stage4_32[35]}
   );
   gpc1_1 gpc4742 (
      {stage3_32[51]},
      {stage4_32[36]}
   );
   gpc1_1 gpc4743 (
      {stage3_32[52]},
      {stage4_32[37]}
   );
   gpc1_1 gpc4744 (
      {stage3_32[53]},
      {stage4_32[38]}
   );
   gpc1_1 gpc4745 (
      {stage3_32[54]},
      {stage4_32[39]}
   );
   gpc1_1 gpc4746 (
      {stage3_32[55]},
      {stage4_32[40]}
   );
   gpc1_1 gpc4747 (
      {stage3_32[56]},
      {stage4_32[41]}
   );
   gpc1_1 gpc4748 (
      {stage3_32[57]},
      {stage4_32[42]}
   );
   gpc1_1 gpc4749 (
      {stage3_33[24]},
      {stage4_33[16]}
   );
   gpc1_1 gpc4750 (
      {stage3_33[25]},
      {stage4_33[17]}
   );
   gpc1_1 gpc4751 (
      {stage3_33[26]},
      {stage4_33[18]}
   );
   gpc1_1 gpc4752 (
      {stage3_34[24]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4753 (
      {stage3_34[25]},
      {stage4_34[11]}
   );
   gpc1_1 gpc4754 (
      {stage3_34[26]},
      {stage4_34[12]}
   );
   gpc1_1 gpc4755 (
      {stage3_35[6]},
      {stage4_35[8]}
   );
   gpc1_1 gpc4756 (
      {stage3_35[7]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4757 (
      {stage3_35[8]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4758 (
      {stage3_35[9]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4759 (
      {stage3_35[10]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4760 (
      {stage3_35[11]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4761 (
      {stage3_35[12]},
      {stage4_35[14]}
   );
   gpc1_1 gpc4762 (
      {stage3_36[0]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4763 (
      {stage3_36[1]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4764 (
      {stage3_36[2]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4765 (
      {stage3_36[3]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4766 (
      {stage3_36[4]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4767 (
      {stage3_36[5]},
      {stage4_36[10]}
   );
   gpc1_1 gpc4768 (
      {stage3_37[0]},
      {stage4_37[1]}
   );
   gpc1_1 gpc4769 (
      {stage3_37[1]},
      {stage4_37[2]}
   );
   gpc606_5 gpc4770 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc615_5 gpc4771 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[6]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc615_5 gpc4772 (
      {stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2]}
   );
   gpc615_5 gpc4773 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16]},
      {stage4_4[7]},
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc615_5 gpc4774 (
      {stage4_3[17], stage4_3[18], stage4_3[19], stage4_3[20], stage4_3[21]},
      {stage4_4[8]},
      {stage4_5[12], stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17]},
      {stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[4],stage5_3[4]}
   );
   gpc606_5 gpc4775 (
      {stage4_4[9], stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc4776 (
      {stage4_4[15], stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc7_3 gpc4777 (
      {stage4_5[18], stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc7_3 gpc4778 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc7_3 gpc4779 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37], stage4_5[38]},
      {stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc7_3 gpc4780 (
      {stage4_5[39], stage4_5[40], stage4_5[41], stage4_5[42], stage4_5[43], stage4_5[44], stage4_5[45]},
      {stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc615_5 gpc4781 (
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[2],stage5_7[9],stage5_6[10]}
   );
   gpc615_5 gpc4782 (
      {stage4_6[17], stage4_6[18], stage4_6[19], stage4_6[20], stage4_6[21]},
      {stage4_7[1]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[3],stage5_7[10],stage5_6[11]}
   );
   gpc1163_5 gpc4783 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[0]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[4],stage5_7[11]}
   );
   gpc623_5 gpc4784 (
      {stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[18], stage4_8[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[5],stage5_7[12]}
   );
   gpc606_5 gpc4785 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc4786 (
      {stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc4787 (
      {stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[6]}
   );
   gpc606_5 gpc4788 (
      {stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[3],stage5_11[5],stage5_10[7],stage5_9[7]}
   );
   gpc606_5 gpc4789 (
      {stage4_9[25], stage4_9[26], stage4_9[27], stage4_9[28], stage4_9[29], stage4_9[30]},
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage5_13[3],stage5_12[4],stage5_11[6],stage5_10[8],stage5_9[8]}
   );
   gpc606_5 gpc4790 (
      {stage4_9[31], stage4_9[32], stage4_9[33], stage4_9[34], stage4_9[35], stage4_9[36]},
      {stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27], stage4_11[28], stage4_11[29]},
      {stage5_13[4],stage5_12[5],stage5_11[7],stage5_10[9],stage5_9[9]}
   );
   gpc615_5 gpc4791 (
      {stage4_9[37], stage4_9[38], stage4_9[39], stage4_9[40], stage4_9[41]},
      {stage4_10[7]},
      {stage4_11[30], stage4_11[31], stage4_11[32], stage4_11[33], stage4_11[34], stage4_11[35]},
      {stage5_13[5],stage5_12[6],stage5_11[8],stage5_10[10],stage5_9[10]}
   );
   gpc615_5 gpc4792 (
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12]},
      {stage4_11[36]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[6],stage5_12[7],stage5_11[9],stage5_10[11]}
   );
   gpc615_5 gpc4793 (
      {stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_11[37]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[7],stage5_12[8],stage5_11[10],stage5_10[12]}
   );
   gpc606_5 gpc4794 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[8],stage5_12[9]}
   );
   gpc606_5 gpc4795 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[9],stage5_12[10]}
   );
   gpc1163_5 gpc4796 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[10]}
   );
   gpc1163_5 gpc4797 (
      {stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_14[18], stage4_14[19], stage4_14[20], stage4_14[21], stage4_14[22], stage4_14[23]},
      {stage4_15[1]},
      {stage4_16[1]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[11]}
   );
   gpc1163_5 gpc4798 (
      {stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_14[24], stage4_14[25], stage4_14[26], stage4_14[27], stage4_14[28], stage4_14[29]},
      {stage4_15[2]},
      {stage4_16[2]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[12]}
   );
   gpc606_5 gpc4799 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage5_17[3],stage5_16[5],stage5_15[5],stage5_14[7],stage5_13[13]}
   );
   gpc606_5 gpc4800 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], 1'b0, 1'b0},
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13], stage4_15[14]},
      {stage5_17[4],stage5_16[6],stage5_15[6],stage5_14[8],stage5_13[14]}
   );
   gpc135_4 gpc4801 (
      {stage4_14[30], stage4_14[31], stage4_14[32], stage4_14[33], stage4_14[34]},
      {stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage4_16[3]},
      {stage5_17[5],stage5_16[7],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc4802 (
      {stage4_15[18], stage4_15[19], stage4_15[20], stage4_15[21], stage4_15[22]},
      {stage4_16[4]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[6],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4803 (
      {stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26], stage4_15[27]},
      {stage4_16[5]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[1],stage5_17[7],stage5_16[9],stage5_15[9]}
   );
   gpc615_5 gpc4804 (
      {stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31], stage4_15[32]},
      {stage4_16[6]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[2],stage5_17[8],stage5_16[10],stage5_15[10]}
   );
   gpc615_5 gpc4805 (
      {stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36], stage4_15[37]},
      {stage4_16[7]},
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23]},
      {stage5_19[3],stage5_18[3],stage5_17[9],stage5_16[11],stage5_15[11]}
   );
   gpc606_5 gpc4806 (
      {stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12], stage4_16[13]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[4],stage5_18[4],stage5_17[10],stage5_16[12]}
   );
   gpc615_5 gpc4807 (
      {stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_17[24]},
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage5_20[1],stage5_19[5],stage5_18[5],stage5_17[11],stage5_16[13]}
   );
   gpc606_5 gpc4808 (
      {stage4_17[25], stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[6],stage5_18[6],stage5_17[12]}
   );
   gpc606_5 gpc4809 (
      {stage4_17[31], stage4_17[32], stage4_17[33], stage4_17[34], stage4_17[35], stage4_17[36]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[3],stage5_19[7],stage5_18[7],stage5_17[13]}
   );
   gpc606_5 gpc4810 (
      {stage4_17[37], stage4_17[38], stage4_17[39], stage4_17[40], stage4_17[41], stage4_17[42]},
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17]},
      {stage5_21[2],stage5_20[4],stage5_19[8],stage5_18[8],stage5_17[14]}
   );
   gpc606_5 gpc4811 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[3],stage5_20[5],stage5_19[9],stage5_18[9]}
   );
   gpc615_5 gpc4812 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[18]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[4],stage5_20[6],stage5_19[10],stage5_18[10]}
   );
   gpc615_5 gpc4813 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[0]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[2],stage5_21[5]}
   );
   gpc615_5 gpc4814 (
      {stage4_21[5], stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9]},
      {stage4_22[1]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[1],stage5_22[3],stage5_21[6]}
   );
   gpc615_5 gpc4815 (
      {stage4_21[10], stage4_21[11], stage4_21[12], stage4_21[13], stage4_21[14]},
      {stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage5_25[2],stage5_24[2],stage5_23[2],stage5_22[4],stage5_21[7]}
   );
   gpc615_5 gpc4816 (
      {stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18], 1'b0},
      {stage4_22[3]},
      {stage4_23[18], stage4_23[19], stage4_23[20], stage4_23[21], stage4_23[22], stage4_23[23]},
      {stage5_25[3],stage5_24[3],stage5_23[3],stage5_22[5],stage5_21[8]}
   );
   gpc615_5 gpc4817 (
      {stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[24]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[4],stage5_24[4],stage5_23[4],stage5_22[6]}
   );
   gpc615_5 gpc4818 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[25]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[5],stage5_24[5],stage5_23[5],stage5_22[7]}
   );
   gpc615_5 gpc4819 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[26]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[6],stage5_24[6],stage5_23[6],stage5_22[8]}
   );
   gpc615_5 gpc4820 (
      {stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22], stage4_22[23]},
      {stage4_23[27]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[7],stage5_24[7],stage5_23[7],stage5_22[9]}
   );
   gpc615_5 gpc4821 (
      {stage4_23[28], stage4_23[29], stage4_23[30], stage4_23[31], stage4_23[32]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[8],stage5_24[8],stage5_23[8]}
   );
   gpc615_5 gpc4822 (
      {stage4_23[33], stage4_23[34], stage4_23[35], stage4_23[36], stage4_23[37]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[9],stage5_24[9],stage5_23[9]}
   );
   gpc606_5 gpc4823 (
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[6],stage5_25[10]}
   );
   gpc615_5 gpc4824 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4]},
      {stage4_27[6]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[7]}
   );
   gpc615_5 gpc4825 (
      {stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9]},
      {stage4_27[7]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4826 (
      {stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14]},
      {stage4_27[8]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[3],stage5_28[3],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4827 (
      {stage4_26[15], stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19]},
      {stage4_27[9]},
      {stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22], stage4_28[23]},
      {stage5_30[3],stage5_29[4],stage5_28[4],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4828 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[4],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc615_5 gpc4829 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21]},
      {stage4_28[24]},
      {stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7]},
      {stage5_31[0],stage5_30[5],stage5_29[6],stage5_28[6],stage5_27[8]}
   );
   gpc615_5 gpc4830 (
      {stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[6],stage5_29[7]}
   );
   gpc615_5 gpc4831 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[2],stage5_30[7],stage5_29[8]}
   );
   gpc615_5 gpc4832 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22]},
      {stage4_30[2]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], stage4_31[17]},
      {stage5_33[2],stage5_32[2],stage5_31[3],stage5_30[8],stage5_29[9]}
   );
   gpc615_5 gpc4833 (
      {stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7]},
      {stage4_31[18]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[3],stage5_32[3],stage5_31[4],stage5_30[9]}
   );
   gpc615_5 gpc4834 (
      {stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12]},
      {stage4_31[19]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[4],stage5_32[4],stage5_31[5],stage5_30[10]}
   );
   gpc615_5 gpc4835 (
      {stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage4_31[20]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[5],stage5_32[5],stage5_31[6],stage5_30[11]}
   );
   gpc615_5 gpc4836 (
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22]},
      {stage4_31[21]},
      {stage4_32[18], stage4_32[19], stage4_32[20], stage4_32[21], stage4_32[22], stage4_32[23]},
      {stage5_34[3],stage5_33[6],stage5_32[6],stage5_31[7],stage5_30[12]}
   );
   gpc615_5 gpc4837 (
      {stage4_31[22], stage4_31[23], stage4_31[24], stage4_31[25], stage4_31[26]},
      {stage4_32[24]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[4],stage5_33[7],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc4838 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[5],stage5_33[8]}
   );
   gpc606_5 gpc4839 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[6],stage5_33[9]}
   );
   gpc606_5 gpc4840 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3],stage5_34[7]}
   );
   gpc606_5 gpc4841 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], 1'b0},
      {stage5_38[1],stage5_37[3],stage5_36[3],stage5_35[4],stage5_34[8]}
   );
   gpc1_1 gpc4842 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4843 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4844 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4845 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc4846 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc4847 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc4848 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc4849 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc4850 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc4851 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc4852 (
      {stage4_0[10]},
      {stage5_0[10]}
   );
   gpc1_1 gpc4853 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4854 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4855 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4856 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4857 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4858 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4859 (
      {stage4_1[12]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4860 (
      {stage4_1[13]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4861 (
      {stage4_1[14]},
      {stage5_1[9]}
   );
   gpc1_1 gpc4862 (
      {stage4_1[15]},
      {stage5_1[10]}
   );
   gpc1_1 gpc4863 (
      {stage4_2[5]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4864 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4865 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4866 (
      {stage4_2[8]},
      {stage5_2[5]}
   );
   gpc1_1 gpc4867 (
      {stage4_2[9]},
      {stage5_2[6]}
   );
   gpc1_1 gpc4868 (
      {stage4_2[10]},
      {stage5_2[7]}
   );
   gpc1_1 gpc4869 (
      {stage4_2[11]},
      {stage5_2[8]}
   );
   gpc1_1 gpc4870 (
      {stage4_2[12]},
      {stage5_2[9]}
   );
   gpc1_1 gpc4871 (
      {stage4_3[22]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4872 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc4873 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc4874 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc4875 (
      {stage4_6[22]},
      {stage5_6[12]}
   );
   gpc1_1 gpc4876 (
      {stage4_7[8]},
      {stage5_7[13]}
   );
   gpc1_1 gpc4877 (
      {stage4_7[9]},
      {stage5_7[14]}
   );
   gpc1_1 gpc4878 (
      {stage4_7[10]},
      {stage5_7[15]}
   );
   gpc1_1 gpc4879 (
      {stage4_7[11]},
      {stage5_7[16]}
   );
   gpc1_1 gpc4880 (
      {stage4_7[12]},
      {stage5_7[17]}
   );
   gpc1_1 gpc4881 (
      {stage4_7[13]},
      {stage5_7[18]}
   );
   gpc1_1 gpc4882 (
      {stage4_7[14]},
      {stage5_7[19]}
   );
   gpc1_1 gpc4883 (
      {stage4_8[26]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4884 (
      {stage4_8[27]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4885 (
      {stage4_8[28]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4886 (
      {stage4_11[38]},
      {stage5_11[11]}
   );
   gpc1_1 gpc4887 (
      {stage4_11[39]},
      {stage5_11[12]}
   );
   gpc1_1 gpc4888 (
      {stage4_11[40]},
      {stage5_11[13]}
   );
   gpc1_1 gpc4889 (
      {stage4_11[41]},
      {stage5_11[14]}
   );
   gpc1_1 gpc4890 (
      {stage4_11[42]},
      {stage5_11[15]}
   );
   gpc1_1 gpc4891 (
      {stage4_15[38]},
      {stage5_15[12]}
   );
   gpc1_1 gpc4892 (
      {stage4_16[19]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4893 (
      {stage4_18[23]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4894 (
      {stage4_18[24]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4895 (
      {stage4_18[25]},
      {stage5_18[13]}
   );
   gpc1_1 gpc4896 (
      {stage4_18[26]},
      {stage5_18[14]}
   );
   gpc1_1 gpc4897 (
      {stage4_18[27]},
      {stage5_18[15]}
   );
   gpc1_1 gpc4898 (
      {stage4_18[28]},
      {stage5_18[16]}
   );
   gpc1_1 gpc4899 (
      {stage4_19[19]},
      {stage5_19[11]}
   );
   gpc1_1 gpc4900 (
      {stage4_19[20]},
      {stage5_19[12]}
   );
   gpc1_1 gpc4901 (
      {stage4_19[21]},
      {stage5_19[13]}
   );
   gpc1_1 gpc4902 (
      {stage4_19[22]},
      {stage5_19[14]}
   );
   gpc1_1 gpc4903 (
      {stage4_19[23]},
      {stage5_19[15]}
   );
   gpc1_1 gpc4904 (
      {stage4_19[24]},
      {stage5_19[16]}
   );
   gpc1_1 gpc4905 (
      {stage4_19[25]},
      {stage5_19[17]}
   );
   gpc1_1 gpc4906 (
      {stage4_19[26]},
      {stage5_19[18]}
   );
   gpc1_1 gpc4907 (
      {stage4_19[27]},
      {stage5_19[19]}
   );
   gpc1_1 gpc4908 (
      {stage4_19[28]},
      {stage5_19[20]}
   );
   gpc1_1 gpc4909 (
      {stage4_19[29]},
      {stage5_19[21]}
   );
   gpc1_1 gpc4910 (
      {stage4_19[30]},
      {stage5_19[22]}
   );
   gpc1_1 gpc4911 (
      {stage4_19[31]},
      {stage5_19[23]}
   );
   gpc1_1 gpc4912 (
      {stage4_20[12]},
      {stage5_20[7]}
   );
   gpc1_1 gpc4913 (
      {stage4_20[13]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4914 (
      {stage4_20[14]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4915 (
      {stage4_20[15]},
      {stage5_20[10]}
   );
   gpc1_1 gpc4916 (
      {stage4_20[16]},
      {stage5_20[11]}
   );
   gpc1_1 gpc4917 (
      {stage4_20[17]},
      {stage5_20[12]}
   );
   gpc1_1 gpc4918 (
      {stage4_20[18]},
      {stage5_20[13]}
   );
   gpc1_1 gpc4919 (
      {stage4_22[24]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4920 (
      {stage4_22[25]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4921 (
      {stage4_22[26]},
      {stage5_22[12]}
   );
   gpc1_1 gpc4922 (
      {stage4_22[27]},
      {stage5_22[13]}
   );
   gpc1_1 gpc4923 (
      {stage4_22[28]},
      {stage5_22[14]}
   );
   gpc1_1 gpc4924 (
      {stage4_22[29]},
      {stage5_22[15]}
   );
   gpc1_1 gpc4925 (
      {stage4_22[30]},
      {stage5_22[16]}
   );
   gpc1_1 gpc4926 (
      {stage4_24[26]},
      {stage5_24[10]}
   );
   gpc1_1 gpc4927 (
      {stage4_24[27]},
      {stage5_24[11]}
   );
   gpc1_1 gpc4928 (
      {stage4_24[28]},
      {stage5_24[12]}
   );
   gpc1_1 gpc4929 (
      {stage4_24[29]},
      {stage5_24[13]}
   );
   gpc1_1 gpc4930 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc4931 (
      {stage4_26[20]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4932 (
      {stage4_26[21]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4933 (
      {stage4_26[22]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4934 (
      {stage4_27[22]},
      {stage5_27[9]}
   );
   gpc1_1 gpc4935 (
      {stage4_27[23]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4936 (
      {stage4_27[24]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4937 (
      {stage4_27[25]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4938 (
      {stage4_27[26]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4939 (
      {stage4_29[23]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4940 (
      {stage4_29[24]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4941 (
      {stage4_29[25]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4942 (
      {stage4_30[23]},
      {stage5_30[13]}
   );
   gpc1_1 gpc4943 (
      {stage4_30[24]},
      {stage5_30[14]}
   );
   gpc1_1 gpc4944 (
      {stage4_30[25]},
      {stage5_30[15]}
   );
   gpc1_1 gpc4945 (
      {stage4_30[26]},
      {stage5_30[16]}
   );
   gpc1_1 gpc4946 (
      {stage4_31[27]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4947 (
      {stage4_31[28]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4948 (
      {stage4_31[29]},
      {stage5_31[11]}
   );
   gpc1_1 gpc4949 (
      {stage4_31[30]},
      {stage5_31[12]}
   );
   gpc1_1 gpc4950 (
      {stage4_32[25]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4951 (
      {stage4_32[26]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4952 (
      {stage4_32[27]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4953 (
      {stage4_32[28]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4954 (
      {stage4_32[29]},
      {stage5_32[12]}
   );
   gpc1_1 gpc4955 (
      {stage4_32[30]},
      {stage5_32[13]}
   );
   gpc1_1 gpc4956 (
      {stage4_32[31]},
      {stage5_32[14]}
   );
   gpc1_1 gpc4957 (
      {stage4_32[32]},
      {stage5_32[15]}
   );
   gpc1_1 gpc4958 (
      {stage4_32[33]},
      {stage5_32[16]}
   );
   gpc1_1 gpc4959 (
      {stage4_32[34]},
      {stage5_32[17]}
   );
   gpc1_1 gpc4960 (
      {stage4_32[35]},
      {stage5_32[18]}
   );
   gpc1_1 gpc4961 (
      {stage4_32[36]},
      {stage5_32[19]}
   );
   gpc1_1 gpc4962 (
      {stage4_32[37]},
      {stage5_32[20]}
   );
   gpc1_1 gpc4963 (
      {stage4_32[38]},
      {stage5_32[21]}
   );
   gpc1_1 gpc4964 (
      {stage4_32[39]},
      {stage5_32[22]}
   );
   gpc1_1 gpc4965 (
      {stage4_32[40]},
      {stage5_32[23]}
   );
   gpc1_1 gpc4966 (
      {stage4_32[41]},
      {stage5_32[24]}
   );
   gpc1_1 gpc4967 (
      {stage4_32[42]},
      {stage5_32[25]}
   );
   gpc1_1 gpc4968 (
      {stage4_33[18]},
      {stage5_33[10]}
   );
   gpc1_1 gpc4969 (
      {stage4_34[12]},
      {stage5_34[9]}
   );
   gpc1_1 gpc4970 (
      {stage4_35[12]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4971 (
      {stage4_35[13]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4972 (
      {stage4_35[14]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4973 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4974 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4975 (
      {stage4_37[2]},
      {stage5_37[6]}
   );
   gpc1343_5 gpc4976 (
      {stage5_0[0], stage5_0[1], stage5_0[2]},
      {stage5_1[0], stage5_1[1], stage5_1[2], stage5_1[3]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc1343_5 gpc4977 (
      {stage5_0[3], stage5_0[4], stage5_0[5]},
      {stage5_1[4], stage5_1[5], stage5_1[6], stage5_1[7]},
      {stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[1]},
      {stage6_4[1],stage6_3[1],stage6_2[1],stage6_1[1],stage6_0[1]}
   );
   gpc117_4 gpc4978 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_5[0]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[2]}
   );
   gpc1343_5 gpc4979 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc4980 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc1343_5 gpc4981 (
      {stage5_5[7], stage5_5[8], stage5_5[9]},
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12]},
      {stage5_7[6], stage5_7[7], stage5_7[8]},
      {stage5_8[2]},
      {stage6_9[2],stage6_8[2],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc606_5 gpc4982 (
      {stage5_7[9], stage5_7[10], stage5_7[11], stage5_7[12], stage5_7[13], stage5_7[14]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[4]}
   );
   gpc615_5 gpc4983 (
      {stage5_7[15], stage5_7[16], stage5_7[17], stage5_7[18], stage5_7[19]},
      {stage5_8[3]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], 1'b0},
      {stage6_11[1],stage6_10[1],stage6_9[4],stage6_8[4],stage6_7[5]}
   );
   gpc606_5 gpc4984 (
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[2],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc7_3 gpc4985 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12]},
      {stage6_12[1],stage6_11[3],stage6_10[3]}
   );
   gpc207_4 gpc4986 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1]},
      {stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[4]}
   );
   gpc207_4 gpc4987 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[2], stage5_13[3]},
      {stage6_14[1],stage6_13[1],stage6_12[3],stage6_11[5]}
   );
   gpc7_3 gpc4988 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[2],stage6_13[2],stage6_12[4]}
   );
   gpc623_5 gpc4989 (
      {stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[5]}
   );
   gpc623_5 gpc4990 (
      {stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6], stage5_14[7]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc623_5 gpc4991 (
      {stage5_13[9], stage5_13[10], stage5_13[11]},
      {stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5],stage6_13[5]}
   );
   gpc207_4 gpc4992 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6]},
      {stage5_18[0], stage5_18[1]},
      {stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[3]}
   );
   gpc207_4 gpc4993 (
      {stage5_16[7], stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13]},
      {stage5_18[2], stage5_18[3]},
      {stage6_19[1],stage6_18[1],stage6_17[3],stage6_16[4]}
   );
   gpc1163_5 gpc4994 (
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[4], stage5_18[5], stage5_18[6], stage5_18[7], stage5_18[8], stage5_18[9]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[2],stage6_18[2],stage6_17[4]}
   );
   gpc1163_5 gpc4995 (
      {stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13], stage5_18[14], stage5_18[15]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[3],stage6_18[3],stage6_17[5]}
   );
   gpc606_5 gpc4996 (
      {stage5_17[6], stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[4],stage6_18[4],stage6_17[6]}
   );
   gpc207_4 gpc4997 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13], stage5_19[14]},
      {stage5_21[0], stage5_21[1]},
      {stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[5]}
   );
   gpc606_5 gpc4998 (
      {stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc606_5 gpc4999 (
      {stage5_20[8], stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13]},
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10], stage5_22[11]},
      {stage6_24[1],stage6_23[1],stage6_22[2],stage6_21[5],stage6_20[5]}
   );
   gpc1415_5 gpc5000 (
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[2]}
   );
   gpc615_5 gpc5001 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[1]},
      {stage5_25[4], stage5_25[5], stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9]},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3],stage6_23[3]}
   );
   gpc606_5 gpc5002 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5], stage5_26[6]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[4]}
   );
   gpc606_5 gpc5003 (
      {stage5_24[8], stage5_24[9], stage5_24[10], stage5_24[11], stage5_24[12], stage5_24[13]},
      {stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10], stage5_26[11], stage5_26[12]},
      {stage6_28[1],stage6_27[3],stage6_26[3],stage6_25[3],stage6_24[5]}
   );
   gpc606_5 gpc5004 (
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc5005 (
      {stage5_27[6], stage5_27[7], stage5_27[8], stage5_27[9], stage5_27[10], stage5_27[11]},
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage6_31[1],stage6_30[1],stage6_29[1],stage6_28[3],stage6_27[5]}
   );
   gpc207_4 gpc5006 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], stage5_28[6]},
      {stage5_30[0], stage5_30[1]},
      {stage6_31[2],stage6_30[2],stage6_29[2],stage6_28[4]}
   );
   gpc615_5 gpc5007 (
      {stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[0],stage6_32[0],stage6_31[3],stage6_30[3]}
   );
   gpc615_5 gpc5008 (
      {stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10], stage5_30[11]},
      {stage5_31[1]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[1],stage6_32[1],stage6_31[4],stage6_30[4]}
   );
   gpc615_5 gpc5009 (
      {stage5_30[12], stage5_30[13], stage5_30[14], stage5_30[15], stage5_30[16]},
      {stage5_31[2]},
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage6_34[2],stage6_33[2],stage6_32[2],stage6_31[5],stage6_30[5]}
   );
   gpc615_5 gpc5010 (
      {stage5_31[3], stage5_31[4], stage5_31[5], stage5_31[6], stage5_31[7]},
      {stage5_32[18]},
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage6_35[0],stage6_34[3],stage6_33[3],stage6_32[3],stage6_31[6]}
   );
   gpc615_5 gpc5011 (
      {stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11], stage5_31[12]},
      {stage5_32[19]},
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], 1'b0},
      {stage6_35[1],stage6_34[4],stage6_33[4],stage6_32[4],stage6_31[7]}
   );
   gpc606_5 gpc5012 (
      {stage5_32[20], stage5_32[21], stage5_32[22], stage5_32[23], stage5_32[24], stage5_32[25]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[2],stage6_34[5],stage6_33[5],stage6_32[5]}
   );
   gpc606_5 gpc5013 (
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[0],stage6_36[1],stage6_35[3]}
   );
   gpc1325_5 gpc5014 (
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], 1'b0},
      {stage5_37[6], 1'b0},
      {stage5_38[0], stage5_38[1], 1'b0},
      {1'b0},
      {stage6_40[0],stage6_39[1],stage6_38[1],stage6_37[1],stage6_36[2]}
   );
   gpc1_1 gpc5015 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc5016 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc5017 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc5018 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc5019 (
      {stage5_0[10]},
      {stage6_0[6]}
   );
   gpc1_1 gpc5020 (
      {stage5_1[8]},
      {stage6_1[2]}
   );
   gpc1_1 gpc5021 (
      {stage5_1[9]},
      {stage6_1[3]}
   );
   gpc1_1 gpc5022 (
      {stage5_1[10]},
      {stage6_1[4]}
   );
   gpc1_1 gpc5023 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc5024 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc5025 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc5026 (
      {stage5_2[9]},
      {stage6_2[5]}
   );
   gpc1_1 gpc5027 (
      {stage5_3[2]},
      {stage6_3[2]}
   );
   gpc1_1 gpc5028 (
      {stage5_3[3]},
      {stage6_3[3]}
   );
   gpc1_1 gpc5029 (
      {stage5_3[4]},
      {stage6_3[4]}
   );
   gpc1_1 gpc5030 (
      {stage5_3[5]},
      {stage6_3[5]}
   );
   gpc1_1 gpc5031 (
      {stage5_4[7]},
      {stage6_4[3]}
   );
   gpc1_1 gpc5032 (
      {stage5_4[8]},
      {stage6_4[4]}
   );
   gpc1_1 gpc5033 (
      {stage5_4[9]},
      {stage6_4[5]}
   );
   gpc1_1 gpc5034 (
      {stage5_5[10]},
      {stage6_5[4]}
   );
   gpc1_1 gpc5035 (
      {stage5_11[14]},
      {stage6_11[6]}
   );
   gpc1_1 gpc5036 (
      {stage5_11[15]},
      {stage6_11[7]}
   );
   gpc1_1 gpc5037 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc5038 (
      {stage5_13[12]},
      {stage6_13[6]}
   );
   gpc1_1 gpc5039 (
      {stage5_13[13]},
      {stage6_13[7]}
   );
   gpc1_1 gpc5040 (
      {stage5_13[14]},
      {stage6_13[8]}
   );
   gpc1_1 gpc5041 (
      {stage5_15[12]},
      {stage6_15[3]}
   );
   gpc1_1 gpc5042 (
      {stage5_16[14]},
      {stage6_16[5]}
   );
   gpc1_1 gpc5043 (
      {stage5_17[12]},
      {stage6_17[7]}
   );
   gpc1_1 gpc5044 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc5045 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc5046 (
      {stage5_18[16]},
      {stage6_18[5]}
   );
   gpc1_1 gpc5047 (
      {stage5_19[15]},
      {stage6_19[6]}
   );
   gpc1_1 gpc5048 (
      {stage5_19[16]},
      {stage6_19[7]}
   );
   gpc1_1 gpc5049 (
      {stage5_19[17]},
      {stage6_19[8]}
   );
   gpc1_1 gpc5050 (
      {stage5_19[18]},
      {stage6_19[9]}
   );
   gpc1_1 gpc5051 (
      {stage5_19[19]},
      {stage6_19[10]}
   );
   gpc1_1 gpc5052 (
      {stage5_19[20]},
      {stage6_19[11]}
   );
   gpc1_1 gpc5053 (
      {stage5_19[21]},
      {stage6_19[12]}
   );
   gpc1_1 gpc5054 (
      {stage5_19[22]},
      {stage6_19[13]}
   );
   gpc1_1 gpc5055 (
      {stage5_19[23]},
      {stage6_19[14]}
   );
   gpc1_1 gpc5056 (
      {stage5_21[2]},
      {stage6_21[6]}
   );
   gpc1_1 gpc5057 (
      {stage5_21[3]},
      {stage6_21[7]}
   );
   gpc1_1 gpc5058 (
      {stage5_21[4]},
      {stage6_21[8]}
   );
   gpc1_1 gpc5059 (
      {stage5_21[5]},
      {stage6_21[9]}
   );
   gpc1_1 gpc5060 (
      {stage5_21[6]},
      {stage6_21[10]}
   );
   gpc1_1 gpc5061 (
      {stage5_21[7]},
      {stage6_21[11]}
   );
   gpc1_1 gpc5062 (
      {stage5_21[8]},
      {stage6_21[12]}
   );
   gpc1_1 gpc5063 (
      {stage5_22[12]},
      {stage6_22[3]}
   );
   gpc1_1 gpc5064 (
      {stage5_22[13]},
      {stage6_22[4]}
   );
   gpc1_1 gpc5065 (
      {stage5_22[14]},
      {stage6_22[5]}
   );
   gpc1_1 gpc5066 (
      {stage5_22[15]},
      {stage6_22[6]}
   );
   gpc1_1 gpc5067 (
      {stage5_22[16]},
      {stage6_22[7]}
   );
   gpc1_1 gpc5068 (
      {stage5_25[10]},
      {stage6_25[4]}
   );
   gpc1_1 gpc5069 (
      {stage5_25[11]},
      {stage6_25[5]}
   );
   gpc1_1 gpc5070 (
      {stage5_26[13]},
      {stage6_26[4]}
   );
   gpc1_1 gpc5071 (
      {stage5_27[12]},
      {stage6_27[6]}
   );
   gpc1_1 gpc5072 (
      {stage5_27[13]},
      {stage6_27[7]}
   );
   gpc1_1 gpc5073 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc5074 (
      {stage5_34[6]},
      {stage6_34[6]}
   );
   gpc1_1 gpc5075 (
      {stage5_34[7]},
      {stage6_34[7]}
   );
   gpc1_1 gpc5076 (
      {stage5_34[8]},
      {stage6_34[8]}
   );
   gpc1_1 gpc5077 (
      {stage5_34[9]},
      {stage6_34[9]}
   );
   gpc1_1 gpc5078 (
      {stage5_35[6]},
      {stage6_35[4]}
   );
   gpc1_1 gpc5079 (
      {stage5_35[7]},
      {stage6_35[5]}
   );
   gpc606_5 gpc5080 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], 1'b0},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc15_3 gpc5081 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[1]}
   );
   gpc606_5 gpc5082 (
      {stage6_7[0], stage6_7[1], stage6_7[2], stage6_7[3], stage6_7[4], stage6_7[5]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc5083 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1]}
   );
   gpc615_5 gpc5084 (
      {stage6_11[3], stage6_11[4], stage6_11[5], stage6_11[6], stage6_11[7]},
      {stage6_12[4]},
      {stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc1343_5 gpc5085 (
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3]},
      {stage6_18[0], stage6_18[1], stage6_18[2]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[0]}
   );
   gpc1343_5 gpc5086 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[1]},
      {stage7_20[1],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc606_5 gpc5087 (
      {stage6_19[2], stage6_19[3], stage6_19[4], stage6_19[5], stage6_19[6], stage6_19[7]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[2],stage7_19[2]}
   );
   gpc606_5 gpc5088 (
      {stage6_19[8], stage6_19[9], stage6_19[10], stage6_19[11], stage6_19[12], stage6_19[13]},
      {stage6_21[6], stage6_21[7], stage6_21[8], stage6_21[9], stage6_21[10], stage6_21[11]},
      {stage7_23[1],stage7_22[1],stage7_21[1],stage7_20[3],stage7_19[3]}
   );
   gpc15_3 gpc5089 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[12]},
      {stage7_22[2],stage7_21[2],stage7_20[4]}
   );
   gpc606_5 gpc5090 (
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[2],stage7_22[3]}
   );
   gpc606_5 gpc5091 (
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5]},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[1]}
   );
   gpc15_3 gpc5092 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[6]},
      {stage7_28[1],stage7_27[1],stage7_26[2]}
   );
   gpc606_5 gpc5093 (
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[0]}
   );
   gpc606_5 gpc5094 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], stage6_35[5]},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1]}
   );
   gpc606_5 gpc5095 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], 1'b0, 1'b0, 1'b0},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[2]}
   );
   gpc1_1 gpc5096 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc5097 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc5098 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc5099 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc5100 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc5101 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc5102 (
      {stage6_0[6]},
      {stage7_0[6]}
   );
   gpc1_1 gpc5103 (
      {stage6_2[0]},
      {stage7_2[1]}
   );
   gpc1_1 gpc5104 (
      {stage6_2[1]},
      {stage7_2[2]}
   );
   gpc1_1 gpc5105 (
      {stage6_2[2]},
      {stage7_2[3]}
   );
   gpc1_1 gpc5106 (
      {stage6_2[3]},
      {stage7_2[4]}
   );
   gpc1_1 gpc5107 (
      {stage6_2[4]},
      {stage7_2[5]}
   );
   gpc1_1 gpc5108 (
      {stage6_2[5]},
      {stage7_2[6]}
   );
   gpc1_1 gpc5109 (
      {stage6_4[0]},
      {stage7_4[1]}
   );
   gpc1_1 gpc5110 (
      {stage6_4[1]},
      {stage7_4[2]}
   );
   gpc1_1 gpc5111 (
      {stage6_4[2]},
      {stage7_4[3]}
   );
   gpc1_1 gpc5112 (
      {stage6_4[3]},
      {stage7_4[4]}
   );
   gpc1_1 gpc5113 (
      {stage6_4[4]},
      {stage7_4[5]}
   );
   gpc1_1 gpc5114 (
      {stage6_4[5]},
      {stage7_4[6]}
   );
   gpc1_1 gpc5115 (
      {stage6_6[1]},
      {stage7_6[1]}
   );
   gpc1_1 gpc5116 (
      {stage6_6[2]},
      {stage7_6[2]}
   );
   gpc1_1 gpc5117 (
      {stage6_6[3]},
      {stage7_6[3]}
   );
   gpc1_1 gpc5118 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc5119 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc5120 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc5121 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc5122 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc5123 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc5124 (
      {stage6_10[0]},
      {stage7_10[1]}
   );
   gpc1_1 gpc5125 (
      {stage6_10[1]},
      {stage7_10[2]}
   );
   gpc1_1 gpc5126 (
      {stage6_10[2]},
      {stage7_10[3]}
   );
   gpc1_1 gpc5127 (
      {stage6_10[3]},
      {stage7_10[4]}
   );
   gpc1_1 gpc5128 (
      {stage6_12[5]},
      {stage7_12[2]}
   );
   gpc1_1 gpc5129 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc5130 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc5131 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc5132 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc5133 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc5134 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc5135 (
      {stage6_15[0]},
      {stage7_15[2]}
   );
   gpc1_1 gpc5136 (
      {stage6_15[1]},
      {stage7_15[3]}
   );
   gpc1_1 gpc5137 (
      {stage6_15[2]},
      {stage7_15[4]}
   );
   gpc1_1 gpc5138 (
      {stage6_15[3]},
      {stage7_15[5]}
   );
   gpc1_1 gpc5139 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc5140 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc5141 (
      {stage6_19[14]},
      {stage7_19[4]}
   );
   gpc1_1 gpc5142 (
      {stage6_20[5]},
      {stage7_20[5]}
   );
   gpc1_1 gpc5143 (
      {stage6_22[6]},
      {stage7_22[4]}
   );
   gpc1_1 gpc5144 (
      {stage6_22[7]},
      {stage7_22[5]}
   );
   gpc1_1 gpc5145 (
      {stage6_23[0]},
      {stage7_23[3]}
   );
   gpc1_1 gpc5146 (
      {stage6_23[1]},
      {stage7_23[4]}
   );
   gpc1_1 gpc5147 (
      {stage6_23[2]},
      {stage7_23[5]}
   );
   gpc1_1 gpc5148 (
      {stage6_23[3]},
      {stage7_23[6]}
   );
   gpc1_1 gpc5149 (
      {stage6_27[7]},
      {stage7_27[2]}
   );
   gpc1_1 gpc5150 (
      {stage6_28[0]},
      {stage7_28[2]}
   );
   gpc1_1 gpc5151 (
      {stage6_28[1]},
      {stage7_28[3]}
   );
   gpc1_1 gpc5152 (
      {stage6_28[2]},
      {stage7_28[4]}
   );
   gpc1_1 gpc5153 (
      {stage6_28[3]},
      {stage7_28[5]}
   );
   gpc1_1 gpc5154 (
      {stage6_28[4]},
      {stage7_28[6]}
   );
   gpc1_1 gpc5155 (
      {stage6_29[0]},
      {stage7_29[1]}
   );
   gpc1_1 gpc5156 (
      {stage6_29[1]},
      {stage7_29[2]}
   );
   gpc1_1 gpc5157 (
      {stage6_29[2]},
      {stage7_29[3]}
   );
   gpc1_1 gpc5158 (
      {stage6_29[3]},
      {stage7_29[4]}
   );
   gpc1_1 gpc5159 (
      {stage6_31[0]},
      {stage7_31[1]}
   );
   gpc1_1 gpc5160 (
      {stage6_31[1]},
      {stage7_31[2]}
   );
   gpc1_1 gpc5161 (
      {stage6_31[2]},
      {stage7_31[3]}
   );
   gpc1_1 gpc5162 (
      {stage6_31[3]},
      {stage7_31[4]}
   );
   gpc1_1 gpc5163 (
      {stage6_31[4]},
      {stage7_31[5]}
   );
   gpc1_1 gpc5164 (
      {stage6_31[5]},
      {stage7_31[6]}
   );
   gpc1_1 gpc5165 (
      {stage6_31[6]},
      {stage7_31[7]}
   );
   gpc1_1 gpc5166 (
      {stage6_31[7]},
      {stage7_31[8]}
   );
   gpc1_1 gpc5167 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc5168 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc5169 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc5170 (
      {stage6_34[9]},
      {stage7_34[6]}
   );
   gpc1_1 gpc5171 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc5172 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc5173 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc5174 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc5175 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1_1 gpc5176 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc5177 (
      {stage6_40[0]},
      {stage7_40[0]}
   );
   gpc606_5 gpc5178 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4], stage7_0[5]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], stage7_2[5]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc117_4 gpc5179 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage7_5[0]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc623_5 gpc5180 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc5181 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc5182 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc5183 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc135_4 gpc5184 (
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1]}
   );
   gpc623_5 gpc5185 (
      {stage7_20[3], stage7_20[4], stage7_20[5]},
      {stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5]},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1],stage8_20[1]}
   );
   gpc117_4 gpc5186 (
      {stage7_23[0], stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[0]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1]}
   );
   gpc2223_5 gpc5187 (
      {stage7_26[0], stage7_26[1], stage7_26[2]},
      {stage7_27[0], stage7_27[1]},
      {stage7_28[0], stage7_28[1]},
      {stage7_29[0], stage7_29[1]},
      {stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc2135_5 gpc5188 (
      {stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5], stage7_28[6]},
      {stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[0],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc117_4 gpc5189 (
      {stage7_31[2], stage7_31[3], stage7_31[4], stage7_31[5], stage7_31[6], stage7_31[7], stage7_31[8]},
      {stage7_32[0]},
      {stage7_33[0]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1]}
   );
   gpc117_4 gpc5190 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6]},
      {stage7_35[0]},
      {stage7_36[0]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc615_5 gpc5191 (
      {stage7_35[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_36[1]},
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0, 1'b0},
      {stage8_39[0],stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc1163_5 gpc5192 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0], stage7_39[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_40[0]},
      {1'b0},
      {stage8_40[0],stage8_39[1],stage8_38[1]}
   );
   gpc1_1 gpc5193 (
      {stage7_0[6]},
      {stage8_0[1]}
   );
   gpc1_1 gpc5194 (
      {stage7_1[0]},
      {stage8_1[1]}
   );
   gpc1_1 gpc5195 (
      {stage7_2[6]},
      {stage8_2[1]}
   );
   gpc1_1 gpc5196 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc5197 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc5198 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc5199 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc5200 (
      {stage7_11[2]},
      {stage8_11[1]}
   );
   gpc1_1 gpc5201 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc5202 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc5203 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc5204 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc5205 (
      {stage7_27[2]},
      {stage8_27[1]}
   );
   gpc1_1 gpc5206 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor_CLA512_32 compressor_CLA512_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha72cb0101167dbf738854b082cd636562159187ccd87c9d564e711c2c3b19ddf92868a4c2ed952c080b63d08ebf6b3ea74fe1baf41ebc7edf9f159f4325b3436f91a2bb415176faeb0fcaa9a6bbf80c9698f33824689a7647a3f52b816ceb1a18566b86a9c6c29d913629d326db3e5c48127663420cded5d865ff4ae6ed619584c22e161b4fcff980802e8f36307d1390011c64ccda22b728836ce46142ddae4629abd1a461b23ab1e3b96d9006b846f584d40b94b2227068f087ff151cae7e97bdaacae9b1edd9561c4b1b74c106b55c310baa62d1a6ec396c0bac86673d8f14aa7ce9d82fc74d1432fbf67a5001f21ccb91ac9cfd6ea9bd5c2d4ddf408b2aa16385e0376602160d23809776e3aa54252329a3485187ccfce923e938739dd2ca8eac7ffe7c8fb26a7d5fc3775ab8bd56b3b410e1ad8829e4a23a85253df55f9fc409d6e34976edec73f0bd48db4d3de6d01f75f94cdad60586c123968bce25c28d7243c1801dc563ea8bfa8333f602298f16cb99a7253c26271de733154bf3af412d71a562a2b0698f599653a0e6e0ee213c3d3fae0dcef7c8a7254bd8f976fe08ca8342ef22045014c576fa2628ac7297d665e7a2daced80311976f059f555c26f7d461eaf5078728fe33d8eae1d7163bf5a1dd6aea1a733f80908f803c0e10f46b67f45023ffbcccdec3182aab5f41112ce32dada82709a249aced347fb4db3729a31687a021173b7d03d96cb8a4a195d75b13bb7d13a36c414e5e1c4a9cc240ec12625098c836280dad62ca8d5043a12542cd980d84b2c510bfecf7b4bad8d5f50e3ee5f031657495a4ec179c61c78ac1a66c55887f4592f108e43970ee747db642def7cd758a0396ab70f8b38be109ba9a38453f5368892459690b9fb549e743cdc43d09bef22b6669269266f51ba72f8f08da1d776f7f8bb77c2e623f7df1aa2d2c60f539b3a496ea77aa2e312bc75f2cb5a28ee53f0e0ffcfc30ac94b1a35dc94dc1e372292c32c51ee7d46735d6afcee67868c434805328b11c9755638d0294435a4efbf4182ee9a62aae3cf786476936e7aee424d48da7334f1d7d7ce9e397016765d67b02f4214d70cfde2d010fa29453008535c60b02c12a1f253cc247f73c3dc114bb17fb729a739a26e8436f2083b772aa4798cd4eee11c99d3a0997bec8f9fac9f918374838435b381dfa87c739825822e0ba5c26c976e86b82c22b0ba68b06a4cef2963e14964c4c8ff4f224faaf055296908d57ee69f33347fcf5581c54c040fcbc6375134494c8def815e718144e12cabf8fd093ebd4aa34aa9a6988f191055a1846d1028b824f89a5c0e8533dd8a1779a7e51dba40611ce61e61fc42378fe2e9818998936177cd59fb3a9947816b713a0d069d8f365aa89233e8d0cc0d79b1e8b35df701ef593592ce8331bed0a6348d4f98ab7f00490d1a5f3f81acc01a8c513a869d304469925973648c63d3b9bd356ffcda973004d9ab72287525dacacf028bb4f41f86d57dc0b7499d10aed2b788a967a8c92736d6301eaeec76147dc9464c565d7cc093f69ddc6e55f7823b10d3b570ec25c0cc75be3f7cef3925fdee3fc930692cc9f90a213d693f8c382f6e31cc56321c0929828cb9b9aa496452103a5881b3eba5c38de8a9be37a9dc60d7b18240432563774554d6f8634359842551c66457fffa52ecad7e672e9b37d9cdf36b5c51f81bca168a2925970e27cca7529a0a54b4cbc28789f8efa907ce5eeeb7ef77772c75d24cc862dafb15e7c526e9e59b89ce85021935ea60696b5f28911c99a94013130712aa5de481ee8e78c9a0a078d98e5b117cde02be680ca29a795ee45332c54ce9d02fa67faa784cad353d514be196f588b0b2dfdb9036821a2763ba65286d18974da4bb9c98799ecd27f9f21711e87620242e417f5f19ec4d7eb08de95084758c9bb5d355c1313e8eee3b71703aad333cad0bc147a4ca9ca00ae3d0a91bd935765356179da7948159dc4d139a9b540ebad54cb59f2ff49d229e5ffad35f8d3c7c76bf92ac25bdec6d18c7092c0cce109441ac4686ae1afe36d68c2bcabb3f578080af8b0f6a6c97e2e684d636517cbcdcf7f5b3081c60c778e03b29f063125e64995d5782b28e4549cfa180fd184f77261fb66f53e486ab782979457efd6e93879d7ae81d664bd224871fe883283854bb6f039c385873fac4a34194219303f1722ae36afed410250f81b3a255c4ecb960e7619f21b6fab58a84548a7689f7c6dfa93f8910cb57096ecbcaa350205d28613d9c9cac6afcac38109f05faa8d4dabaf94a8ca11490e0157b6252bf4a5ee89bd9c31d37f66949a16d524fad5aea9d4f4ac9b060f2d39bdb6428c0bb63562d886779a94dd2ab58933a5a1c35ef90ac5e8c1efad9cd1fc26283e3131487fcbcffe2cf41d89d5bbe99f6619078f39cde61692dd12f65a7523d975dd83cd69e0056d00f231566ecce84f3bb6d1922333ac018448983494bad0f0f8901af36fbcfdd95db1e3c684d99ab053b3bd8d112a7ca8056b14110dd4927e4ba9f87d36c8161bdbd75efda566e1840ead4ffa370b32eb730af482e45881d2f58140c2935412f74f9be2d1f63e4fc845d89bfec3f5950f179c99bbdbc4853f4e3e0541086fe4f67d5ab0c6ebad50fb75b05f2a7652790e471515b0bc7df1968ebc22877d73165b2e8f94e76b1592807026579e1a17e85deed483647a158acd7962b14310f03d28b222ec41b34b3271c3382c1eccf2d7e9cb4845b9fa4fedf3d93cb80fb355228157c20445ef224f94ccc48dcdf665617d5d2649bf8d00d1a50adb4ae97fd89b278a1dc50581387dc45dc5ea74b45ffa67569f2e14d6af6f63e82d354c8326850e0781d2a9f8f3794d2163eb2bdb5368da7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h370d3513fd2d1b33145ebfb4d87d34c7d9400bb9c4a774b1ec672d248173bf5e74d41615da4278b35d707194217d85227e7d0c56d31640a90224fd0bbd34c02b21a2478cc340e1c08282d02ea511c317cc733c637d186c972cd9b79dea20ae5df827f93ffe346c66b10a8a7de270dcf9619d15480f6816f6eedcf1d60bb3a1dce43962595d44135c49f5e44fc22b91f978e71d70a8bb729ac984d71178447881d790f536fb61873dce8390279b0a0bb792db8faa32370aa33a8cd755bd3efc47a85efd4b92ea8ce5e1c883852e1d44ce133b75c5b42fff980597f6fc906c7c5dec8066984ae74650e6650c9ba584e8985989692785f90c0a9ff4552e04e2675a399aaf8c60b3494189af2af9c226b00d50cc672bbb5154e9d1e81e629152dc5fe52a39780531d457cd65e534427b4103e39b145102983f1389bfb2ad416b3121bc9ead9dcba0ca0e284f94bca29631f3ca424fe5b4705f0a7783f549d5baa30d2c67f30ff38a0f1f59e544845264bfcf3935243d81aaa45779036b96e6eaeea1e85001c45f4040577fb81579d80ef3e89e16d73f1b32682d9295e16dd2e3c18c64f7cc5f6b0f908c6ed2dbc8fe8d2c8a548dfc37f438bbaab36b38a0bf779c5a2b3b5bdf2c3b3f24e4f27a62a04c1233355b763e9debda10d756401e985fa98b81cf7f69e14572d25274a3ff9afa0294ba1463d9d7621fe57b75804d61e82f004afd9e9c228d5139bb2987a2ae7f38d42fa6af7e0fefbbea9173d940be347c40d0c41b8c1a82d928ad833ab6da05225fc444e4d0759e3424c1bb4e2d1d62c0d4e5083f1dfdd6be8d6120b3aa92006edd63c5fe04ce979aa607412c7fe3cdc5bcde731de780a3bc24a93a0ffd2f44f114d9328aa9186516a358d85911101d9d046625b9d3f6367b9133c7a8a86ed8b2fcb2af3f766818c7c03c5fecfc6bed497ccd724496eb1b8c5535017c22be1e1f1916e894491823efeeb095b0be0ca7307d9b6bed5af6a2a0fe1fe4f7ec22ed6d384e4122b0eb96f692af313e891f87a38fbd935f93139b56c8d76fa4cf5f9f18b0d9640d0a0e940f6c313cc3c31495c90adb48b87059964f778b5cd24dc61c327b1e5b1f9e1a1fd6b50c24544dec3c46160e1806366faf4feceeabbd669b77d4a1fbe177cd107782c6d43febebc0b8e7f38de68d2561a43ad0de2f72aec5e23aa99f2cf5dcd857d74b431ddb6ef836696fc7680de020a8b24afd6eaa7ce2376b80606397cba37dae5531dbb478100f41e41ce0f7824ada14acc04ddc4dd2ccf4957ac4d0f96216365ea8ffef579ece6c2dedc0c6daf8a1e297e41e8686efe79d84f9887f34bde4b7d751235b48f71050e1f8a2eea3fa149db15926ec60edfcc134e83579753846b9d4b89a384ca88c3403c82f57899c3d7ba806f265af2700df622e22e2907137eb9401fee065156d14ababa4cf598bcbeb878443fe1bfddf23b49be67728211d7bb8738a99b33acb6f432215c89b673942662207dd396ef78859aab75d0dcb1b32bbec7761d3ec5e662fcb4f2814f83889ea75190f9db0f8ae66aac266a0530c7b86e62573521d4012e5005b6fe92ce9b100216c691f6f20d2b16eb1e60ebb80d6737c0b163e24cb418d3f9605ebcffe43f30e08487c209fd03b53b6fc123a688acd49a7afb891097eb6e03c7436e1939d337b585650f6cec93c7f5bb8b350912f5a0ca3daf2ae864a1c6f54a3044a213d0ad6f71f63781414b16bb7f831dd0bca103276f50aed1db925963475865752a2edae445e0dad7c96dfd30c46f887d7c960a10f9f6a3f8d907dea49e32a4cc7cee356c3f13f2fac1f01c5ea394e2853e64adbd84f50cad4123f6a1878953062a8fb7b1ac24ad1944adcc21095aab3532e73ce59f1cf38d8f48b03d64fb4198c53741725478c1ecdf629700cd4bcefeae0c6dd2b23be978f2b9ed1ab88a24752c71dc5998fa602b08446a691255e9ea94c13b8329de297c92c1c9ba44b5f56a40acdab8f2d42bb95c693ce33c22722f230f1b68879add3d7af46f24bac2d99182879cf03006cc0eb2fb9fb8145b3982b7e3efc82bb5ba19af2ef59f8c1ed147b89b75f608503895d968a53d8d16382ccd447a27415edd78007bf76786baa8723c783769c8d05b7a4985f719675955fbd2db320c4d17527567f1d6d50ea2f9179392dcc3fcfb3d9f4605fdef21cde53dcc8cff79adbc9e4c1dafb1d695a3a449458d89ef010a863204d31f286a192c1a58434b55d41ea9b7b6b6e1233e50801144ee3c90af68c6b8984d574aea9198c08ae0d8b19cc8c7c868d603f9b16f44c6383d63eae019de0c9818d1d601e26bb0cbb32977f462194f546bfd7dc57f0cfaa9aa20fe95e7ea00e9a042897d6d6871512e1d787434591cd81c04b1672f47614c17d3381ec772766e04cc51f13b700ef72822e095267dc24c7dfd5f11c395ff19fed47b8bb6654d297ba35bdc9c2c1b03949958fa01d3d36999ed6b7ad846c25572052f01a1c53ce7c1d2f12d92ac6ac15067101dd088a79662036c991d3eba91acec362cfce24166c968346fd12e6e8142043d1be15c1593f505803084e081fa362104649fba305d0be1ee3e00844af8481784a2558c7cf70ed586f02b321b299bfbc910e7e5d7a2e1e225ab3f893fe867e5739bea957d69b898396700e16b77c2f9ff27abd36569f2b0b5d518ea8c12d38913680dec96ef7ca07d041b884cbf04f927161f027ac9952b78bc5691e5af1d0254dd41938d3b400906389502352d3cde0968925f22ecac14e8fb27e89bc7b0d323b63104013f3edce89844de2806d4f8da55b129c33de7d150f8c8e8392db405c98c77271450a23b2a7a12575b7aaca6db47ff1cd884ef96b495415b120942c04942de0a845d410;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h24c24bc1c72cd4e295e85ce92a75a9fd6ca48a3d511ab8053eb314aca77495f0ed87e8e90988e28909d9ef5aacf3a0fca3afb033630b3921cd2cf660a86933bf07c71a9ffc2020a83363b1c4df3154c04d30cdd46bc610101e2b442a8c7458880919e985faca30165772a4f4b22588b9c26e2568c95766cd5ce8f3ed5a8b3845d9bca9673ab8e192c24fa593026ecbeb36e6a0441038f02b065169a04437a527b5cdac74fb857a23e86cc1ed55ab9315955a10614b89f48ed615b7d73547aa21814bfcfcfe0421ff193bf9d0641fd9281cd282262ae85370c912452b5da39a9a8a7dd970a7f45ac538d0a01e43f1d5fc4985ec0f2ea2e2938556fd6ce995ce74f1dd68f89e627ba1f568100aaf4eb808bce21b1620887b4e0fa6276495cd7001fde89c5aa801c3e77d23c48a0f49bd9e8547be3a3cc0c1aa34788a2c0c2bdfdbf9659aa339b0679bdf20b40f7aaf432d4f55cc618a5b6a05a0ea0b0bfff61f5a06673c6b745978302d30226773146129ed4b7825fac4d90f718b3920a1fb19780e7eb8587f03b15a82a864d3e5a10fb098abec86e3f655ed3e31e4d2487b2d30e92ccaecaf927b3a805f393c2160cac3e0dba82c997d3083e3bb6b51fe1c8e708df4b57bac271da8f8a744bb19c7b72c8a2b32c8560f536bc23b40501daee524d888081012bd68463632690d0aff0a5b3ab9e216660eb24a3f1aca2f5b75770ff0d068e92c67bafeb1e4f05716c31d2f08e8063c0a81e0123831f813eb95f90c30a4fc68bb88e7d06dfd59d3e5ce14ff1deaff98d6476b2f9a1a29d4662b2f3ce92c7c6748bf2081d4212ce6d73aa0a79895f03e903456749b72f471f55d75bc25dcb26e33a6584e08725b2dea244123924b81f890a84c0059fb7cb81a941c1f544c416b90b003858610c8eb1bfe64c9e2ad3b9b6564246a310b7f93a3c820c235d97d25a7196d683b88f81ecbfe04d00627113383b2a9259ec981ca1847278cd5a478bb19c147f054b621a86e16187f3764de183a5cc6cf77f25ea9f6f6567f15e2753facd1a44ad2bf63e8e46900daecf44b4f74f0fc70dedafacbf31e90733da9be8600b8aa2f39cd1e0e4c64707e204184c66ea1fc386640fac2c0a72a4edfae4b27f55d1e99d730a54e8d967238e91f9904fb6b20dcf724802f4248c0c350fdb3ca0d95a829f918b5f3049d82173b3d8200f7f77fbe741babfa41567c7397c3192aee7f4490a74aee10759a70b64bbc2d5bc66bffd97e78c76e1b32ae8adf999417b732e6fcd1594ca21e24068c89c18a13086e620973a02d1d8b9f12955f36ae9ec284ce158b7338c4ca435e745aa781c56ee01d99882b0c4b45625ff80d29ed75d1ae57a7a1d0dcc680f40552c307bd15fcf8b9ba6d11b0054e1194e14021e38c523500a66faa4d7ea91f7a0a8fe155fa5637fe3b59eebd8f12cd396282b71e933f4504ef86966b23aca33bc18588cc98430166669419d28a75249dc50737e5865831454b4b86128a5c0e4913d59f2b8b6d1c9c052dc69741ff2b54e44a3898c0d598254f7b091d6f32fb4b0ad67887a1ec4d00200999e447d385579febe667166ae0b17900ec92aa9a15a1161de4490b6989ff2da8b830a76355068a51cf15ce98f93b77864758f3c6467adabdb4bffe35c870ab47674c60fe3556e9f41169202e112ad0bce121b1fef6b236a5230b186517673c91553a8ee3c2ff583bd83207d20b0f90a8dc358bc6f093802091ae040d493a0d1825e6cf94bfa6566dfffa5bff4590e4a70dedfd7f6c588bfd4100bae29faa1daf9d08817b107a9ccf55e51c93e31d295d932486aae2470d344a9d2613fc02a8c95f19933caadb1d6aa12610dc5545c9bc3260449327acb3aa51097bfbad355dcc8161c22d95b82ce470324fbc44ef87adf2794e89fa69ff4dd9dee4e99b142917f16665ef7ac833c087ca13f2633b6205d435de5ad8477952aaed450607a61cce6f0da9caa314d9414855e5fb8b8e203a4bdfde134c62c7acecc50e4a6da63046e415bcf9d16f2683825afe303f07aceaa826a82721ea3c93533fbf9c95628113345b9b9057ca3e7b18d6e04d2af9dd3e2c96919fb8c0062f3dcd995660c7e7c7e7e82306c18da7a231c45455aa6e2601aeacbf4a3a4a36a6e844ec0f05bf7f3b92b09a9b5bd0294a42ca481b976aba4e1b610bc30b2d14830965f72f5c7e1baf6cbe56874dbf4e9aab9bfce3f46924784550c33722197f710bca3fcd5a2f9581e4c7cb0f17a79448048334c0d3001d364681cc33b15de9595bfe493429e8413fe7e04c5a0f9d3dc733c5d36561e6fb33b710c4ff28106c2972155835a75072ccc278d278a4bed1e9d975f4d5ce52fcc786882397360c4cfb46e94e8a617acd54068127325af5e68294ef6f6b89e897634b7dd57e4a5a55cabbc8d1f0fd71311d8b61e34610ed09ff50ca5bfc79426cdb3c1794d45df47fe1043942c6adef8be0a7f439f71297c504cea4cc0561bebed780ba693bd3b234036d4f11b49d2a65d5f4c75536b27d5e9b000ed6f019ffe17ee5ea2535997bfb7349a7fc82afdaf6df30accb61cdf53bbd44d30e726691ba58dd06db5789ce8286d4657fb734d9b188e5e0b0a97152508e7f8a02831db47b5e9775d0da7e2d9e0ca648db0465aef0bd3a89da27684f9e0fd2b98223d813a23364739370bb3124191093766ddd5d35a3c45263ab4e794e17a0215f956047c5b5d864f44f95866f518da710e6a9896ce21ce67addeb5264fb35520cf3773992a547eea7240baff18c3b89ef4638f2b674e85586c31e9bb3330c6993b1a3f8a029653c10b0699bf6149b1e6b2acd0d633d8e6fe779e07f19fb70f337512abf5abf5d2eb57355cea4d347eb7ca5424d71abff019b1406c0b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd4199da2ba7ab4fda6af9e02200af91fdc311ea10835d2702b66eda6b8d11ecd1571681559b97584b51fe0c85f1f7a765e25a7fe4270bb1570c5d683ada15ee5ad8e7587ab90f086edec1e731f31c387cc86e22a6b9c3b519432106023cc500ed928db259fc001780a7380272508a42d8fac6870300e501197d0f4b702fabdcba858aa19817b731daa39eca6c0ad0940c692cdb8e43c3268dbb29f60bc733925deace3d3aed7c5ae0e465e21b5b5e67bafecd99cd5ec5f18dfb1cb84615d8f401b4ad7bc93b41e079844c980adb05276b2d3ba7ecfdd65d857a675e1b1e5bbf332b74e00c43710efe32be9bce4e0ab2b6b4dd88b30894d654de15b9a23126dfe41a5c2628adbc792a84e6c27e40b7895cf0c9c6249a00f51945904adb27e0f0e6091c3062daa49073e5c6bd0a9d6753af373d129dedb56d3643f54bf0e3dc5e22fa366c4f7c9ad027bfea39ee57e45ba0c9c8654783cd527845819de4b53206892f0f3e876c2e45403d58f43fd0b190fd888a54995fefcd2f7f76d192da173f5cc98284182c9056fa32465a8dbc3bf3ef8acbb5afa388ca64f0e27212b3f694b700f862d12351227800876596fb3bb31b8bec0efe65026b7437d366ec7b223bebc9637ded003b768322d0e7cee0b13bb52bef669e8a80c64db903681535b859a1db223c297449bfd7e7f23dbb9f1daa6ffbd8a7d8e53f8c7fdc06ea40a4002830101d32428ca5500e4cd26a5985c9ad0755263e23d0db22e1e3cb843a3b16e0b4dbed18c1148d862640e50efd1e778a59b998236d017f2c30095c52ad7c6cc872715b4f4896c41d0b541c2c53dcd61bcef5f4230fe1ed873405fde63638283774a6243d4ccd9298ff0d68dab840ea0c752df939924c32135afa71a3beeb73b2f3d66a97c3687647cdfb8a0801c86a348ce15e75eb2020f2b19de0ef11c8ef84f6d08325eb97fe6c87708b1532cac2252a0b13ba55eb603089615ab195af70f0835b3a44561fac6047e55abcef34590b46f9687eff03c6fdfdf04f4e25496350d62cb82728b58cd019ecbaaba06095208e9d518e15169c9ee234f4ff057f455b55294537c3447b7d88a68e3ef5971429327d6fd5d293c2b426f63124bffbe43071e4391a8f81bd5def441279a91f235868c4d943c2dd9a3523385e4df28f45dbeb8fe0ee8c1cf1709f44ba545ce8e95620907d44c0889e5d475e64517b899aea51075e4b08af6ed22f4adbd4afbed1ab82990b5e954a2d05386ecd5cde83454f88d5b61412cffad136c24400fa789c1e0dfee867af9375e61a29d750c63e020b7d979acb1c754706a2306d180a461bb2dcc53300185eff67a9345c553d46a5f2db38c77cd39a7a6b296b28bd48f18ba1fed0503b7d1ed312dba45bbefe647ed481283531be1be6dfc5700d11d42c99b422145b06ec01cceba70a3b61473b3e4bc2722a5a35901a7b6cdae54b9e68938b4f5681244bc8355870d8527198fb2b1e317219fc960a83e07391dbf7254624df98a4d7b57cccf4337dcf34ad377c50ca3dabebfb6a04a2e14c9bd423182437830a7f3c0ec5a1fb34f13c23471cb151b0f9ba280034c1b33a867885644d8848baf14f976147f1fa1cd78739e14e2cdab2052843ee5c22ef9f0cf6267d0b3479befdf6ad1675de72ab54bb129b4c56d0fc1e360c928bcf8ecb3bbcde793630ce3fdd3a889408006ad745428b7d64049a4948ca9e651ee29346cd2339adece10b0eb8cd1d918a759a34c537f7faf4cf817eea5d6393cb1b13bf08194e3c8504d4a49c9c3d08195b70dbe79aeee0a0ffd3cc752d08f20d7021778c5e82bbcdfa81a9a49e5dabd17eb79f9285fcabea3784149ccc787c860b9090dcea3bbcbf9b6e0a4c091b7e8ddd45816020fa14fd20d742820b1730dc24815e8f937eaae422f1be012ed8d0da0ba84cbe6bb788869c7ef164580b1ed1d31062c15eed26a244387315d2c64f58a78c92b0cd04bcbecd096d10165adcc5637b5ffe38ef2f29f888c862554e9ab98350e9631bb37bf71858f2eecd9a0dc011b6601633d96f21ca384a389bb0276313e5c5a875f25d4dcd3caa9216b663453bd1522c282d7779116fe8d92fbffa60f46490b60141199397230ec9209f14d593979f1d64a3de4cc05a729fe10e1a9229a85dc6d728f4d1982681c95745c9948204bae52b54a3453cc498cdbbd0ec8e7c47350bcb0d5c2a0ee144c6865125ac396bd5e1d2e651acd510a83d4ff22dd43c66fbbb682b6b368a28134cdb6fd268f71462d2ba489d006cd84faf866d604f4c44f588f08a30f214207ed42f99f6949a48490b85f4eca3c361926c77a9a76f29ed5557ed299c56d6ae2b9635d21caac2a9f00beedfdd69c52df349d4bede81dead92ff361f6c708b3de91a2bcb67d8767ee58eaf9018c9f383472022d67748b98d19c95d1d6fa503a5f1aa9cc546130c74636367447801ba50be5170d48e49caabbfbfbbeae4e546459488c7462359e6c921aab9fae9fca7139b869eeef16bdd1836fc2502cbbdb533d857b0bad30390ee68e3dce112a0ef7efeb418eae85019ad5f6102efd94e802754d1a04a884ed7dbbd9de2ea159391ae929035198c83b7e05b9cca4323c7ad3af6e6653ec3e411d46ed711d14c4f68982f155b78837d029e0239b3c6904dab8af71fe7e57e39be09b371b2f6816ddbbda8e15fef581f36f40bb594b310c31909b25fe471850085b90f1a30d52dd0619643b68336f8ec7bc7fafbb5fe23e7b5b3d32825ef08edd0086eef339b3663f3dac87fb114f42272b514cb8aa237cc37fe1529231c1526ec69e02a6f06ab511c88403968ed1507ed4c2a371287f588918d7d39f81ba72201e3b6374ab93a5ef8eecf1c685465d5f1674460c79c67d2ea1c31a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4d6018e3ac80fc0ccfb67764a1f57cd26c968bb6ca6a1a6ba657dc3479e3262f6a396cd2414aec6fd11bad27ec5b7b5e5de5b7794b01900a966ba560a87b62bf5038d8ba94f6a0f9eea8f939bfa082233401fc0d51aa5d01da0e69e0e7d868927123dfaca59a321cc158f51d281f22f8dae71479e184a12c0c5622a96736457cb37bc0620216d71f542d80575190d0f93ceed11dfd7e3264e24e74364f5f440a401dc336e9f3e8f7571b952f515ed5f67717ea37b421aea1dfd909358b0e4945d50a8a351175c6a10fc5da2a07c1561b0f4d41686db40df6c3c10ddd508af9e79b0d7c9fc280003c752d861fd183cdb9ebd1f57d32f12a420db8ba7788a59668cd194c25c2b919e2f5aa73f1c3eac7ef3e063c8d58805bb5e2805bee5ae58d198a745fc10a3cc7efb9109076084678d77f97d01bed76e039531a29dbfc63e7dca791d77def4151376284a7a010f6b5dbc7cab35610b41168f1622644f1772cc0106439bfeaac566a49c8505ac796296a5c576d12245312e27a888763cc9dfe92329cd32b03ce7cdd639379dbc695ed128e4aeb131131febf003bc8842fa77a065235e7acde66b4bdc70f7e5ddd77f77a9051a7bf38b15716494e8a0e12a22c90bc0ab9146204d6f00fe4a0a2beeaedeca0c1e5f996cb15c6e35ca2d85a80321427ce102fb05eedfd06526c8765ddf88528e1e80220aa76bb42fda8e1bc199a39e9504c848040243e35c0a3db6d0705fc1d9ed9aa29784b7a6ffaaa415fbc734d2c46b652c9d1b5a61d54ba7a73d406c9f451807dc0aca83f93cd2dca6e7edb45ad77ccc1fc923a89d194b4f1c94be0c72767556c7eec805f64b9186eb70e01cafd7875c3580763ac2e8d050ace5ac7ac1647a6484549876d35464c1359763f8ffd96d74e2399f42d174c633672fddb90a6885aab71abbdd90bd9a94a5cb269e0d98407a618a2c2d489cbb0073c8659033129a5c0266c16926d97a57d9ca13d1d41a55c200c9dd4c990b7cdc5c3aa1c110f28eb94dda24d2aa3c972ab5dbcd2ea4f7c37b8d321b50b9da5704e98d3fd1f8239a9f3bf2fa5ba5a65c381754a8819e96a95d327798370940f001657978789ffcbec8af01a3f84bb7348f45120ebae053a3dfb0d58cf94bbdf71790e536efadbcbee60e91eff1979fa6f9535eb99dc7324a7d68d36156aa1856b7f1cb03e82c923f83bd7d93c837f1b39be02ce05d0b0bd953ce2eb2fa9d327fe940fe0d32ec789134309d35fa9afede2b8f3746e1aa806243122cf00e7f89751cea470a1d40d6c3310743b5f5eefc2d7390841873fd712bdbc7d5bf66a2e6c54f9da6cdc10b6f69606b9e50af4fb24caf7228f4673c54c96f067ed963a581bce915920472dad0af89c93b2728d54893e597b4a4fc5cf3107bf8d062da9cbba17ed6e1fa0c37bea3bdd00900b3c252090a7df09778bc3a26b01c303c80be60129eadc8a34736b30c67094ab90f47bbf02cc35a35765c7737150efc02f8a50b44cbdcfe657d959fc5383387243bb21d4c50b0bce9634ebde0cae881c2c8b5b316e134e276fe2d8ceb908e37797e185bdd92787d3e59e45c3324c5bfde255e3a0dcc8c4d0a947bb154ecba2a21bd9e335ed191ee71f8eac081fdc16316e085786774962d0fdc0cc3c832aa38e49e93037f7958d8034977f08d584fe826e006b96e6ba35376879c67c7ed9c2d1a006844774442e2301a183afc780089a998a4c9c316e6fa80604968f1b336176974a1566490ec2fe6537aaba38886e387fe7412f273d0cdaf9b992fe06f62cf88674f69b22edea162d93180aaff958912a0d85e17a001003748b26a0cfee7d39a91470e11786c3b1779db3fac4c7b33c902272d2157ce2e24e8f3ff1d1a6912de9d7ea315f9b9e1205c880b14543da6b486cfa0485e0dffd78de6ae467f35d571f5ceccf76191dcb72c2c87f17df0d34b27bf80bfc392e2f1af5614e3eb57cb57676ec9d2471823166765350e2a687d3cbe1d95ef8bf0fc25036654dff8d598ec5a5c1e77b36b272dd88d92eb9f558f3a702521656fb5c1f66c75e2526c076c421d217a9ac9b3891013246e8edb77db7b0ff7a11727ccc1eac211ab7707379aac69fb93da60b298e38b02a31641694b0caeba86a408c4bcec060a1e07508735bd0f2d30c33e2d2c4cd40d9ba50f936d97cdcb0de8687243f1b054c2a9104e96b6399e7285fbadb72db28b3c7182a16e42e60c6939dd334f2a1defffb23d3ea8f56acdc85a64e5e69cebc0c2bd868843cefb1d6ab4892ff4ade7828daa3b265a187f098f27d63b0253e3ab6be432bc83c9f23a555ddd703be01af5b2103c42179cc249a9dd2924db79e3eb37400ff3a0a93b0248839a1795603e9968ab788929665c1c4df1aafed9cf7d91ffb006c89222724a4a059f8701bd1c79e83a23e416c3c4234d9e1c4bed1f39f864f7d84f7548ddac2604f8613bcd1a1ce997677720a496b797a49a441affc9282f048b6777ed06b56367a5c68c8933d55faee50321520085ab0eda1d1d808c3a525cec1479209c43c78315b76178bb0e1cd3259111404e9bc19109a13352e327837ea34354e5a85fe7d28e0148a0af5c8d2cbb00f580e2cc85772ed633f28b0f6c3687f69820fffa3d0ba26e8c6f150dec901387801b00c26b952b61358e1bb0a61b86b5cc7edfa5de9eb586949f582431ae896d0da0fa99d8ebdf35d4c1598dd721be5a19c6c6ac9075306329f02ae244ddab8c37ed6764323cbbfb6bb091636ddbec99569527e85e85566dd14dbaefdb432d8e92c3a9ae4ad62dd6592dacb05d7cb8231d27292d867320223b04c43773f17853a4bf30c7cb2798721149915a4f63bf48c447d038e08c05f2c4586ef1cd070470f1f778729bea877bf396dc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdba7798466ef7ecc8a0099d481923f52b8e7a65c3c1bd5f679ae69e893625a2ecfa9e6b3af72ec6509a1ed212bf0e8d3b756c73ccf4601ab28b5c8e9b9e5b702ea51a60682a39df152e80509bce7ce5be55620f7b022d2a9fe23f59f931d44114b209910de17b4b18315d53a8b79ceae23a9a30752815ef3fe5353c90850c14fae4477c1c6cd70327b8d8a4faef2544ec8dc128a1ea0320343a248d0bcd0d18172dfb64acbb07821fe8290d64badffcd537bd95c515b236375b96da602a13a9b8c01f3d7219c63c2ea097c3042288887145f32e66d07f5be6a01913cd1002f379bc21fce1ddbd758ec70893ae3b24ad0a0a0ba926d2bfbd4d62c966eae895d26c077426a21c995f1299d7344dfd001e7781cac8f207907107b021cf35d5ec91ff7906a9438e80b9148b9dd74d982b5cff556b93fc221179bba248ca3f633c2ad8b61e01b4e3fa7c6f3586ac2cbd420748beabcff1f768831865ad6fb9714b98625253ef441e305dcec9f8778179cd0fc694e96a9d0f656d037a51fb185188c26a441bf1a2d2ccc27cabb7860e5879c3755d038a189eb283d4e8173ff1906e10e959a634e47c74347475241ee64632deaf16bbf37b5109ce15efdebefec802efe18fb3e42f035c7068faccebf419ad80677a3d40b4e0d9c61ce3bc5dda0426e4b3cee870735970f1e7fa0fa7a7a5b674e85f258ac336bbda8ac83729117c46d9896129c76ac2cf50b0188aa0964c7c9b8a7ae901784fb9eb1f58cf23cc30c7a238397ff5c02472b4a4f203d01c868234ea9ecdddaf6687bd3072e6e38c659df5bfe0a74902cdbf7ee6b5c3ac81533a07c61bec0f9aed68a9a3b9227eedeac85ecfc87aeed9cd8c22038d059b7637bf62f1ab406a6f35462ab17d96e41cb654588c21589692a469439d5563f952e8177edd8d508a49cd35200412e8e10a2cf1f4e70bbaf85e40ae876d46d029e57edfa962619b79aa43730fc9468c6e0c3c00f4f0e80aca3d6224ccd4582ba24fc7c3c4badff9164ca35a390d3f4bc793b247d69576024fd294582c43871a05b61f1c35d288b9fe0285a9900d6f14e8dcbf6823dd438af73cd4fbdde1b20bb10c5c2b755f3f7a8950e9a12e0986356e3dc987aeb12b1773bb872633344ea3ccfaf836499d21007fad40f9465c2d05bb4fdcfbc4ad3b7a1d665cadad33423939839f813e95af67dee2bd0a7439d7f526fd17465c0ca7eb7700b9ae8d76228bc9b7e9bf60976af2a9796e5e574aaee4be0f41cd54a6f38af99c7aadc3acdc6f261c3346fe48b8effea6720e82e773db9011a512e2a9912f408ce95fa73ca6d2f2699d5814c8d76f30d7d55053eb469cb94651daf890b73cc90e186637b1eb8abc58cffc27c9842ddcc5e0f315a0d8aeaec5eebc592715937b9459c3c9d0a69e57e35ed06a30a24f6835fa7845dd01512f33d6ff556587ecda1e2bdf51b0c2c105e91f577af9f4a1401b6227f91eca5224662531ad1ee4f31f92f370e7a6f4bf5824ade9219bd2102ead72edb367f580f889c7e62a9af125eb43d7339d68dc8a667ac1b5f46d88087de0bd339c68acbe29f019f365e89c750bd4ce5d549f3c8029cfd98829520b92af2991be5b7274c2380db1afcae379ce27e0b66ad0e11a5440e0b1a4ac0af398067e650173bc04443291f9f9343a72dee3af217816549545161ed47fbfe8d294abf8b5f8c5c5f5afcb0588bf95c67544ee788b55b9bdbee59978be0d823b7fb9b46e8dafd0debadcc63332f922133e9a56189887b2549d886aa294a59c4417e457218a3b80ad96ff5d33060317cd2a21c2f1e7b70ecb22d1b04d903fb20f05ecc421a18520126aef65e168234c3964d4bf49016152b50b3b183b958d25b7e410aa85c561fb3e7d35d05ca8bffdc63c0ea88242400bf793cac3e5baa5740b43f020c2c4c7fb1f536215d4ba0d86ddd060dad22e29759ee346d52c70def9dcc08027bd2e60ad67dd7faf263cffba7c48d156e56956cb7686df863057cb798c4d53278611a369ad4f93eb7c2a947cd90603c63157aa5ec70321d72242994d4f9aad044312e64c91ad5f344a796cd9a953e477942632f5418297432d1f52c1c6b9a92437bc98e8222fe97ba12522ca39d528510cd9da70c5c7a419a056a5ca4be6f99a0680df765da468d67accc346ed562f36dc9fce7efbe7321d3774ada125fae200f79959b9ca160b719b971c9e49e20f7359318d99f8a8911e2ad7a24562400df99c48bf8a6318604f7bce0e931a26ce1dd6626f691c7549bbaee4719da23396b3f547d54be04e010b16f9c2e1fb74ab6f388066024c4e014437bc02065dce922b7917db28231c24abb898a4021d3964d495ffa5d0b9ab6062bea7b6a53eb74ce9f8415c3071dd1c4f79ab34815bf5c9dea18170cd2e3756cd4e14b633d0a462f5c1ac7c012f0cc7f69e3af65b6bb4391399051eb3c319843fdc5afa8583355d0a48a864f1698ec1dfcbb5ce22a4bcff8d042623877ef42f68eb6cc1d608f311c6ebc5cd5d465abcf09bf2d47402264f0306c1f4f464b7c3403cfb95e0cffbb0aed260dfc0fc4e8819c1b797ef132b84ed9e3eb0f1809588081379039b072429c0be9b68999daa6bbdbc80c2357a36116430994371ebcd96b3b31328594c7e173740122041d54f51cfc2fb3a2759ba24994113ac4744024d27929732fc289997f88d0c74bbb0129f33d6886695abb3d63775978f07e92c3430b1c77b8a8bc48ed504a3a3931b6277f6d76d448d6089b0a45fcfd6d8bab59f21278b89ac170481dca98579f23d882e68492466da3a772c095e0aaa0d5008f4dd9b383167245e2c3ca14e9bc3ad0b86145f0f711ebb798c9704b3d359f8f65e5c377f532b5994fb1acd063052c51c6157f101241f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2b16ad213225b7eac9194592210b92a5838f78e770f5c7c0f902a5f8aefb983d6e6b0fd2b6657a59f544faab10f2d07316ed908943119c8fa5c3ec1b0913dbd3967f67019c324363936d31e208c413e0a34685974143f47049e887bc6f102ef7d8887d3bd2124d5968b40ee649392bd730547f40a7a03205cd9858516d73c10921ca22c22a4957cc1ac0bae33466e4c3184fe83d1051f7bf465bf2f902e1b7383e3093bdb6dc2c47cca8ff90fd86c11df1b878ba5e596afcb046065bb83e3a410d3dd9bc746a237d4fe0ae3765e9f80979865abd9fdd8878b4cc0165f37b90106086ea38d80c36afe79a3c074603045bdea9dad4f07efd3f79764d6895809dd777592c9e786f8239deabdff8e49b4c25b316074eabc2d997a10b555c9e6e456cb52d7221b1b4044d1e8bf5018d36601a8d5ba6c20623a64e02775a7ff969ab6c3e81cdaaf67d7b622325740e6651eba2b8eb7663b76ac63fafc5aea9cbbeb47f9fa059ad3701493689841c0f8ea1a24027333d2f7a67f1adaeefcb983e1921bc38c8e18dc9d471d50f412e28a72e78de13140b122d04a31f3c3e0d377c46c1102f3d129c0afff99fd75d187ae88844fcac5f8e1215aa2d3e7f8930bd318b6be88dacc6d026a7e11d98c04994700b08dc2383678050cd9012eab706cbb060a32ae97e0f1e5b925875267c08174908609a1c09a8ace2613117614bda8afcad76927d0571bcfa2f8050f25b2414bac345c2435599a8ab7eb1448c7338d1892c9efa754e439a1150ef1b91b8e037347e72d6521c203070693f99a8a6d219d78310aa868d7ba465dbcd40d0cfeffc58bf0ea037123c95b12c084696603a9214d3ed3ae4a42ae9282da01acae859d8d72f1836edfb8e21fd5288562d90387a0ec340bfc19076339cf2d245bc24173770e6a40d0248e96e684c673561f2ea9aa65af960354eb2081360a859f432671013df558cb3b9d1811804a86ba4561be3544cac4bce22567b776bcd42b9a6ecf6707044ec0112a8491de8849f83481f3ce532d7355aef1562a1576b1b2b1e5df71abbe96972f0dbcdb489d3c19ba38837bf1542e9d35c50017d08eb1d6078551f5b0542806ee427b8d33136c2fa440e65a45cae9d9b7534155d2b372506ce4c5ed2be1c09f574ea0360122673a8bfc19d5a6274e45dd89ceac45081614ac5c7bbe1df072909ccd0cf973e9e9127772c99d324fb9adfbdf8f4f61c55164cc3600ab970a7dc19747e0368076040ea38a776baa9760c7d5fbe6feb1c7b18aaab5211425e5d5b878f30a6d1ebc290227b0f3ccef99d5977156f41579ee727f5af3199210506a9a9886a4ffc94b1c17c72a3e7f9ee6849b60dbc6da80372cadaddbe50d91f4108ea4587c3afba1eae7077b785a7f8e94d5f27cea4aba89ed281ae8b5f9f217ebe3fb66b40307e6e012ffcf34bf9799f66830eb3cd9ce9aad4194fcf627e3c8b4f9f769ca5ee8c33b08e12d57b71b4c78c366460aa3443a7b4af7ba509b1ac3116626ca4c176edbdae6108047ca53fd3d3b87ab84cc3dbef300ec3254179ae3c8374dcecb81ff91fc70bcf519d2508adb71e9e274e5480a27ea910a4590be78b0d1351178f600f8cf74cbb334f6321fa7d843cbb901ec25bc283a29dae4a212ebdb3e8e2c7b091f337780926e30ae3f8d8926e561fd29d653d65d60305665bf6f7ff99935f4d2a903b1b9384b97e8fa99da966dd06d47d00d5613654394460d783901e0a9a81062cf8c77d05efc56543ec0732807bb409af27203ad7bdbef2200d89e1c461a8a1e84dcec42847e6e146e1d1200080a4a28d3471f7bb74f4b2a713058fef1f7af140509fcc8a3f5c9bf3b9129fe7f2cd1ca55fc4e1f422f68107222ce748de6034fbdef6e31a3e2fe80dfe3ca34f226c5be2d7987765f8b8178fd38f828e3297bef0e9b2503aa2184398b10455c2e05ada24141d265c41fa263d66a05a0a11714465ff4405f2b2d8105a3456bfa3fc50d37f8d65ca30773c78b324226789ecbb59c072c541e6660c7be4964ae109420a42c4fa3687363c19404dde830affd009770a33e1ce2dc7e321868df936396bf3c4be44f55a698f416531ec8c50fe2d77a013318beeb1ae648681d3c0b2c94801b68707a0d1183f3bade85cc1952a16a00dded4b551cfb21be0508f18e4d8ec8c7aee51d854ca6d5fe699486528a368193958c861af1b9a7499d3102ad1ddb2047803cedc7d36f0f58a4b6fa1a4e6fda278fae4060e7a891c16fcdd2919735cdba07539b25d2877b34dbd80b8c356d575e1392213045e1a6816feb271296f65d24143a35c79e7f0aa46899d079e74b21394ec6d972a6cfd4dd86dd42e64c9a4c097a2097578a7f7590a5ea759259d60ce19ccd7f130b95626885b15069f6a046c25dca1b3dda420183c1aca9b6ef141b37cf13f6b316f09da8d9e93025a72aa6e81b3c4a54e49f7c3ef3aa3a96bdd9d44e804faf0a13106e8b332977e92cf035cf57f131e59e34656e22d50231ad56f393126ccddb2effb8ee4c0f0c217c0cb5883980d6ce6bb05649dc36e4e393c27a6e8e174e0331c9b40bab15a2749622452bee44c03bfbcd9f39f9122cdca70f9ca9f1a23d9fe2f2756e76b3bbaf28fbe85f52c333bd1ab78cba0c54cc6ce189a0415ffcdf094662a22d08d9356d2bf1eaa0c71fd43c2f22d13711835c62a92886d5755d51b40237f2a6a33081c35de7c754d4e392f0cbe3a03e7e00621501f0c0805f7abc3219fa78a762cf924f36016d4c35b942aebd02aed37adf51a2a40bc0fec1847e78503209cf0912432202aaba2c3c3531bd5861389194126503d646ea4df419caa5c06b78da1b1499ad42d6ced36df98a1ce123a4f83d9a0b53405cfa115c346744d9e0bf215e67e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h84d9ec1c6dba43180320bd9790b1cd4c7941c6983bf66ee02b2fb6dbc74903c8cf411fb2038dbd6bab4de6334739bdcaeb02c70e877583f4f30f325c8d1f7bb50ad04cb6fc069ed4a11ae5965b9ad27e99df0a173a80fda039fce179e4001e194883bb99da0d65df4e2fc13d6c7170b9c4092534e913d3ce1b4ce4d96e3172a712aeec9e6758bb9f87c1c5de02cf71c7e51cc6975cc91be01e0c140a8bfb548c9a436c10c1c5184ebe640be04b5e3eec780bb3f86a7523f0b65a4bf9229cb5ca35ffec6f26fb5db8615bbafd956695779bcfb0adafdeb484026ea4f37b8acc523a27ab25930b6e08237788f3d71bcf2c0ebd6ea6c7010f925311d302635e631e6cfb31df01c15638fc442220f807ed6bb404e7b16a6eb86e116e6d733c55126593dfe633e894042a14a34efda4fcbc0bce97889fb2611c11a89ca13d3d8e716802813da6358f2db4c7ac9bd00567c7eef915a587b5d43388df7d576c9afe9e1b33a4cc4684783c8445bb84c0b625b9bcdb6d23c78c57413c5c13e9dddbe1aed20347a841b6605930afcd194d4d6b314c51d351bab04360a3745ea2718cffe1223dddee1b89ad16d77da7bc84912de2b02eaaac95d44e7d50b5ecbef2cfd2b243c257c2c7ab23f7ee68301df98dcabdc8c98c6f0ad7d3b9a143231c63fc03c492b34400d6cee806fee679ccecc032a2de3baab7786622e12d0cfd7a7084992a3a88c4cded24e089b32e0cdeacba458fb51992e91d753d49e2f63e9f5e5225ee0fdd7594035a35f3d2acb9c466f849ef6ba04f7a6f12beaa1b76f49fb62aa31cdec6570937540d7610161b63950238a967142422b92fe1b8fe904a4272c80e31f31eeceebbcd433ee296a9965c825da360bf8266221f70e12a8bdbbd29c883327c5e3e2c167953a60b49c90760c0d0443f83023c8cc89fca22c57ad9c6b669b65b105464140e28870ae8064778461fe4d58f809853ba65d3b883cef480cae7bc01ecf205dc3803ee70516ce5230509cbe7f60a3185ff87454396b989415eef62e91b7373e3d3ad273d8c9e02d12292ba41a73c44b11bb96a1065a609aecf83fc6597c93635e3670330ef52033bc1ce6d32b05bee5715fc893f7bf45aa4fdaa8b66bc24bce25181cbfc708beace0a5b50d71c767e89c1e26b9505a8df228b0232b1d92bc735548213440a431152358da283cbadeac807679b53118eb99b748a9a811d889e51d7422a3ec8ff6fd060862838381f5d5882e512e2698c1c5db084bcef5914faa1cfa8b48a42c03e8d7d64b484b6181536cb00ee4e6d7e2794a48b4859ad00a135e76d6a5452a443b03f360c0c966ea98ff93a5ca609378a51fbe60f77540a7577d6f41e59d8a27eab98cebefc8377dc5cf3bf06431ffa6d26bdda9b94f1fe9cea59d8b20ec311470fc1afd3bbfa7598d97f7dbf2849bd2b2f32f0aad211c497b51dff5cc3a283850055056862c7c7b1eab79845facabd6ef6fe57423f2efe8b8806a588340af6943b4de669a4a86b5a51c13d1ea589d05ac03a6e70764087463ca6d3b922cf72aa318d28c2a14cf4c34420f490bf08365de1676242eb829a2e7c99a149729cddc4b439a224f96d8d0e115f9a35839c3ebde50fa0fa90d53dccc8e8eb0a857c260b0f3199293e9141b8d48211de227b1b896a14e2c778b2709d7a924819d6baf8ac700755b0f5cb613b11e061bd918aade1718fa36152f3f57ad4fd5c0bcf459dc0e21a12c5e3956ce87f0b1e164d328d2078238d2bbf3482e141a001b82a57e725289256739d8398c9283d130ca9eb90253b76ab33dc96965ab6d91ffef6e6014e19eadcc7b0d5df96a7e98390a24cbea69789065342c2cddefe7a69a414a2037cffb70fe21af66c7fb6d6afe2944b5380331c886559e792693c2b3d03b8a748fe6752f5c926085bc20981757afc527c98d2fac8be90d6e913140f3085d00fdf073daf1972d8ed97651245be34a1cdb8232c393198409d2b28aef9d046c6810f4c79473015c51f2daa4e9209f245547e3a634bcea6bf582c3042e27638d12772995d4ed378b4e9cf822f8fb3d3c3374dfd66ee30f4c3b73fc45e60d66b588d7ea945d0bd8db8847a1f5e00786678c93d78461dc1b9d4a6782809519ba9c9f98ef10313aa861568be980e081240f6308d9e6118af255103e719e8ae5f9e9fec3deff0fb706827a8de56848da2587eebc77c5856a66efda71052154ff5ff80a13f62da0ac67550063d76ab16f6bb88f4cf2a94e476e64685d257638c03e1a1ba35c30029d5a70fa05cc9c2ad85867b4ef8f28a3cd4e59b5f7fd8d1c270ed0bcc0572c440e532979f926734857dc48639c2ecdf61eee6879abd61cd90f581ada4edada659fbd7c6994ab44bea3024932522f25399e54303aa468a9dc808822e4685d0fabe7389666006d2a745c9f62c007803efe93b26d22c942949f866949585e322baa1034a1fca915e94193ce75beacaa5b7cf97d78f8d007435af7ce15e884fd6403b27fd0feecedcaaef2b7c1a6aa05a7f81a98776c1cd5e3f585d878884e7a36e619b90b639043d96bad908d5469c707c2748eedb9f94b9456c0ec15346e800fab2ad5bf57d513dd408a2ca0646e48f68ef843b27c61dd016a674adb64e0fe3e7e16189b72eead54cbbe08c72d5b37463bd6e1b60961936f9d79300915edbd2eb55da40cdc20068bd9a03d20885c4ed6e7d44256d1ab5b6bc87f3fcba85781c4f0461af7e3743704a57a55978328ee4bb3f2b798d871904ef63a17def48c949c0cadebc26cff135febdab3659eed772301b61facce981bd33601aff214f50c78e8e99fa84dd00c867c9a44920a9b4a96ffdb14cded7229cc33ead5dc5b89b99233525d811a361fae6043b162099205a5ea10c3ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6808216cc8e223ae81820887789754f236e3844ee8e232b886b482568003cacc60207f5e90bfe8e4c25556fa2034e2ad462c6fdc2f0ac698ad3b6f64cfba22a8c47cb3c252b6ea65db9499de3ea996e3260cd870481a7587c44eee160c46306f33b2b0efeb11a2a9198661c750533590f49939622a9dc4a1b88e8f38eb5b208cfd7617ba4b0bcb7d6065dd0cd957dc77a1e4116b485df01de94e56c413d041d969e1f4451c95b1d6f3a84c9aa0eb1b60863c3d511e85945bc0a42afac7c84e420e4a3a943e44d2613f920837b2f3ea4f4fb1f4e94873a10c44e9a8f860413c9d570adf0dacd3cb4a3e783e2122ccaa351fab1b7740f7953fe4859b10359f9a720675952378ff8d6e664c2127f3d721f7e5930096204f6dc1bfc899cebd53a5a5323991aeb41df80a6596dd5fe0e7430855d2ae816a57be839d1482d9653427de188232b3aacd4912fae0e19a8e8c53b7e4cf23b8cdf16b6c4864fb5a392453689e784e2c8dcacfb873622eeb1a75653e761618a580f378331c25727fec0bfc7a408c7301b0d652195f92969ad877b4a7f524f91c39dacb7f460d5ba2bd26803979185ae242c6fa88fe5a759e7fc2f3e6debe8bb79c480ef7100ab3a2c2b00e206ea2d92bd71db555148b38a1b1ff454026f978101b7aa08c7202b05a5e8894aa4c7464c576f07c818004d2d4d4a2180e2d2d9f5f0b2eafb0475bf48fc3e984c32a2b394db6c363e4354fbf016dd370b08da159d868314a36d068cc85f2e6924d9eb32ad9c7c79c0d34ba66aeff7861a5759d68704d5176c0858c8a2b4249ad60db1d0408050cf453d0eea8dc81027ab2deb77af4428654dbf00e69b2d3c31041f598f9ce005cd58898f2f802144ad3a7221f3a39f8720ded1cd2197ed8111c9c28461266e23620ee43e910627c675eb29bfe6c21c1106ba46085e850b04a67edb1ec28936763074167596e58678d01af9530bef2a08752eaf8ffa86bba0d985bd6d8419fa2c0f1000b46744e07cdb6c530cb50c4d1b9c1edbc31a250b8fa0e9a26fccd658b6cc4f49a6cac11c9912f94a5b587233b76d063b0d42e55f242b540107320c7db813aa6eb52d858e7c44fc1b96c1ae8e6d81f80a046c28c65b208b647e4e4f823e8512efd453470d89deb2041cc0f272d8bc2447bab20615cf914b04f4b0f4d06093278ac165e6bd914d374c8b97ed749dd64fc3bf76ba2787a6e5dce58d2cca32e690f9b1aff2565dc9124d225630523d0fbe758a56a5d3cb707374f58f0f84826fea096f84ae30e191074c6c094ebdc0e1a7f8dadd89c877509d44dc605c45e226651e5039fe7835eb82ddee47ba71be575f66ce4e93306ead9866d9833eaeb6a737cd2ee97f1d5962372ac01c499cde7b27c8e04a4cc2f973b760d098003c77abb29fc887930efa25fbd08bf14dfaee8d246e8985281ad69d96440bd2c2bd5e791319816cfead5ce72cd9b8d922fddaae2735c4e61207164c63bf49335e161beb24ca2293e3feb9f5720d6bada823adb3b8e33ef250ce374005ce3f072d9086d2f8649e2d73fe219943e8a8e01581068731cbc183977f3c9f11fa57549ed07cac7d2e5079a0cb73ee14d39fdc3dfc47f60e9d81fc8a55903adbf917feefe2c9fea0bfb3721f87c009cdd03cd625e0dd2d1b753442f1055ff2ec6793f1b4879fd136a6bcfc957e3555f12d94fefb43a0ee2994ed56b5a7edb6a8c7597b22df067b8673020ea3c0aa992f6178d583e5ae4134c33edf7f98fc4c93d3ff0460694c71f609c02a143352ce99bdb8dd7895fc19595b1d5196a436ede852c1d09d39970aaa62e6e74f5fdadbcf209dd091878a4a71c5e0543c1397b979575338cba020f97aab220126544c173bbfc995eeb53f85cff5505962845363e3adfdb9a9a1978e36d07b9baf9a484b753fc15155817b565c020653a9d9a1a8fd06f2e8f874e6de30d697f36fa7e0321f7cba9251c460ffcc525b2dd9fcdab24cf7dd5da59fd72a625c654947296d2a673418029b82a03115838143257ae43a42dac69adafd9d9190d0e2cf163cfcfe2907cd7efa70e97b561d4505ec5d91d5ca79a6eda18cfc63a8bb8c6984d4942691c7b526977327dfde6e9a609cf2a40bd6df84a2501ef38763f8d75d0ecb8c99071fa57fd2e646d0de48ec1cd090b45019293a67b8e143009c4e54e14757468cc683bbbc9b3c4e77f5110dc7411a778964f9f9e3c88f2bedcd4f0efbb00a342fd47ff23a801ddd14a8511e4130dfb7597369aea4d6551fe8d40120fbd8171f8f300ad52baefc7f619e7dae57d83032de3d42d021ca9461429746298c777d2487475f0dd04438aa7ad656f1c26dd56c37ae85b1a2171b6a5ddce8e5865234c8976a708243e9a9c88a6562e06e45550e3414ebe4d963e2729b7be594f6c64a961bd7fc446e9d6cc9000e64c40555fcc67b5c2d005039f8da8e5afb0cb7f6af73aeeef167760d48a01751f628c0f177d08fd0ea28ddfc00ee163f0609087787dd17b435ce7fa3c7c9a41fed208504ce9fbdbd8bdea741ec5e4339c2cee0d5838d6e5457b264bfaeeddb52ca195ce1c4813486b4e2dca5bca40ee6ed9011b556ddec0a08a9413fd87cb03a98022d9cbe034487c660e2b4d6f66cfa910703c0e6bcb64b517b655b2d5d2f3c121ad1430a7c4748029c1dc1c02ec01d37c2e242e0ae8b209aa1582d0ed65ce30dab532b3bc06ef75c7a2654c1b5a8fba9d43c126bf6f1a9aa82b393822a4c903a8005aec4d7c4b832926a99577fcd33e3b1bc75e44cd1eef7d20cc1ed7aecf125f4dc1799631935b55208eee7dcf155c936fbb8de6455a2626daa7b92a41b15f0b5517c55406b79d87f578c59e9349b941975f5931ee873749556fa65985b4fbc7b249cdb56412ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h954fb67a03c346dfe74a1a1652aa24e2bf771e28b226cfbbcb890d9c0ba3043eb29d57ffe649b9dc3c95c81f2b135420e4a2e140fa920e5a1b641ee6f2def9d1986527c8b11f0f92321fd593b9d4a28a1e4bb3fbab4a1278b8eae86cebaa0feab36b109a73e409e1ab15210f4845f90e753252e4fa14070ef6eed15b5d35ca4d39cca01e4d26a64d004d180412f29aaedb777783131c49873a61a9a442c911ac202954d4b102e59ba8f44777aa5b930396d63f646cae1ceb7b8c6f27ca7685093502ae8b35f735c833d11b39281d7b79275644380028115d2237a5b25ba6d4a2bdef1b27c86bb5612c7efd361f0e2c05dff91e9788b8c1551aa0e015a647b8a45638e27bac4bfb84bae4fc1e33236f5b0b4335504a6ddebb9845cb05e981ad82ea19644a593285d54b4ab983e1c261405a8dee01e23dea085a707f97878f319d414baf1043e8d10df579ae460f4532f8e358ed47aa6bad870325c0efd7026fc04d05ba3a57c3585dc748931b15cadc95538349ee53294c7b55dea71b92ad4ee51b38dc2a2d2daf7e85383b75ceb52f405e3a2c45a27520ef1da33b61588c3209194c27ab9ea1fa7d89a2336732a4f38f9667027dff674b048f6363f7c35bbe289fed2fe3284cdde46cd6fb5ef2dcce358f1f979345ee1ac14e120398e1ac22e9591960808325103f667665f0e9968edb868ecd8c89fe4617c673de209f413bcba04a427d6d74d4f6db1dd2da2579c4c255f6af4fab9fafb2611d8202e5d6043d7c1ad14287b76c2a84b0fac6a7c5a4b39647e34dca3cb8012a46658ea4cc31147b5fb3ab5df9e41941c9edf8ae6d905d5108ddea84d689663e3b9e2549613d5ac6fc094915ee8570c0b8909a7a4c3c4ba539650d8fd75334ae5b8c583491eef7576960768ecdefb9818a7f5be7080d66b9bd5b121b71ad49c66831b6a4a8dae4e50160dabe36184cee728dee85b4bf8ef7b1e855b38543f329869f54344aa3ce09585c752be0ad1e4b8ce918f06d83d7f70dc9e22dc1bb02efb6837d5314cea045a5d951418dec0303b41e70c8fccc1b625775b40a77eb7d9f27910a1869ad20d3d1a440c6abf62f5c80f55ecd890bcc396f095ea313dbf26e57b0715061c4849a6820cb6398e21286d9192598e8d509053a7897cc9d8fadf55ebc80a8e322da9674e7290cc22175738e8d998f984ab18e1af1d9a3cd2467cc3b35500ed6b6a2c41d47cbabdb81186b6589d9326483d2168a4b58924f49c5cd5e8ca023c4114ded36c358a15c26fd97fbf16b194d73e3bca8574394c3677552ef15737647272c3f89e0c6e394d6cc28659e2f59420fe52a2d8b41ea83b2767d661c6325bdbd2dc19f8ac34adfc58214bfea341a6481a4c9dfe7fe93eb35cded2a059f6d9fb7ee16972ca4b51c7a498ceeb2a60100458fb09f860c8dd3d344f4a6a88180cd3a5b7779e2e109fae49c41b01aa6a6b7572db7cbefc63daa9fdaeb489a4879cb089fd8736aa5aebc5e7ffb5601763d9a3520aad8a83cada7d93e62bf5b7c58506e5a0881b6b30ce1136aaa7c0dfa65a1a50647c9980bc7b2c29315d440fac796d8447274309608b86ab7160c9238201e2d6aeeb9c4eab8b8e273ec199bcc5134e76308e2a92ca66fef79cf61da010f75ff4b5dc6fdc2de80f7536fdaadf4e88ae6640e798cece3509372690537a220b110074dfeb9b44070eda0681d19e06e7653b379c33e0ff35e463273649b31b8b65d16afc80fa4403bd0f2515967950f7886096c0a7e4e286009ee80bcb1fd46b9c8db6671fd15cb9a8aefc18e6527a1ac4dfc4f04c4334b37fa0b0f0c11d74498810ee4287d78e07aa9aa82520c4df8e066c4cd44f0b24d5640295e855d472272ee0b6254cda1f56ddd30320d770e0aafc4372f60daa5bac771117adf8d001b3778a64f4e91e0d8943b1067c2402fdef3144f04092a881e0e31f2d6b3b1d9050702f5a31a793d7dafb055e333e0de2ece3d0f7f18de1a6a56d6a6bcf2eb6066dfdf14eab6941877eacca11fb0526af0fe5261be1651522394f465f294a02f6dbe32848990f32a5693aae70fb7d6143857ef4055ff4dd289322f627920d2d878f75b9b7cafcd9ad70b82036ea9b701c44f00c51cdce13b597bb9daae8fdf24e517166a212efdf119cde6acc2616f912400c359227c4a34472a5ddb2ae7eabfa871968b355ddd5d49e6945bce19d4ac31a56a77306b5dd3f1cb71637a524210898e99c83fc98785e1e41253f87e1ea51f14a7d32ed022673fedc1576b9061432f958217cf39c15ed7a123039e9321feac013dfba8c48eed08f6d7f235b27be1ce2db61386dc0c4b6665310e3a82c607e031d5ff7433c3868d5320a4660f157da1c01d73ea8dde72f9768eced7c807aa3d42764fa96a04423031890f6ea141c76feca0abcfee5820dfd88251f88ab130bd5cf026e99015cf28e823d8d932c6dcf6c3004b608a48c8462ae1d3b5e9eb99bafe9ad7ed1fb25f8f190ca6dcbbb3e3f00ff0ef5bac212095b6d65f6b44e307612e85ce53c81d68502b4a5b37adc55e531b806e63107c158cbd780cbf95440cd40bf520f670f929ebf29b5a9d0351e2a4827e46f1e10633135bcbc62539cd30d2392a56d6551fb81a50269c8edee59fdd92fb79dea3220ff2f3ad7860f47ab5b32b27398adcf6eabdd4794c0420546d304cfaf2c2b2ed3c2248825c612d63b0cb1e0cd1c5d4513413014da12a882fe16e6f850c615e73c59055505eb89a089bc39261a77f98e3f0d48e33e1c4d9a3272bc6f352a60e8fa48e3aa02ddba7a35e69e1f8239a26ee76d5d70ef29c9c1d9f13ff4b70b013cd379b6457cff78bb7e8c9a5e4836b6d08d48b3324e4ee7f6d0a4bd4da24700a6f13b218cf4af13a8097a03a7817;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h28f0038faefe1d1f4694ee36309490a9dd58a51d66ee68a471bee8942bbcf6aeb93af1a53286f113668b0084bf1453265babf2e42c39b8a0e4a1406f66b3547a339f131feb7c2b5e82c98e8d7ad8bdf0667363167f39dfa88e604a2a932ea1382ab2b5c264901c0cf73d045d288b19c257c9d5fc8a9da2bfe8f8c941a184cb3c92867e58e04930459dc1b9f970393d1326797ffbfc73e2a08fbcfea4c43b5269281b595e50e875b96f95f18a97a6b03f9e5bbba81e7bbcb1f376989fbd649b63f0b7bbbf19d7f07401d74c985bbe918bb588af5bca108e446cab488423cfdd4c7066e305e46c34a02925f50521b6f2c79f4bea7a1fbbc890bcf38edc9c5ab2426431486fb04fe8fedd36224c99d39dc4cb35c84f8f7aad112ea02b995810501b3b517b23107f606d2065467732e2e06b13c67813a7e290e946cdca8a5136d29d4524954feb334c734a148a54991b2d5e062fe12cb260fb3bad1a3a83f559a5f64cadbbbea93b1ff7fee65a480a10144fe0017eac3a1af0290f99a66abc12323b3c5f48ef65b32ce1b7c3db207a0996bb3ea2869eb9380604b74b2db1644b19b465c97a18d5bb2d72f7780cd2866d908181e4a893339c46511409e30d1978e6ab441f81dfb99c45328eb5914deb2fd5cb2c7369e6eaf602f6d2696800eef158ad94039ffc11a3895d6b8c326fef341ab3c196b8756dc24422b32d93c86db8c2faa595b42d528de3cd854b27eaae127d02ef266ce7ec6eacaeb9bdee21494913d73c7d2a1951aed1d9adeaf105f90a6aca352940e8b11694d1e63f43db047a89361d9f03bc9cbd1c47f4363b214a3cb511ba1f44cd44752c54a21017506e38e7c09506908b238ef112ea43522fa5ab0b40972684176b2fbd841153c2c405ae8e0caa141d869e92ba88deb4040784866418676fe5fb4c1effdb11656699c875abd530b9851d16b07c8b4004aa2726dc9834c135b1a99a2f7ce50ea5ea2c01e03b12b41e24aafe14992cd9a40ae5fd375ec43737983f03221d34b0440f25f58bb56290d75b57fb2e548a0fa010f3c87df9c7ba2cae4f3589eda5b023628e7a2c2a06a921f5032a9dfda304fcf687a942a801683332bff3be2ede79e7ac3d15baa7a948729886c6d3ce50e291f754b2dc390e3c90687ecbd7e9fa85ea4e7e318f5b7393ed0b68328ea7c3243ddbab9b01209588fbd57dca03a8aae389b9af8d765da39d21843c34a302346b3778c9a55353c96dfe27fa8cce2eb2773f20cc10065c6e3129aa4cc2080e37143ce7d64c1d8bc7e97a961ed215599b29c46668e40643e133bdf356ffeab28421d433f0835ca8b148b1d05604251df383cfab8776c1b53da739bd2f32cc78988f7633565e8caf0514b19c3f31082484a5becff586f136e4459bc4b82b8557020a306830a0758be0519e507c0465a168efe8e4760afc4bf08db49e092e4d81ca4d62b7deef3c056a1d70caf79493c0e60ffb1ed8b53cd6f08c6a86a2505d008601461cf14e269187a706f68c1bcf68f25d3f92dd7b720b6b52198ebb74e75121bd7c5c3505cdd272c7c525b548432fcaeb1fa130956d52aa383b0f9e450f6fc2ba7aa3ad2db2574b010648e02af3e2946c5cc7bd2ab6961ab3f68050ca6aa8c992d75459943bc76b01280c7bf93ca8917ce29de5994c9ba3c063f317e3a7e0c4eac070692e4a9cb2818bd66609b7e3c898abefe3c56cca8e38c4689065aafe1f264bc90aa0981d6395a12dc1acd6262e3fd04e573065d4a9a9fe807e0056b4a5a8346f0174a8e8f74b1d1871bf194e425ff75983cabc92daddcb563a5bedf0d395c8b521f8d5c4a30627ae1a829c2ef36fb0c5e789628fd5a79ffe4f95f3295618187bb15877d8c51e3a8185f7a5ab72ce892cfac45df5d6a0dc6c74e08f93de43364dee9795abdfabdae167ca7eae68723f018becd0ff5534330bb3aee5eabf4f83f9ffb5301ea6401c0512766a3db390629b255f531c20eb49f62d82bbe1bc5a839234e3c58a021cb96d424ab6c11042ad447ff6dcc889b3485dc18c6a4ac8f7b058236b95a3132a0f198a5e1ee1265f40e032e0b6baa67e99ff05041f693d81ec3440dd222dc5c8c1709575e05dc036f0b1bbcb6754ebf8703b29b009442f8effbe81ec65b65f7ff14cf8619627153f8367ed0d96e2b77a8b6abe7ebdda54062fab517c063ba1dabc73befbf97a8b0e918ca01543af8a109285dad156fe29c78df11e2cf3961a12b6f463cb2fe9f9b7b09b4bcb2df8df6e0ac2ee35d4afebe0856c792d6ea6cceb9359784c87e202f86ea8eea94943ff53c2ae48f2940dd6f70924b3a82173e7e2ff7d4c8948ed458e578bf110d65d29937a9e3bc7aab39919b35623d4fbd72383369ffa5aec201e01c2956b5b9275d279ccc6077cb27a469b19fb8bafd16235d3bf293cef6c5897f6034f0600c09d1b49a369788097d9247883349d33dbfc5f52792bca9d350114a4c30a81aed2749888b07941a466ff0b79262af629575f2061652f192e61627bbf1ed29b32cf4b524df3dfa32dd48b6bd84b535f7e16af46df16a737190020548174576494be78f41cada163c85d9588dbb1f376825ac299c5b77de263ed97d3b677c9c30e35dce0640c2db2c2ca8fa9af20cf090314a9b9bb70709c93f6bb9c0c1f75df46257968ac02dd421259c066e9e13f64e5ea1ebccbeb91de1fe0dd599c0b4fadd44a2b080d56a04d498bfb7cb1136bd6e7ca7fce4184675a934a5abf54ccc153c80056ad1abd1d9d582f6497acf3c02a290d5675fd3d22a8f5bc3f16fdaeb95dd41fc75395ba407dec20ffc0f2d36918895aaf87d1c955f3aef278afa7f51caf259936680f4e1a63ac6d1f9bd991ead7729c4804b1e7353c13021e406bcc746a0c2f13c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h77b87ef7cdb319ad0bb023359d0c4263dd70b578803d29e9090479884e44d28264552a81d3985df8a7146740e75d23014aaadc9b6799b1dfcbb6e895fca702935252978a797f0cd9376f5d5a8191c36a29bd7ecdacee5db5783b5fd0bf56615a4e35a594bbe008e425ab7614a95c61ff2a736150ea581c62e89550da6ebb404686959768ae7d1cc03a0cc563628b9525532495ea2f1aeadb52f1cbb2fee5f0534a7b2d1ed56fe1ad24d9244d5acde477a38031610e7d63ee699401e7a4854e81643865324ec0aaa0db5d6181654c8fb502658ca09034c52bf8ce132f4b481e052ea7ddfff69bf5bff8931b32be6cab757fed6d5c9b44225dabef3dbc62a22c0638f7df8ad5224b644ff66aafcc3ba48245b8efabb854430495bf013bd651cbc53089f8f75c385864cf699a428963bcd2c33758bf4ee1a93abb4440e74d0c22f357de34ac2d00eae1a04c859ada91cdd8222f527483d70b8aeff099425c4485412d1f3f2414b3c685726b6b0575d13f55337328d156b458c93a091c43d3e0ce5affc1c013e9e70335d41826371525d5f097104e152c5952c84c15911f974e649534171907ac37adbecf7d447cfd3bd48159faf5599662c5dffaa8975296b3d4c6745cb96f2cfb90c59f959e3fc12a6fbe8e344a5bd877b91999f35893ff72737c83c7932fe59c802dcc994747c9427b70a52156f27aa73be5ac6c64af97b6039113efc3e0e4b94858fbe6b377ad546b7a465721eab4c4b4b067b3c7ddcc00590544ef0fe3b44cdcaf2add23ee5c8d3d778e615c8b8d587cd636ccbca13b1c8f669ad7201f94abdb9e3d889fa1c3309a8f6eaa8ffb60d2c50d9c335b867901c309601553b7b49ee036bfd4fced7a82b2951603af9a903d28c6f936111cfd67bca1d6bdb3d1a4057776053ea44b46fc9b42477e834089fa18b0409f53de62a3bd59f4592550415e22b7170efb90c42d12ab7f394f9257f8f60b3b9579aae4db69aecf45bcad06ffac37510e097afb3973696c5fb22e99abfdfad08428fca4b539113014911268474a1015202abb51e9e23a6c9d1f0c6503b549b963b43680417cc23c2fb33e2cf2ed10a947aa73fc69443ed75b083e3028bed625aafc593b8850d4326d6da2b484168d7a441e2f1b62ae24c37b3a6d317ea4c10997d70a89ee4733c6c3a2a940158a7baf42ca03e347e490ec77b19c4121e72f1fb4bd0edaecbe48794dad84babb206953170463a472e7a472855e2733a175e830d91ae85441e53f0c85e5ad91fee41740089dbac89aa9d18ed90e4d6b72a95b119befe5102245bf9b9ac39574dfb925cd28289e7883d5f804d774ad2e7b02fe31342b37e5f8232e5aec2d7e041fcf644f50dcf44c98a427644cd73d409afe7372699cee38268f675b9118c50c9d63866d0ae8f26448b5777a41b43d9ba97d3ff19306c56229a82c91f6f25d17fa4a1e2f7dc49377e33d05c78a87f158b5f71a5e38d5de9a86c6ec125555e4165514540597f45d490e036f4a6428810895dd91e621945d7ee91fccbf2796ee548b0ccd7b908ba4c6e57908ac81f5089785923c7212e793d93e7bb855bf4d146892963173cfa6c0f78ebdb0adeeb9bc0a3962019fd9362050043b0850d8c43bfaa8625ee714928f2513944dde07daf91cccb3999c9f81e17babd4429ae903e13838595c243708b0cb801b072339533204765b9078b356a3028ca89534977df172ccf03ec4d05abac8f43f563e73de5b0fe7d8201de8d423858cc65c6282655b99f419ca31099f08714cbe8595f7ace4b560528bf287a534f79ae6696b6f6ae3abcdcae41a94ace029a41da55cd856f3cd9490cf620a47a62f90b186fcff94de054cb556600d148b32b2d255500a69d024263508d9aba1dfd952555977897d445f6b8e049a663ffb0080004e70fa98b4f0c8eddfeae6107a2e13309839b8876fe886a6c53351a41e947b66908f0f0d85296d136398e2dcef093775d3e6f287c67e234be2017e49fee7e5b5439284c5bc62aab6229f340ab1fa98121da5122df695d8ffd573f028cf4c25a59bba7e717c53295ff62efd16671d10fdbb275dc92e1f838eb40b7304f54c5a6d469e019bd3bb66d1a68bc30ae5c8af1a4a527ebc121292597f78e6f1fe63f8e27321f1900065c6a7ac63d740defeee6434ef1abf743bb74fdb22426bffcb7904abf8bec5709601056898264c3a2067dd46f5131b8027dbacb5c622a63a89adad00508d09d634edab798e89e49a7a76ffca26da977cb1fb0eaf58e5c7eb30fdfa82d6453532768ab1f6bef0a810f0f5c2609b99aec2e824835561fdf22dc6afbac34a38799008282985566636b099fcb099942fa4943eaf75e474ea58c3f9a9dc8366e335373518a8f4529514bafd4646769c817f4c437df030c9a15c154296e419fe37953e37eecddfa095e552c34c820ce56c2b26360c95567a4d3365a48991c48f5d7a9cd1604b5a56576c01e5703d49aa8045eb6b11c429e781072a22e9c73a3999f8c9ae1252f2274a6e3d8ccd449fe183233f1773bbcaadada3947157d489abed9c0af2eadf111ded83f8db4f3e3668c184fd16a876a38fa6d9e1eb28f30eb0d8ef2d7262eeb2f1c7b303d6388ce4390204e5e9fd7535cfab2cfe9bf2644d8c0df65eb0edd8e75602221f30fde229838ac1b53f6f98564446d99615d5e96394d2e0fd538de3c2b001d26ad054eccda2f364d70112f23f6b5c1b796ff7bac31e4dd0215eb191f143856d58cd2ba88d326b795ed2de235867c7bc7ffb1f07153953f290c7c039614974d61c236cc335ad0d86cf9141d533b343c3b0cb8ddfafad0660af161be025d64edef9801fa0f165491f121e484498a62553d99afa0277061107d983f319a2e6c9ba023051cd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf65fdda04434c976d671b23079735b0a0aebf52136567304387944e184d874a9d5feab4d89e860d54cb90349060acb1030d76b265b07f61f43b40cd783431c43c5f3feebdb70076a4f45f21d571231fb10e54ae523242c513090a0ddac9776769b4cd3dd9fd1fd56e78419694ccb4027457e617aa3e615ebeffd76d5009b88d6c96e3d06e72c3497eab494f9d6263333c562001ede988377647f0abd5220a1093979c7c9632859e6a4d15af701bfe546d4fe84a6925909fca3f74c503b5cc5fa35c128e2f0f341c6d2111cab0ba4921316980df2e4510bb77b4ae18fde8465c545eaf0ea8e0f04ab6105af3112d907bf0c6c753708643160fdccd6a9c0b2632701f6f80fb0c6b487088cc2fcb88b5fbbd35adc4cdedaf84786ea386546655b270dad618de25d802ac48eef8bd7a2a6413f0ea70875a82e00b9a49c86008e8045fe8a914bd16779444a7fca8894c1ea840ae506fd0ff30512f6fc1a233908536bc803bcc84bb156c1f055fe4eae3f53620f3a80ffd4e356aa905795c7cb7e45d31f4b416e055a3223b92cff63ba3434e54d9940d6f765ec29e3412081a697527c074535bf749a7fef3db1e6fd2a34364448aeeafd68b4d81bb45d72996eb1a8743daf3b3f314f314d63793a21eebd6c778956b3e41bddfb9dad467c77905c5d571035848161a96d4a57d24e5272b9488d6fe75694f6e56089ae8dd77c4cda968d4796f3fca29996809130a1a248b996339ee10f512585a4f5b2eba493ea8825149a56950be6a26084c677361e96caaf0c69b9ef5953190dc700273aa4dd0b9bd92d0da3bb4728ce69b6201155402d06cf4a4493ea8eb51677aaad2aa74902a967e85de5e57b45b8d3fb2e48a4cf35d012fbe282016b32c19db7f89df31e25a2658294ef1d44b7eb7d58af0055eeb57e7dd1c44e1d68cd87170931f00f6327a137b39b7a2bde3c122da3f6b387b208cd97d22e9de628bba16504002be0c341bc4db2529fb3f563d5d79847a352d0ecc02ea498330d166f0d7af51053c0e03246b2e9a55477b84c9864c9020417abb249d65a82f6fdf5dae136cc8ffa142dc588802bdff79ef23eff24bfe1e20825486cb1ed87d6e387e8b73710e0614a1ce8a2257b379ad8e064fc654a2078f4f8694cbd50edb6843a1327d2f83386db1b03c1d532cf87993b120e3b2d5e1d8f8b7eeeea4d83e591a70457d9af403331da847fee86d414ac94051aef425548823c7fc5b3be80e9bc8f7e69a6792661a02fbf28f213b4e53c81195b68153134e992479a2950d3c70daeb274e3d84629111228119f880f98e4d0bfc4de2b281c641d5fbc5b697e295cdba86e53c32b6492124d36ea7d33c75b17ee9bb5b996ef950cdb6d55d69947aad374956966ca93c65e9c4917d814be1c3e76ba6e011d09d87f9b2cd9bd89c49087adff9cf30d6a9b4aa045ce0c1942067f280b588778d49b5bfc146a42152a1d75afcac3fddcf5b13738f047433a0a4d63b330acf44a5cbaf820067b1442e69f60addf751090d86cc00c47425a70f11e40656ba42d560d1e3f285f2bac488a7ea9d800e3846215981c923711dc282b7787d9467f58c529cae414da03ca58f418c1b63cdfaeaa90b47a529d43332e8f66a319a99744f8acea97aae86b2845e92a551c2d6a73a56b55b2133b7e5dd532699dded521052c45690785d3e8a9b8429258afef62006d387b88dd430a4c8620f96bba44a05403754f83bae95462d1d74693d9008984f1a8702f6ae6568851d0ea958667db5fafaf5d4bd2b355b22d6097b8bd7ef4f36ad823843f6db27ad177a12c8c6264dbf87bbf1acf7c6d773589db5e0eb07363d820c402f6774331c94129471f488bdfc6d35ac051d62d4a9409eb0154f91a60e718cfb56e3f8889e0bdb2c2d9452c6292cab4e08f78c88daf4174e49ae7a4685e75056e1ad49abadc5ec211ea58baa2164710a33a98577a6b823e1fec75ffe1aa7e605c94889f120456af40a7331a267c6befe5d85b94bb351779ce68a6aa66d8465888726d457ac7229d1489ddfaa510378978ab133e47b6654a21d9b1044741afa261a5da03496a7bb8d312f0f5ce5b829366f35e11324c017c56e20a1d204feb282eb245ad364ed3c7c934c0f8d40907ec201d2ca75f809be01a6e72f6f70deedb801f8adeb10ed91b1f861535c480b1b8810af5d474b994bdf42fbf7586d99060a3884c6de29d524fd1b075173d03230919ba467238b51f69ef1ddef7baf996c2097d496adabb1deeacd43c43eeb06435c8912ecd415830e88a74e417836504a2cd8dbd124573ef55049f5f080bae5b70af7ab3f6ad4be9f0d7627be5f459369f3c6f6b8bd86c1bddfbceab92f8d3b6584f3581a96c72bb36fd4c2265e1d408f2ec00b097d1402376e1015ff58eb5366573f86678b22cb50e925110c73dcf43a06b40adf562ba6dae892a2891ee9a7f440e6fe63dca2f55e1ab72e00cfd9f6f5baa74583e5dd414d3ad1c2be1b9231dd3429215c48308ff7faf77af15d1fa023b418a821a2b0a998ce6a34aef5a3e7472bd87fecd434a3fad3972b335db3399faa77272e7436a8d5fa361effc685ed144f4f3818d22e139d1737bfa3875ed285991d7b130baadbc0e175211fe9cda33465d5d97d6d321737a79d7c0ff0ae92bfa8d5c839608245651d0c56e44231b2302d71a0d746eea7dec7765aea3ad65ba33c559f48cda44a3124319dfe134f504c2c0f1c092183e07c3942b098811bad6b8e18e8a4a045383479b9269c9cb16a377d3d9ee3c79a8b1a098ce5396260c271759bf34d717b5a42e7c760856f6192671a091d8ae7c83b30866c3265778ae0d4a0f8a7f5c757099ba393a965471fcf1849a11116855c0f85a7d6eac96f70516ed6c206ab2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h98188abf5964c5be6bdbc0d358aacbd7fe211abda5ce632fa7be3050c764ad6373e27742ade4f4c98600e4e488fb291a36a832f5d7754a25092fef15c358a7a449692147d27b1b3a4d15d887cea362f03b57c69c5e0b4e1d5a54f181c405d720c6a9980fa34c29866b95864ddf082b9590d081c3280de5e2b54ae80ab9b2ade7b513a504d3ec6d961a8407e5bdda496bde74440516eea1f19ddd3e00729a62084e663377d991f4563e58a58c61a7524b8304bee49cfa36fa0ec917c0605cc0453599e85fe75892d58f3efac1347def8bd265d18fbb89fdb8f4cbdf9f8a1ba0408d31681627f079194435bb82adf5bdf0629b6f78009c8636a9f15f4f48045016f4d4eda632273bbd63fd3e4e5845407ba941995b3e04ee51fae42a86e1c6c95fbd285f0125f4badc13461b900ecd630e141210073b46578414fa276e9360a60eb1d3b347972b1cf4cef6ed61d1c565b60951d45cbed37c8e6d1a0b5097624dc8ede043801b09530a5a2a65f3dc7c4afe35c853b0b477543a47132c7a4cf64c996b35761aa4fea6a60053a3d328da352bcf9bc987370c450d1737e304ed660cd635b3c8ac5683f9678fe3cca911bc305df42aee16db562d872ab0a9645c52cb523ce0924cd13dc6abb49f0f74ec4744e9aa222f8fa3c6f6c656fc077e25c82ebb5bdb15d4ce0ca4fa191e96ae085dfea9e5c89ca940a94b2bc6b68297ce78ee434425b708b7ae5239ba22b8b4e8d21c653833658c8fc063401aceb875e7af92d6c5901f0770fa496b19c1d68371d5920eed50327bb6b591d032abdc0a25a1009fb88e19b298e0aaa8f42d5175d745e436fdc3c67eda9eac1d52eb710635272d0cb19b8088f586966e4aafb5c35f0127708f9eee9d495bd1cd3baf99d8fb205b769f632620702c9f81567070881634ca206c6b8c0581455d49788cedcae184ab4e44d97484c1b6a5cd0e1cb49e3b7e22531aea2576061c1aa4ff3babc51312a4e5c9f1ed08887cdf44601d02d6c9197b8b6de9cf21f2599c7f110544a8b891911e91366e7fa87f31fcf4ba30263da7204d5457185a57ae82c0c2e65cc963920e8d1aa0441d80660433177c5f01d1cffb1b78d569db1c2cec283a98ea2fa0d2f8885bb35bbb435e0cccb7199ed0802443f118c48017f06ae0a0591b051b955b6e96bdb18c3c7744e770206dfc60bec70e0502fcdad4d87dfa9e647604f892f4750aee5553a11a2ce39e06ecb0918b6d2c5344312e4cfa313f6d85413d323be89505cc3557baaf3881acf0722d7d0dc2b4c761b7b32fb68178afbbc22802326f705846235171fe0ef7ede9f800f17e07c36181d89366a09cd94c4637e839123daaca42f638ddafc8cc13da34436723e705026d45efa18eed687caa1b7804f6011bf7c5f55ae5d7065ee1ecd86edd35f99dc627776ad38a6b827da255841dac9c98981f2055bf07648693712c7300163ccc905b3048655b1cffff478b85a7efd4960a9556ee34048b2428bf236a421d39a6a694e3d35948a7fe03bbfa621416cd4c28993d93a4f5b66b232c63caa2335490aae0c4ed8def7ae90c3c07d1f432f77f141960d6a35932d0d78c562641215e5fa5e1bce9f5504104b9450c28d64c8675c29b2a6058655d4192fea3d8dae5e6c49ad180c05a8225366b7a2fbd66d89a374c1d5fb9cdeefa0a54a653448a8e8b45abdf0a96bcc25c4810479617a34ad1fc15134320981089b655a437d5fba57b3f36525a65598224ade88c0a5bd0d530acf5e290d4e633138a93e300dfbffb53fd5c28086885da9377de1eecd02dfa509d21eca527d41fbf338748af59edbc7c5f2a654dc5492cd625e7e8b6188fd788f0efca83e47d33620d291d65de93af31fa3c068ab802b09dbdba6ec5c9f46bd0956a2a7508d0a2cded75eef42bce9b5e095e90e8f7595e59116dac0775a7589bc2b3dfe4cfdb9d39b0534c5a6ab8057a4dfcdb9a1b1cf545bc42a59e31e1d9ba642b77adda6c4fd9d98d990d0ecbbe2437a46a94c00bd55c6aa0bece574537ebafcb36f817b62c930de4a308be2529527c0d1b9250e976fdad0077b540e6a22e35e29e3abae50f295a13fe18e48adb1cbe7a45e9efd9c031bcf244323b6b1e56f5790cda48cfaadff64797e75321afa906ae78975ee7c4474eb1d5cd54aa4c1b86a83215efe7b6c05fcdb70bfe53f38e96765bbd0bcc0300769589391d7d2210ac7e14e94812251626537c479c344c504ce63ff57a4e2c1f8f60bd3d250e95eec58acd6f187b0956d49923378235ced42187e50f057a890330078e360be1d21d1e7fa0817b00694bc7e61d048d2db85e67b2f41d04d01eca087d8e22b54e8391073a38db8510541d7009fa67a4140c9cc5a26e0de2777f14fdbe465e3511bd8a0c223f3fecb1882188b13a6b71d9e1e8e08b94fffbab647c6ef6f0948749ebcc4d0e419401066b857ffb8779d6b3e90722644c7b97e8cc95c3dd1ec26367fa956767bc6abe3d9a81f4ceb0f0873a02f7781029b2a90608d9b438ebee1c9c4b9d827b133dda7275df887b22b64b7cb5bbf42284f443bfa44fd25e57c27c0a0442c75a4e3efe355f4750a505e832781eda3446032b3f63f19b039391c733b800f314efea8d97c48206eb2eee4d789d25fb029b32dcc80b836f75a650ff31d447f01d7dac61692e8db680351f8ef245f265d43f472efc4ecc30f1f171b354b895438d31e92e8c6f887fbd048d1610c32bee9b356dce658c5aece0c8518e466d84a4c642a54bffb5b3cee781a106c32c6f954dd9c65813dcaabb150eb6bef85dd301b71f3b068df26f87c4421d734db1508f0c449ea865810250ef821fbd72b32b0f6e7af7a53539c98ab9d70605ae9738517384838fd5ff7c3a972e8e5dfd51ffa74817;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb520343680848485f808a2925d9114475c1fa7a5545851c5aa2dd820e1cc786886f7306e3b9516a5f996ad46ee9204b089e9e27104e8a4e0b9bfa787bb570c1c4e18784e2014f10f47d18ff41228c0d0d44b52d451683e0d35754191e825aef0c1d81ac80cfec1775291dd493ceaf681c019d77583228c1f3d6e33c9d90480eb5416ca6e1112f9e177989d580b49b43a7d52e0cf83701f7151af79dcc67bf4ffc1b65eb89136a63ef3a08f99fc3eb3fa4f1c55f0792d64fa1b70f4ada328176f5311b10b7dd3ab47f7e4bf8998951c665717e5abf68c00b1785e491c50838f3892d62aa2839a45fda3cd54187115900c11d1cf28ac01d5f3306bd18ed6d5b58e6e2eb5ac92434be210515ecd4b500ef791264c39bc998c6e62c53c3e02afcdd9c9eac2cc9f4d1e4cdbc25e21d0d999425dca0e57e026a61da653019d2d607a5d288637ea619f978fe1c9d6f083ad99d8bff8a11d1c5123da7866a294bdedfa59cf8f38904af6941d286e13dafb43a2b25db16b66d59aeaf20b162e43c7dc6b5b75323f8de5185209b6840181e29dd76687339ae55745a09830a3f6ce20c45148bcb3de1f4d9281b47d41ad1b3507259775c50a56fd75bac82fb6d3c6b444371a9118ca999d5f3244988fadb0858a6050ea2a99fddddcb1d918cf16653c8a8c4d83005abce727a31e2e452fec34def46a4081d79f6d480afc777103130738fa48b889f20dbd0e07c8f44111157863ccafdbd68527f4efad3018332c5fc49d8b2f273621c0b34785445cb573dfdb2ceba1b6bcf03e8629ffbc368b64d5f45cfeb03ff1f76cb01a723f9df065aaf9d92c676d639529dd5464c682b0cddc66b6053fbc45e570d507968162513591284eed8d6cf1edae7c8b8af1015ba95c48b73c4272f41492694d1cb7ab32eaeb605ff441c3e00324f073f42eb6df1bab7a1363e59686fb46d336c49de11e2460425b18798b83bb4c4358f72ebd468c47c1292b7579e432b983fc65cf1ecc5ebab1ea96e3ca08328590f22eb649e032e37baba36e92cce0a6adb307ebd694ca42fe8e230f311422a8331b82910e4bcd16c5bc32b4069d3f74844f64e20ebed638b8a505d315c972591a3481fe1d9b1008f399d72162b340e28bbd66ce62feeefed3d2ecf0e9ab1efc4b1240356fe5620690f30ec4e508b06f61ce2a0056727afe06e29ee34d1bec106c9ec7b2e184692e030f131b2cfad40da3a86b74d86a3e2fc1a71266d319dd6532c1bac8da8387bd8d8dbe9174e0f3b488eaae04e519b90fd3c72e77df7b181dfeee52da4a04303bc5bf5e0f4df02ff8546070817a5fe3d034d532c04741397910561d8bf7670768461f1b0639177e4fdb2f724a01c9edf6a2f19c3fee9f6e523c8afe2ecd17397e1e6ea9f96ba2b0170c9851d42f07c44497218ec01c067ff229ddab9637090ab69c8bb073d3a9d9728cf586f0edec786e378a6de0dc17dc35f1b7983282a8e1532a7248ba1e3059a0f1e98faed70410387eff317ec10aaa09ec12077f0a330ff79531d2b40912ef18f3e899ddd437f36e6666aacfb4dde54eee4a7c349724cab3fd12a8ac9bbb14bf6d80db7b0da0aa6d4d6f61a9323e7c6c8d4fd75990922238d4d44dee7e9553cdbbbc0a6e9ffb8fe115d25a9681b3b62bf65ddae7245d173a39e7e69e7f4667cc1e295c45cb396ae8a2e16eedf007b227ef82cab0a0bbdfb1e3277438b8728750620f8da7cbad78f55e7e52dd1bfe11022f268f5334632f0d032d9b966eca8fcd5a84b8f4958f8ecd7f53aadb73c5740b792f062c7be823c014128e03b0d68810e52dd3472c805cd27e829c3e2e2b4fcc28a79a15ac8fb7f4e71b3c6250d7da56f17f8c0c714e1b2cf7fb0c0bfdd3955b76b05855674493cbbd91c38966c59b0959f4f092bebebbcddb3f1fa033d71406858749fbfcbc46165f6b7cdbfb21e0da12fa015b8c566330c1c2491dcd0013a3974c9abe075b0a08be6a73213775cfd634ecb921ad18a8f73a387ce639ae01d522a0409bfc9699add6e1d1238d6a203e9adc6f79c9557372bb74def93cef94e55464c4b707b777081de9021578e7322e03b4f40cb862be8f496f532ea6ba44d134215900b618b7cc16832f34fcfa782eeedbd3f475192015c7e861e5fd0519cb649828b5d96378e0072ea9d90a69b50955bc569627cce61ad3ce86469ae1603cd9b06db495b63279bcc72a0cbb50d080bf8a396f1098092d95fa5ff33fec29866b86e3a9395c890b38f582d07b439f5b74e754fc457bc0b3e9e78f7f9c1c850ef099b24ae61e968c631df8820f344716ad74bd6152e974ec9f3761788aea2f05fbc6d939e4ea7ba9e3eea5f6adcc6f6b53bca6b63353584bca71f8f4a91ad2acf3f807e5ced6cf7e7297c65677c2050a0bfb4ac051600e85ab0cfe7f75acb864689585a68c7aa3d261cdc96523841e4466e529013138d1c060e7ee4fb70b6e84ff695f35a5f2c8e0c578f025cd78bcb8e1f18afe59148e95377d49b36b412f1815fe66a773df81981d78bfe096b61cbcc35bf5e2f152204d71af44106372ed1a309bc8a034c80e5035b2916c9ca31ef03a343c6ddcfecb95b18c2f663ae1c2509f3b322c4ee682c0a63f8db7073a66d6317271433e23342940511066c6d9ed9c6a0564887f74cb7762a685039489de631665e3204ce44dbb3d07bc0bbc962e854400bf329ab086bab7166b7445accdd5ba6f9f98c5ded1acf3541746be80471c93e45a11d10210d6427cf2df3ffe16d89782198a0bf5de2d5125133e530bc96afaa6aec4719e8c34ed9fd1d4cd83e27c4e71508ac9a37b196a0cb436928d62bbe53b6a08214a426703592e7a5f35b0c9ecd78ad058bab98ec257db2e52a1380a2f1a6cbaf317b0986658c3c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5f1c6f942e06c95e29a8b724f64b07f3f99d9eb55be0102e79d5ad2178d7ee1ea0fbb3f0724b4bf69655dd4cbd6e33f9bbed9896608149086fc3b5f5089d3541b990fc158b4df09454d33caa5771a85d30075aaac878a1d3d41f979a9aa6a74a708125520ff75fd11d9780015e4ad9f4e7550bc4594333ca6be8f1193f6134fe7d8c7673122d4c383b75fcd4774e7a9a189c6f78b19ff43e51974c66c0d8328fbc3dc672f17c7f349d7badbdc8d61d9c61a6885c0c4150194208867bc589a6476603705aeec43ee3498e292c88c7e54b5c49839585be20606ff583e6580270cc596c046b5560ead587ed138004ec5a13ce3649178bd2e034bfba562dec41d10289495261c95d445c921ed9ffa42b2705a596a3d7b318d1acaf68f46fb6132bae2fe3fcb16a4f5c5b793ad5d718276414d8f13fa8773b54585dcdf2d9e85c5c7fea24bbf0d9045566a8901d099493609e154144178b046cf414440b0f9560cdafa50cfe3c39f95ba8e7057592106f6267dd52dbd9d466a9c334f2a114d28cfc123eb365621f28190f19d5dd3081d19b7b898fb3dfdbcc7e68de0bd868b4233e46379902b8ea48982e4314970fcbafecc602b50d619dfaa2bedaa8c1278001bad37160331e106e1e6c6d7693b703344e2664a24f942ef982a71aaed68a8e5c9b9ed955d40b5393701504c9de89fc5039cb3ae21cd831dba0e93b6950f1f8649de387659d8f71d3686b46072d8606dbb595343de95f159f20ab4ea26f334158bd15eac2272c7301a1f0ca8a57748f5d6335b9e15c8bbfd9d4326ff0782753108401cd1f7172aaac4d632bfb1c19040445c33b421e872190c3a68ff867240ebbfd184e4e2347c10aee3f1910848524d401caf5c3bcbc46fd131f0c6cbdefa0901c7e01787e28beff5f1439f32eb1606c7577c8ba5665ecb58d17add8658af4baf2d894730a0687f720bb5d6fcc6c3c01ce8a56ac5bc459e8eb7ea73e30e78c43ca0c485c2c5c2bd272690fec61c78a12eb276207d16cc806ffec33fcf2487af384ec688bbdb977e14376e5165ef834f75a295a0ad87bd9eb748fb40e0a08c39ddcbb1a221575bc16bbeb403974da942a2af54c7c746c0255c8853d800927c599e444deccd2b6662f7e159911d659fd6e38ba14f623ce226252bf970119a1cc045d78450dc06b9f77cde493cca35ece2bf25e8c7636ffa3de8e4882775037e7f0407c03ae78b36f0782b84b1e2e3b77214f299c449c2786c5331589fd08a9eecb93287ae03b715e09b03bff4562cc5d252bcfd9e10c2bdfec3d538b30f6e4bf83db72ebf9503114aa4f4c16609f6449cec15fbb6094827f5d1279a8ad3b6b78d20727e3deb5782ede0bad994870630c434fc6e19af6625ef4f9f46c8b676fa9a31ec85c0bb51d9c20a8fc3021652eff46a74ada0462e0c79783c7ed6664b5f6fc541ef138faa8a83f3e2d539d1813d106942a67cdac1a471ceecf7fcd7be68c015eb4df6742c8800f56316191a29d36cc1b3f12d16d1673ec9e21e9526154130ab67ca4a36c6eac3c623fc500384c984cdbcc494cb9f69d38e49ff150415c65ae11767166fefd2b30fe39e5cdb726e21161f39de31e053ae29f3938c339303c625251261c56f04ae0ceadbee9ca541290b5d54d9e8533d4493b437c56aacbf5652e662163ac3e32a22797800fd6a5fae008352e01f28ab571a18f69823ab7e977c0b31fcf6933ecfb05ebbc2ebb88041d9375c7b607e7432f7906139f6aac75c3733ca2288fc2b1e8f1310b99002104000448ddf913c2b218083bba2e17ee6d85bc8c3a34ff55664dd739b9b1d3e57a36957c697078accf62c54b20e296ce056cffd6dad4900af1e6acf1ba648394478592916fec91e28e18725c41815f4bc388c13d4f6ff395e4e1a7ed30da84900f034401eef693b3f5923681d1a6311de7814a717f76ef4ed2f123bcaf3e087fdebc3d65ff4961dad79d0057d7c390ead9b17e2649967c40d6e3f7876b270535b27801d0bee90bec845ca595acf43d1eb54d8b88b038060a14588e3722ac9c6e0d97b724e8dcc8b6d10bcc623be28eaa346e0c23e6fc82b61d92914fdc61fa24389e92a874c210592a218ea398e83417acb17fb1208df360e7d211ff4a0ade92a00e246ba87d09b838847fbffa359a98ae65e4e9bf20aa48a41bea17904732b6e8b7be26e9f418633152da7ee1e96e4507de6b0494f44a6506074248b376a9785000c56e3e71e867acb98838e33a68c0f94745fceebb4353bdd116ed3c8bc9f2879819a350c64401952b2c0bc8ece9980b92ef8f05924eb1434bc1cf9876c6bcd729e14e79c1ad4dedad90d1a90f5439d6528bb74696c53af47901cf84e0e1cce5aa9498fbacc5742cab6a58828cacce866a332f7c257071e24dbd23be4949349e6076d70c8edc53b381ab025213710f63ea825e6632f8ec851a4093fa48e51804b78218f48df359541ee9f89911c6df8ac5b56391dd73ce8fb3e0e5b10e90dd75b16bd696ac8249d70803869c6299105e3ed2c6a30a2a9517780696f8a7e80fda2452cdf84da3d54c3ba34f9d19a43e0d566bb757a8f235d835729c32a668f6eca1013bae02616f84118538d68d6874bec29cb885a0bc7998453fe07ed0f518f21b942fe1151ac2469a865236c6caa38112e3d8d0f8fb43c7ab27f869bd2616804724035693b994f08ad8ff37dc15425de78a4b2d8b1d1b22593a5c288f62d5f75a59029b9ac9b30ba6689f95c4e72a81a60d42482630fb1a5f29fd4109c7f2b29ed15a14f9c346c1ef38434653e3b98f0ba00957559ac0f13f01c35f22f97f262b12d959d2da8454ef56779ca6a74a2bb88effc3cd72716809e548215059a5de309ba2c1c62b5a3d52eb2be87d696e73f543c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he9d77de4424f688b08327945506c7774ed22d933a7355f3b96e359345bda7515f319cca4c3a6d0b4072fe49b7251807987bac1ea01cfd13d09a0dadfd46dc804f8bf7fee5022964302dc2bca9e348514af03a41f12b096c694a88079070b1c42651894a72da05bd4c3badffc6e2d3709adf11190eb5437508fb0b713c283a619291bda7036be11d4676364039dcf53f91b713c284eb2127a46105bce6518c4edabd6cb308e9d49795e4469dcf41ae20a707af0960fc9d57642ee477f9a965a51e6e417035f946c8686f498cdf6699fe5c85e679e73689d7969d1a39c945c849166a28f7fe5d2fc05b1b973a5b72bdbf3cea98ac145a80f8375fa5cd5f3149a55986cdb090a1688926c6f9fd354e98f1ac5de6d2560c4f27656993bc1ebb4fe8026c91dbb8d31dd4ee2b46d3249891fcd883338c4cdd8500c6e312036a2899707b5810ee85b68a84fb1d15df13cd665708888af09b6b81a024d8f33096aec64a4619a4bc09b5ef7f6c20cccbd639ec4999baf51e3c562d8a0c1cd9515f1a5c0bfc56cffd49e3ffd1dad0e1aaaf35ff1bd2f909f508b5b34a199a46bfc1290b60e9d8934b453389a746d2d9d5b41ff96b696fa600f41f536700611430b67c032556be55b66ecf0ca4ca6afce0f0260457ece18113bc5aa391b6080e6a021f34f23dd0a9d84d7f27dc13afd738c0dcf87792ae4fbeb2ab2b26d730eca134d071a2091dec32cafc7511814db8ee5fc9c8de5024ac14f36941523f48d91b40a85dd76e3cc98e22bad4feeae773e6246211e13d53b39e2d954e434642b8e91efa37b4358d2527d7d60feb14d10121108f1a2377ae7389ee58ae3e686571d3d2142da3b66398fe5ebe419dcb338ec5909e48ffd6942afd3115b1b67a3a11ddd7a6d2c27f20a506277836f9b50c9d98c1feca176f10ee3788ddf23a3bf61d7ab72c59f30b4773c4c00d87e947c401cc87dbee2fa8de424a321059ed99615ece799810f18df4a87ec6bfcdb43aaa1db03e40ab55c06d226aa82bf4fdce08e6144ae61e98b59e13c553c3f9359faab074ff84c711bf6978877e67c0688ea98ae444bf39f1afbd0ae607aa237979ab074d85ad62a809a58a517d8ffba4cc13b76a1b917ab6af15fb087a871f0dabac93e6a512f3904f4559113cdad3020655997fbe0772b797a5f00e43b952f64d85010a6a36050307c288a3156137a16277413f963c66254756a96753e73ca553c4b328fde76cab4f08d84ee083de54433255d50558253ff05b42665e36211beb3f2ae92c5249af735cce210a647baf8374a803b89ad89d121acb997ffaad0fe17816f0162b9ce9d47c88bfb7338cff057cc402c0670126fc18ba1be860ef7a5406bba6e4995efd334070e31ee96e3a854acaae74081d28e814fe8be819b29ad976b2e6e9889eaa26e93b5d66c5179b37826666588864e13ef29d8a6506ea20d4f7f96bba57588eff8bc43e532cdfa9f0834767dc33ac6a0b9ffc52b3d1c99223fdcd5944d722073f097958319f6c66bacb64f190745bc9e7a667b0c1168ee81709dd070b028dfa9f7402e93d88e777db4b5c34ccc652b12d7771268b161ae37ace57f51aafd6937cf97b64fcc49e44d3b91da8d4596eca884b3dbf51aa3a3df44af49cf0eee424939e3187955f979e56b006aa2c63da140ba1300e8cc1d7def829faff6f5d925cfb4ea4a7e0938b6990fc8929372bd33a28e631587681a281cb45011638cdb21faa3ee022487eba27eebacff938c7b7bc93e642c78b3e9b7b0c1933ddd92342b8f41475629e63e15e32adf820191039e4ea104897226535bd607249c0fa56868dbc9b03c1dc35079969f70246408924d5b8ff7495d92a8f668642f0e72c35de3aba664579497ade3ca9a2ad1ab05cf5b551d415d3d356c868f9679fee090808ff7ad72953f9066ae99c939a8e43e96b9a52385edf1d210def1f7c129cd778b8880775cec02742e87a6cbc4ec292dc4e41e14e5ba426e2980c2a0942cd9b60a8a82eece9f03e38802c585c7b1029fc8e471a0a59c88daa652fe5b6254109c25bfcdd5a79481a4f16e353dfe4e949352966e4a4dc51ddcb0eadc43991f92c9e24ee5347fce4b2b69c7c1f75fc1262b920fd9f06fe77fea900394345c76e6cb9089a22d2b32b44b97d3f6c3406c8bf80a385dc183791be3bf3b80b4f3380d8ce4c33f022c9d04d4ff5f4f2b0996b54786b872d36495151f05ea8038176d07790404b3f90064446203092de8dd16cc01ac57515ee08f2a382c66b1d0becf2a6b64023470dd96a8dac44877a2745e78b02cbd4e134dc544746d34cf8943fea7d7407a3b1e80ab34b80e5c4b4e90154ec87b3bc23e77e779eff1aef964af793ba418d64c9492fd164af362b4745ecaee420893d8afe9f23bf7d95d2a4f9b278428a561e3407bb7923fce67a20c0119dc6f165df8377f9bb50e1779b08360e7954b281309e1e00a7ce19b1fd2034787909acb4abe559d2d85e2be434ce9d7608cc53399e7a1ff5238d8507877c21ab5cfe1ec69c64748c1121afe6c3d924f449416bec49f1accf46dd7afe029a3a1c3b4a91143bc2646f5c0d550f0b0485bb792f92e6273cf8294a6c4e8ddf8ddab51585bbbfab4d36ee581f122c5658fb81879110d5d7026923b0141cb970bafeb07ad5cc48df5326eb6ff741174549fdf1f225db049ad5ff4e50220c39e615a943221757aadb48832d32d9dde5c39eeb3f003e1259431b61cb9d5e88a099da0eaa2990533b1bf0d6df29f3cd8b4bd4219d466f84e2f84ed8af015dee20c84fdc8fd40268c5212424620b0d4daa21e9ae71555d033a84d14dfe58923faf0a97b3325b3e2fc206a22cb67022edb1c82dbeda76a303ed24dc996d22a292882d29082183e373d6f23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3175c12cffa61ab7fa76104fa449913f6b599cf0b4a9d40c52f50ae42dddf644061794e7863ce1612a5ebc4c3e431a731c0e2a01a56a6c8a25e7eefd117936eba31df8e7c13b5e3f0cbc4d263f59aea6b484bcf11d451a695f2832f459aaf626f4625a75b5f1918755fe217c647fcfaa4e074c591a06e3373d6c97ffbed61276d8553ef5e00aec701b30ddcc808328570defc2e5051a4bcd7b8fc493497dd483409fe26286fb06348f0575d63c444085cac4e67bf97f74aa8111fabe1d21135e3a228ac46df609938a106ecc2f2f8100433c06373824a21e6a253292dae9108a2bcf68a404bf1a06e3083489dd4a4b10d7f3f99ed1e52b4e08687105879a4418fbaa39b9144678aa6b9cece449cb2f417e38946c7dc68bbcbbd2ddf4b64f76ac2fddbb69438afe27c9cbd94702873cc8a8d491a11b47a4941c21fa16abda121006fa9fae8fd65894621f9221d3b67583aa93236fb2fdc74bb3fec199cf099a3e6cf929626a5872c639157ab8d3535f8e4518647032182e54261f719992a83c8ea59176fe59a44b3ee582d25a1b5afad81e2e791fdd5a2bc6921bbf98c821a938a54a4bbc00e3d2d268839616147115e1f2eb56ef8ed8bef6dfef3d3c7f13440163ccb55446031f24066ddf01bbfbb9f5e1dd3fd0f30c2eb0c796d5188c20b4b6a626322680c66b057ad6bfc767b9011c33da6d30c7c918331e14124c34e39c114ff2460b8776028872b3703fb9d748fda5faa0ba5484a547e8e05324e74f2a6f651c613afeef90b5e4c091ca36099e9041286c2474734cd2cd832720986803720e93a850809096c0236ac1063cbd89e2367fc65a285d07e12aff5c1d01d0d9c1644acbd7203ac0e668b8de102366791624d203803069f574f820fae0e2b22c8ae3c7c7413a28d9c7c922dc4191c18bd41f94c616c0276777ff5ed955d63c0b8050faee90b98b4ca0653393d226912462c88fc4623fe8e75c8ccc44f606d988a98930a9eb2f9a7045abac896228437b19695f9267b996f58620f1f1ef700e6f2a1639b4886d8cec4acdd00d84b2becfc74900e49f4062b25074a364cca2dd8c989ee82fa50ddc2f51dd3a665cfea6718ef7ed6580e6ff23f857cb2fa222bc5d092a38e55e007d0099bff362f2b4583b06c0f02d2c994b293961c5dfc4dfdf8ca024e02ffc0264013f06b55b059590e5955758197f397af150c9521342f83aebc9bb62184937ac2956ff29f99eb6af75bafe68e03083853f30444a6719e46e8e39177680989e0fb50e15a96f83330c6135a36d511703661e4d0a9a4b7aab10e3794bf8b0ab2ad408f2c09ef56cfd5df5753d0019c11308d6fa2ba2c31cd3a91ef80bf250e02b761439a93d8193af8971e30d2291c960b751493d000b0453271430ccc492a15d07d2981093c9ab28fc6b90a27bfb07b92c6e007837de33c94e6ffdf1efcf8983421722df5c5b649d8ca08ed42349ef7ed9d6d273b4e9673bed6fc65c12ad4a5d2d77e83a3b841030999d7e1fb271930dfe73d472a72befd70584802309b0bc61ef0dc99e8d05247f70b90318f5a08d36bf4f97bdb5f512a780610e47443a89234c2395d5b3a636098e75846642567040a7e08afcdb81ec82e79937fb32cf38e4ee3d49bd93709fb44d4338861741cb27437f054a302261c2380b7979b30c4779e96e3c05d691336159fdbb92d60fb981bfa2452ce039b39cbd8c40c07bf5df68219c369c2cb0efd7790c767f630e835beaf116063039bdbdd612847f9e1200a64d103c471f978bc59db98c6abd0ce1b7bb7e32e2bf5a5f9348ed88bd5ceae24056bf8820b934269736b441aa89720efee4b233ffb81360be7a6ed3a657e438b3e444f348c65a48a6fb4f42adbbcd969852533c484765010269b141b6d67368cc3d21a777f210159a6a67b1ef3713e6acbfa6317989c45a9d5aad0f6cc1311c878d1f26e3b31ea61101015bfb4eccba648248e5df44c8e005bf18d05c662c48175da8133c02ba3664fee6ae94bd860ad37c30ebad212f53966864645e0134bd5767b15d47af4f113a59580da7799b4ebdfc7ab332b19ed253bd5512ff3da84181b32adc8aa66a1bd98c6de82292519021c7691b75f81071d6feb08117bbb441f7cb25352c10f5eeb344d82c1256aeca50f070a8c846e4e54bc998fe2b0983fbfab84715532bb02e2801caaa306ea178313b4084892bec437fbd0df7b2634af73eae904882ae6b8b988213fe327c17d199baa723e558ec67a872bb20dcbe1e4da34030094b9805967347904b54559459d3f4ab11ff7834e545ab0c28850da6d96e904937c684f005f7e1ac4f56d33b3a28c56fbe5d9a6b7ae4f17c0b3aa02cfc32d8c2b9f004d785673c21209f99fd0687dece2a416743f34005bec8eb2390e9c3db0a09c3d8c59221dad91a19bfbf42fd76eeaa55ce9e466a0818474e848e82b76d801b57dc74df0dc71927be9927ce81d493cd36f6a1a4ee99086ca361621f6494034b34c8acd451ee4f36cf224d0a5ce799748d24f7f01e7cfa807089620426ecb4bf0007a93a1a5c454bde3301926d9530b37b329699802ee9f842f6db4bb346d7b5d92e4fff393649cdbe3776caee684859c572b30495fd94a0c2257080998e177440aaab678981fe59e060fdc2aaa6f7418e283166bbc25646d5126fa085fb5b626db82f4455db401f1a2c371a99c139efa8f59930d66af7676925a7601ee3ba3b3e3e91e5ad7775d3c13f72604a3bf47a18da9323e47f4a0bc297c2cffea9abc3b0a81a13f72b65bcd3e6eecd2cbf35031448119b35aa1aadf5ca94b354c5c3087bb5feacf4784ac42aa8fcbe428aea5818e18dd970105c6c032be638f77f3dee0f69e20c9bbffe4c80dece31d81084b8322efd8c87999f07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h171ef328ac75814db7002d4084076ffd8a38ad4e6a1c339a5115d607aacef566bbb2930bd1779b38a4e9ea944622f4335bbe9c0c0e6f9419c1aefc46ec5dc25b09675e405a986ce9683c2caff57f79b51478c06d690ef28fa47ec7e7645bba12c895a2a8ae5ccdf675538f88aef4ff884d4beea0d0c5534d7ec370aa4e7acc9a7361115be6558062e4f4c31ae4d8a47b9b5f0d9ac79fcbbe496bbbcba9e388dcc2deaef7969eb9eacf1eabc6c65446cc7ab1a13baee458245a05c74b51e08ce00905a08cfaed95bd3a7c253dee25e1ccbea3953f42f08a9060ccb4d097ea291878fb0cafb4468253e640da8771b2d992421b31b8cac5fdd8f6324b5fa77bbe1ae2ef6e5a92b9194924731af1ac2b5adf139c3632a682fbab69cacce15ec5a8cf7370dcaca72b9648d12ecfaf0c69762908febc316b9e931d4cb913aaa0df29a0232f438f0236caa6627cdcab2e09a60c1bc8f4aeec35c08867cf989f2117c367876fcdfa0c86fb644b0fc8173c7613e864d1ca33cb40ce027ed84d6bc03ffdfc79415ca1616912d545106d510b05d0aa2e759c9ff383b1ca6f616674324952fc58121d4dabe0e252894875aa5faa8359c300f72b0347a2cdc208a6531dc77cb2f894967534905b3ad9e07744d695017b30738f23eec70deb571e9c5a0b4bfc8181174a2ec350eec671f78b601249ee4189a5249656ca8e45d34f5a86a90591b25c1d3232e531a26a5e5277b0033645055eda4f69a9bfa925ee078a7a3fa188f545a41800d0824797a7c1f72af0df4803b154ef75dec4a98f05bf91b3cf72496f3aa096c2f44fc0973df57876416d18e0c68f7859f1027dc16113282726fc208e11eece983a3349591c00e2386d339c5df725c30ee77191071be57362e5d9a69e2f8e1a0cf653ce0aaa0dea287b28e477354f0ec74d9b9106b607fa10c6eeec422746e836b5b5bf361e2d2c3acebdaca8c8bc00b1fb3a4e6d63be1724ec14ad57cce82d2cb9101abb5f301d25bd75b775578ce017794da60f1b26f59369d3bca95c04df47f9192eda81566348f8e3c013b98ff0de5b1868c474279bd5de0b39d560e4943318bb67e9cb93fb06c17fd3b1a6a6267a5be9ce2860db8469eb63a280c96c9834daa4b046076f48891fb2cfcec5ea248737f88a5c593f5d9ace5536eba449994e19ac521951bbdd25f9e164f6b6e3db2e4c1e8b9435cc1906ea24306d8f2b19880eb5164cd4b455b20746312bf572a4295e1fbdb262d9f7c58b564781f394afce3831f49b21b40cf4b6024fcc82d0a30f2aad1538f0b5dc8360d78971c611b3dcba0df39be4830645d8ece4e21aad5ad8fc8e6dd326de8496a9a679faa4cd0e482aaa87e4289b37ca3c4d09aef151e6cfcfa7a73b415130545c40b5a3294571d9278f07b0cf78d16956faf4bd794e1cec96dab614aa6868a881ea603c29a5e01cf293a1400baa04895b288169a5f60f77522a46574e1e39f18cfaccd487c8098da8c73702692596df04491c836569a48d5b3d23a51acb2d9f1998d66eb339e33db7440108eba7074604822cd08f758b480f8e6ed0b48738cbc690dc779b9cd7508252b04e4d24e99498946775560384056e61791111089514265dc86628f622377d4a77a81f5b18882d2fea411f354e2c2d37c1fa2a8bdb2fb84a0d431d230d878fcb3d7954434a16165e6dcedf330cd3b25b4e713e18bc2817bf4dd00679a1d06d6c7570abd9bf0c3cd58183cb29033683c8104070a4ae348389beb781add53d2fe8cf223024ae81bb0c4bca042e6f547b15c7f9bb3193fa1ff333fcf9f718eeafa633bc4ad7f57ac22109aa42ee671613515aa3294eb16be80d2855b157dd4744e76281860f41eafce9b4313b24fd40e2c2a5099e59ac3b64a128e94e9e39f335e949b79ab4538f9771964987d8b1b0abea58244913ee9c8402da42512e696ac914a377f4d83c6668f521b84c5831d3403ee3781e72ddac6d9ddab42c167d635fef72ae71bdc280e04304dffb3ce12924a99049a0a18edbbf53d7e52b7104d63a16f67e8bf68d1b172d1f80e5b5d6e6eabfd0bdf4c8ffaae75988b88c5c11779981ce79733ba3d156466064dd9458fff4c6cf43e630564ef75f4eb4c3c56bc6706e5e8230ab98a9bceb2ad509c89879ca7d4e490edd3c377ee701b190111073fd66997483495ae6311cd78b807eae284171c4012a23166c25689a4d0bf1137a33692413cb25422ca6fb18a6ac1ea4abca8958bfad50f0700f89ac515804049111aa8118019f66a44ecc3301ad2f77ba3ab3d4f62a59594e9924f5c954bee7ef8cfc71c29458f8a82c35c27d17f58013c2c00731bad9ac771e1255d3e43239f180cff2695a34d14f8763611eb796e0552fa9a5e1f00a11732936e22520f8f17122b6689ff31fae6901629a6fa2e1ecefbad4ed9d23ff15caecc4fceaf6e3b3e6a028f978c0ba3cf72c2de366fc765b42c697023d32454491942a98d14f8b77fe26ab98894a93eb4c6a8c1726be016b87b00ce30ad3e63086e2006cc05acf32f8c917c7031078c69700bcb9c520d6abc66760276f3cb3197d178bd8ed0258575088f47e462df0cc7e547ca31296895c9f4ce8b049b596a4d7eeb4e47be9cd5b871dd1cb21f55e17665fdef61da305b1d90ca982672f677fcf41bdddefc7469e8b1ca94ab15c6c6ffb061e098b57d646d977fad6de34d01f75977fb49d2615e0e337c0b28ae735226d3f98312cf5785d047af267d18a4f1c68e04b16c1a501c3d1525f8a32805ef28135f8970f4fc2d495d9392bcfb64fada1b72bd7e86a159d983e8891292fc5ccb3089f9baec083d8ff5c1d82746f3f936b48e68497e259483926dde765d4ef4e0d8dab15993f88123417d475df839ea3cfdd511e08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h51d6cc39fa93d1fa519990be9afeab10f439f1f94abf562da4d3971cd8e79abac0eed052d9386341b61241086c486197ae103bbac22eaa4629d6a1a4fa9a247b626d67042e1651e6c6ed59fd8f9c762c9bf9b57f951bee9fb3e425f0d013616001b01bdbc194349cdc85dfb06a2c8174ec20ee05af3f9f0a867285dd190be42faa5d01a422bd04fa5f2d30259f21d91f67c3ce465db40654b9c35c81b1e9fba8b3ecf8771c1f437efb7274f8120b7cecf8d178c785c92aa4caf6c94ddbb86241a16e3c8c21d7d5791b9bd4a9b8806041b410d75b9eed975c60b3ee2b09834995ad1fd3b780161c3fd779da5818bbf6b3de91016bc3b6babc42aef9813ef448ed3c8fba6be944041b77e7f47e54e1c811656252a44179ca08a77bc25fe57fe6bb13d45f2d0ca90a7674082955bde2b011cd6983128fcb13a7fbe384e7f58d0fe6431bf3c97c6985211a1372e65d746c2bbdf1a2a97ab66efec460da300fe62b85c84f4750021d822fe8f1e9145f6f9704ccf1863f99b75301a3b6d533c16de2e81548eed1eaff5e3d514863e7aba285fee5c919df4222750703a4761f4abf87f6662d287434ef647790da768d42a9365df1eea5364e0d23233aa40a7fe4a4d9017d17707a1dd6ad3883c3fc7b1c13e027ce6f884ec08a9932502f86e662f17da1f3e238bb4b70deac3d5037fa010bf8b81163f23446938275262ef0cc992b195444903e95c243671be1d86000fc6260c3162f3950d34bfea3a64b33ecdc2ba189bd1cd4b016c95cdf4bd3cba1cddb7e04df0779a86391f5f1221c31b7a99b8111ac4c2b7b54d49563ee5c172a42caba851879805c90127e7cfd1166d42178c336bbbbc9dce112fc6e924eb1e7e82b55192485fbac1646aadca40e509b0c0b25b209733c25f2984f66b14e4580dc970aa664aab0ee1dbbd73cf2bd1bc1aacbd3de22dc9b377a218f226f6dd2ba54dabae050a71a8c8bd11ef493b2581e24968bc0022564495ca5b06a83a03c9ea543be90ad6830bd862066cac7859cee616964670cf5a37dce3eb48c28946adcd64c985bf291cac9c47dd2f66f0a3487179f6191f1c3ba34050cb21f003794ba17d89ff231f32017fec71c659a303d1007a897350d847eae13faacf5cbf6dda42965f70cc477b3787ebd253bf487876ecb2c41c725e5679326040012eb49a9eac33c7abda32c9d3f102510a51784015ef7ee52e0c501952c482b087f82498db825cb5ac22461fd5e7e9c173ac664235de875b49e760c4053c87d1dd9383ce5f86ad69dd1428212df956234e1d5eb965ac34b44f24b172ce1c91f203085d7d712a0791cb0a5ec62d42153e92d0c9612296256a6655e5c6cf331613936783014eaf5d215c8b24d22803d614d8da2f82c2fc4de4eedc2b77cd94276203b6e2cdfca44778e9787ee5685d54da1366c90f4c05911cdede052ee82077f5947a50689b30c8000341afa3b723088aa30e7128d989779292d7e6c863fb56287d469d8ad24bd228e7c0be0eb106b5f2d4265a797ad4bed6a946b7b63898da8e3702e469f932a77350e47b6ae5cf2bdbfd77e6ccdb5214e1a9911f111cc1fa91527e3eeaa3e5788429a5aff1839899c319bb482f519d13e0e5140933436421a102a4d9164a54c2d242f1222656b02d4e3b95b0ccc556e4798100ee91df8932f1df94af604776ebb6d5b455a0b6d38e69a84e8c4dd5feb4fce5501c732b8dc24ba413fccd7be1902c6681eb32f7cff0b0d2537d897a3f7fa2c5a6ac8e296974a489a43cb352ed84a6df76f0a4146e3a3527eac7cf177a3986dcc7f0bd376d2714bb5bac9d750eff7f59d8f074d352ed664677a20872777f6a935122638880018a83b04e909a325d60ff05fce42cd681210573cdbfb7151c9b8b04b520689c13dd02a05141937d582046f817f38f1a0ee00ac77c3d7114899afff4a129bb20a94481cbf5e548abb662604be2daf10d174d9dfd5a4b256c2b12032ca6e092f373e6671945fda3819d2d25c336c365901eab771794b83e7b4d9f61b71d78d53ceb5c05edcbb8a0d7f23a1768a32f331dec4e66916cafb295c79f0a5660ce4d7a2c1c856802eaa2dc1bbc8d6a0674ca52ea1ef6f42180d436be372028bc67b984dbd8c33c3d8c7b0a4ec13fb6d32055a3962679a34095501024011d6b7444814f1fdcecc47ddf57242120762eb6c211f391309e780131fab92058f1b2e4cb139bf08d9a657cab6c7faf88a02c4a057e24bf6ee87182fd53049bda1adfc8f778b4e3ae6fe3409ebaae4cc40d80e08cd300a190a75b79767919802e7c86e47ecd69cb2a3da8db26283b82127ce2287ea4ac071110b1543271d7f6b07b434433bdcec44ec1b20d411b92f01689ad9140cc6aef5abe416bb5536094b98445e650bdf340e26288a30808a0774d515dd016521fc557f676795b2dc3ee229d0e3ac85f2275fb1777b0e19186d8d33db4de255a266c1c8485c7864060809c09866e00c4cf2d59fd58b9e0a4e6800aff0b768ab04c981f60ab914a829cd799a25c8054a9071ee373b7f9293fb592bc70cc805d567216b36ce9584c46a32807cce48404a6a70f133f60553799b6f10ef8c827bca8193ca8445e79f09501913cc0afb0a0339120cc0e48d3b4c8c56d30fc82af38bfbffea17afbba8c1bc3b572338cfabfe98752d0fa9f9f8f5d502a38365a8ee1f8c6bd65931e03512731a598ad213812d6049879fc9ca27cde0cb32a116bd2d23ad0ebf77241a6ed5c34d9094e79689314322b6efbcd079881d2816d4c0a90541bcd4e29778eb366bbc437533b4665c207ccbae04a346233745beb07c7221594748de84d111ca7d775a4b0d1d6847388e50523b793208d3cf901953a496ff68015c806f5b9d8c16f0597e5cb023;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h88d64959145a3e7b3170f127d9e808c84e84ddeb03fee8a698922c4db6d2663c619c303c212eabfe0f89b66687c173a6acfb02c9f4b207f3198d312d40832a3bcd22b290632682d3bbfa89e16aa6ab1650e322a0e92e54ba8e87e29e5e76bb867750c3d0ca8d49d959c857b503539faece70224c9311f4c649933ca94306e8bf80290bbce9fac665940e93cd41b648e8b8dce0c4836a79e261dce46af53bf3ec14a40838251b2f1852217520a2159f3346cee39f3203f2638f5970897e78fe6b01eda6adfa2c322396c92b724d264845d84156eb8b291e4a9a4234f00aff0f42f5c9d3a0f2d75650e0367c7d8c5f3dae2181f989355ab6a9a9e81e5fb138f2d287bdf6d50805e049862dae97e4193a5d4799acdbc9fc044af39bafd1e46b5061a921096ab605943ed98e4eaea91e666e62c674bf8956599f724275e7af0bd2a4c2481e75be33fa895ac1429d3b34b7f0232737ce173a210174078f6a0df6df55e95ce49bdbe0e2ec7beea9eb919678fdf5a1e345bfa036caffc312dabd3dde95fccf6bf5c23fd3595c2603d81e1bac5e77935b13cfc82398a8460dd809b16684148172dd0f531e6ef2b68c7df880d62ad609621aa3981877c300aca94bd098082a07666c8fef84cea5553faa4c5d213970be76a52c5434c55bd804f8e349ecee72fddc9c13ade4fde6206e78c8bf31093052b99c08ff8d6668d2c3f3410fc64d5d3bf362716f1b43f0471e7852a3edcff4bda7ca0f824600cf8aa73255b10e1b29689233732d0943d92cbbbde87b64a99e2fb85fceae31c14acd7ec77938cd2889d58f82f4606600c10af9f4eb1a5a0be601c4f1de47b4390ceadd9c93528d918504f73aa217bff2a0da198a1bb5499324cbe77c723c1305e9e1948c177181c0997ed1c13ede2fb26bdb5801edc1e9cb3f9d4a8f9c02a0e6dff983c253985c62f6c1837f26cfa8a7bd67ab0960bc00f8bfb020160152e36ce41c575f797a36cd171e0a2aead7d14e3fa07095b59ee153a702a6795e6f3b8cfaca3b33c0c690561f01d2adbe9189ce2a6ffe832b1fb5dea3c6e57fcd39ece26fafb22104f847c5affbb19dac7bd925e38ac53a735c894f7c3615ecd84d1347854437fb1ca84f4a6f939b31cbc2d2c232091587396c820eca6152ee298d79197b4688046f3e887e68137cca532fbb6be54ce4b1c3cc8add739939fdc79cb965cc60dcd13b153592544cbc518f29cdcf52ed40f82b0026f11a1907e0081cf5132ce1ccaae64c6950d615ff7ab66cd9c9895a004652b09f71a73ad7bcdb83b330313e62316217799f40bee7de8546bc081b39cfb6c7a0aa31d0a1049e28c01dadc28907d841e7a353b03061abd59e22feed0079cc1ff5b1444f14579b5ad72382e7373219f782d1ae3b68e4df0d6caa51110e8f20ce6ac965016704174284b96fa5a0b6cb86142f5a108b18b1284785ddc2f23e1010fcf4386c83cd06b4e8d03cc049902c89303af3243d8d8d566835c4b38c654322b2e9a5642e8b266034239e79a7497b563fad0cb901af24bc66aa89c040416c852be0f2ba90c6a38e8b7677944bb8dc9b0083202af6c136139cfd40ee32d8b58639ab062aa7e5b057698e94db569c3ae48d915c9accffedd086670ea564e19fdfeccbeea57cbd88c32f0a29959391b736c7ab373211f8442c8888a3f5f15a9a4bce11816d5561d6777683e3eb96947591dd6b92ae43f6249e50badefb3df7f827f6411c7caa63d828e123adab71497cc32fd9714c86b5d8bb2341c98985a7bb722d71ca2e44a85fca1d218d789936191a5abd8418d5f96fdd61c6b3eecc8e71f7c27401319eb30be4be2b572354016d051671b5b882a9f9b3e6a1d08f4362db69662b7b03cd309225936d20971844d51afaa2be2f523609f1b4f54df0a502ecc46545d09d1105b73e1f29a2f0669caa41820e5ca8110fc9abc16d13e27fff4a7aa11898425c8f5280371f700a526b4f8584ee510bf09ed550b777c0674f845828703ce8b83ff82baea26c90a8655b7ffbf5f69a748b0d097e9f70149954eb1cd29a7f0046437b71c86dc2b79f3d521cf57ac30ea8acf9604f585bfe4c82449a067378f0aa1acba3e66c54234298b404cbbcf486e47ad2afb4d723eac5a70ff162ed17dbc72ae4f00341514c5ab15b0b1997e15a399cde0f75efee71a1ebbb9fd885c2708d0922eab3d6a02f8035343c8a20435a98b1b027cc9113b1e3a071b4ec6de4b1a9dd0c095684163dc63cbb6d0f18cb7b9eeba91e79fba51a8e71d83c30323e82d2a9f521aa2f580c59548d9ffb30f5dcbd4385d6eee0de87838fcdda09e892856a4bf543f6a10c79ce4709af50f99b28b4dd906142a0065c0afb7cfa7ed04567dc6cf98743010386a2b883c8dd371aba70298c8a13dbc871d493454a347072efb495a010b2898e39545c6690dfba52aa384b5dd5431d6d0ee2901cea79a49aabcf6ec41643055ff6c049b827407a05de1d2439b600e5f55c957f3b4cb44653e66b7f5e85156c1c8b3d5985875f37e926945e058272ffa0d98c44a9c78043b536386ec24f5ff35eb130a446cbb5148596faca3ffaba0218788e6e16b959338b4d2eb2c3a7839fe65d452ca3dbdf2445e62bcc0d609233d31b10514632aa4c8e0875ff3b8ee08d8c54c49d058c9010a06afd3fdd8dbb73896d2ec3c52e4411cc29d19b1a896ab8e4b1aa2351e8ca741a2d2022a3668b61b90ee3c41b6123fa7ef352f33beb23ad4ddc472978d7af8cd8b94de21adf1d1f429a03d5888e36bacdf8410d9648432a1d96b5099a9ab194112534adb077be0f5d52a94b2c43379d8fcba035b2c4a83a1fb275c5f24029cb633283847c99cc22aea6803525153d573d6c59e237b603fb22ae9b7f07d96acff04c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h48662a05a4b1ef703051f12cfe860e6ce1ee74dde6d09c6452866a554e4b4d3065f09a4abdfd1e40ed3911e0e7d816d772fe446f82aa6538a580eb1391f927c55527ad671ec581c84d41a8c815f19cd07e9ffd08dc65f755611456f6112297383814bcee29f12945058a6391960bb2354cee15cb7c2bac57ac282d616b8571dd47ed16dd5506734e1d0df82a384f27c0ef88a5417fa990d5ae8ca0afaaeba41085b3b736e133cdc4bf45b82a45130435a96813d905f666145bbb9bfc3f04b27da14faa7457c9f237b6b1f2d2ca888beae25aae4c0ec6a8f00203f36d59cd873f6d3c4112026928a3c763b27520bf78760c328a879a926acc0142f9c8ed7f26db552f8fc56964402087160c3ceb2d1ba8541f4ccfc001d3fbee6843d888614ce74bf5a0b4907ee07e3f9bf3b451b9fdabcd4e4ea4fd27b305e902dbfa3c753478acd10293adf6ae940af8b7b42d279797160fac36ccda85477d965614bf5711ef4bf506a99fda41f507044fac6dd632c955edd12f47d0ac5383086317460d1727b3f0c54a93c6ded3e55907f22c184628c6a51e9425280066449fff7514304417857a7beb507ad1aaeae8fdd5deae24db440d2aebd9fdd3cf7cb5afee5a6788ab04817d5abc617532dc6a414b839c06ffed84916a1fc69b9702f83d17b4393aab34afbb17e05f7f67ffd86812018c7c397ca48a006471f2e425e7af2e465ea52da838650da1f982cfc262607d76862b7e349f53259ec1cfbd13a824db77b892134bd0d30558d6da2a5128ebf1bd254e55b17d9ee4333f08a44e4a0150fb53fdcadc4faca68823024db0b6b5830a4288d11eb132b5e56a0647969cb68187bc8dd21844e04bf1a0e8200544b2a86048aabec85e1bf6dd4f9caad07db131029694f59a7c74d4653d9006e0f70d71dca96e7261ce17a9816b878e0fd45a9c1fb248ab293377a4e4119c58eb462074be0dc253d0230bc938b2f9dd0018495b2a98dbf52400fad1017768fe27de112d6c669d85b63ccea66fbee6829e2274e774554305e8a7e58e00f83b742a47e0536148f09ad999ea7e7305319f2fea9b276a50785abef66547cb1f60926c75469d9cab0cd90a9e3023019c290e5433c9a1ea911eb69e337d44b975c87ae64fc1fe056379f696af59138e0f88b15ba7d61919630436152845a5c5ed515d363ff4e3ab561844307192c3cbfa695eb1004bbb86474c63e35fd956c9fd00c7343ca21f486f1528a11e513e1dd74540d4ce055d9e90c6570490683c923fdba5b8b0d12821dc461f33d9679d9876a15ac2c4bfa603b60fbde428d904a53b427f46c8f1b1a3c27608f3f33f945127f636b37bf674d555ef348334ad4cd631cd3b16af60b51e9582a8eabb5650be656f17a355a3bcd42c7ed004d7440a7bde513f02dc1c7e7fda063ca876f95ff593feaa6532b1761e2f3a00dde126be99a89aeb441a638fe09c943bd3e362c47da86b38226948c5e8caadcac99d9c7eeaa2335ca7500eaaee9a3e66e3be3dcc9d343202857a571d90b068710bec4ae4cf2d587e7568c7a36e37a69931c3f9f204cbc0030a768a97f3ddc3df91e5bfec61dd112e178a7b94617a40542886275a7a40539a30ea3ca0f3bab6048e3ca30562ec9a5ebaf5dbec08a86ec1dc377dfd4fadb5edef90b3baf9c82544b2ee7113f3f09a6b051609386eaf3e2be7e4946b73ada6060d912114ec526da60316374573bd2f5b3ceab289a8dca7f58e694c87b868bba8b2fe65bcc5449208d368ac6767b098e45ceb3be3c92f05ca720b93f8ae40b0d7be54aff92dfa22e8f9ce25f75cf22c1b229feb3e3d496d8795d5dacfee2e5281f915ccbbb4d6c1301ba55b52ea98f7f0a5ac0cb1135079c52daf26b4b6aceee54211d5b6643bb807c56beeb21df86e8e6554b9eda4bdd21ceca88ce800a85b8d614985aa8f324986f20e65027a0c95da9dfb537a45785894ab88999fbe135fd8c006a3fe3591f5b8413037512955cc90c9841d1ce838b2308375ce30039eea586eed62e839a1856525a8e332ea7f2d01210670e782fc11a4c9734cadf92040f8c0f9452711008b8a80d544e12ca75f05ab4accabc54a78bfead1dd171582c30e0965ebb783e4eeff60757ec3742c6cbef0bbaf10599af8eaddc837ec7a9d9ad6a0ae4a6131b2695d4b297cbe5a4c26a2f07d240fd77b889ce87fba9e1256a86be10e47d31864b9349aedd8fa0bf70e577242ac7d35521a92211e52a2cfef0c5b2307054b6401ee54a9bc38daeaede02a3d474225ce608cfef046bd4d01cf2186ca7b211c825a431574f06e52394ed7de0730fa2db2a23da6164acc1bcfd0c61f050ce80bd5082329d7b190c247323c90460c31d255ab2cd8bbca8215b64c2680ade91eac4167ab8648dd076e6b80c4b415cef0eb75a39e70f72c43b190889373a1788730d6ae2a37c11b5d9428d4eaa2d825fd62e73bc0fef32e45e49f2375894e295467664fad2dc9a51171b4fb993a789c66e9ad5c7743f645de1853f9ac421cb1fb82c77f88e36a3bdde3023090925cc055e10dcfeb6bbb7d56bc8bbe9645d1a383d9a73719cd96ebdd90982024a6afb74ba6af40420eb9e2921e27e12a5d72cd6c3341c670fa2873677b7e5edb9f72d1242bf4e3d094de5231f2fdfae97d147f68a43cd6edcee8685cee28fb634536e929fd0f23728df6d07ac645d6782054f422a7f3692c353d3580d051a91160a410c5d9b50bd2ada0abff83d2b38a09472a91c268d9de1eda0aa766355a81921e4d1ffe4e1612046dcb9cbb6af3045a7f1688aa9cdb99599448efed531b4498e43db89c7b586c93819c00c4739eb62a42afc1f3b1209c31433acadec75584429b7f7e53ec74d3997836867466355977dd1ffa479dd6aee9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h839f5a4a2e4279885dbc73c3bc4b9c5b4ea3edc0fe09ff961df3f7aec12dec422af7cbd245ab1034dadc93d6371c93ec03617d6d9ae86bacf97f1a1c153403c54f587a23ba673cb989cfebacd652c503e02b71e5fced5a3c421a9e00d0f612a3d5420c5d5e248bf4a79450e66e29399874a65fb7a3418a7e3571fa3ec3b8041b245a67acdd5293ca7dcbb8c30d030712febbf6c3051881272da0873822150cd50ce628fc3e245f171477fe686bfe37a049b98ae7c34fcbf3f8ea212fccf5d9872c66a7055166319a4912f9b27947faf44dc383cc1a6a39d5bf97c6f0a8be95be2b454d2f331bdca772e79bf9ca809d5d2d0259a13fd043675c5737317962d317cda52affdb9844e294497e6cf04c1d55fc90e02c8e96834686e7e50cf8ade86e0932f612a7a94cd3661e41d852c07b37d61678f5f8c4dd1657e62f7b4ce61d7580f9747ea82d55f1885e0640f7bb7cfb914819e9d12fe51b1810fc7e04750f7b919f6afc168b9759995e614163e057a631fbcf2fa1c40fd57ae84584c74bf95ecefad18e93b32f4ce5f8a3466ee3f61301ecc54f9c4b3f89f17834f7b1b0856b46c2260ac51d1450b098cc6828e1c196f682a929410886db73c4bc10f6fee96b234448c424cb2f695238569aacf86a4d64c8129fd297e9a62db3abc242d419c73348b71a502b9da9e6ffa82159584a162a8d9f20cbb2f36a85848c8d7e30873b3c274afa4d8d9ec96a8ed7244149404f45ed98fac22fb75175b09155bb2ee1c412e7f033a04fcb2d93b258ebfba303c754d34933cd9a0f551e6838816d8b98b403000cb486498eadf66c225cb2a2603bea93faf692549603cde5378f4e1acc4c6ec9dc17fd220bdb3ef93ebb78758b50f1666820a354f11dc3ed2daadaef100f1151627fc8612688f79498e1cea6343e1d84dbddc48ccc70b981ec9ba510164eb05e644a79e051c0ba29a65123940edaf63c722765b18527d3507fdb5ffca32915e8774ff3430cf0a86ea704aaae938a22a671b844c4dd90837e3567bcdf878de6d5b38a55c74d9a01c40b9cbf7bfc99b54acb9953e694131040b94dd5ea0896244f1fd8f68141d0000853fe952c02d03ef341ca32d13696f65579769de33133b108f1796bf521fcc6b005852cf44a03385569709dce696c3d6058fe9285db3b1969480e06039126e8454bc552844f6cff46f2b30f410310b0f81c2cf2c758f7b7b90cb6c6c8fe6ec3d7198227b64de90274726e0fdbfca5958c40ee9c8a02896cc78d178f572c1a45a8a4301d921415ef935beab5715ce80782e033ad07e3620fb2ee2df2a067cde4494592de87e2f56c8c15caee0e80984f22588019f0fbd25dde4153ada7a112adc6a0768905bb1df6a246e32d70bd5fe1e7c514d73ecfb406dde509b29117b50012fbb33694e84f1856f3cdcd96b28d6fec67b7221a3a10b4ddd3a4809e097271c361f09342c04e112f7d327096af44fc5680a3f35ad32102821ec5d2b956992199c1a10e707702c8d8740b410196c43d8178fdb925613da4be6456b9d05cdfc3431cfac3b1c97d7fa02ffd3d65b6d72e01beffc042e6da7c684a6efe771dbb28a2ef39170f8a76e2aa447a34b5575fc463e5492b5c1fafb413bd8620e0c32a97ae196aa41d81291d0d18a8b231b4bc8de4f747d4dee0b847e08a3064b4606b4ced34a05230997920efef515204b7e75f33e5e9b081f9cfa23724b21c6178a98029db8320d22d8892800c02ba9639f35a44165b40059fae27080a258c1cb9589130369223f78d291a7e811eccbf71c93c9a401c27d514580f33216e980c123d963031971960ae0c69d8e1bde4386aeadb3b2f35344a4c63857a0680b255410b99768a90863073e0d2ba3a4ed9e23bb55888fdc98392322814f741b033822f189b009b4ec80bcfff830671d4ba0a87cc2a296ea1f2d3d430fb9fffe6c014fdd16709676ee180a82803034ab12328366f2f3a1d8f4164d342dcf1eb23291834cd8ec027a3e455e29a0f9be961bbbf20c6f93a6fc87c3b57a7fe983941aeb81b6b41483bb3c8658465ef87076bfaf79a849cc793784c14bc297413394e4007b75a0d5ed1783155435487c04f9cc259431318b960dcac8172e54144c6c771e37702302d0dff35d9c376538934bc0789717feacdade6fb885dbbe5ea462780f0c0d3449b342ba25e8f905fdc10cb722c30fc5d504b2ea650fb3c7d7af55740a9701418ba8f4b4ba14877333f338e1c82009a45c17c7d8041d205174c103c3b3c5c61300b8da3717e2e5036f80bf54e69ee7b5f0c1891b387dcae8e3efd425ac2102f497e47a42a8aa07cb7ec10f67174face8280ce13de361b5822256c20aa61fb4948ee72c0c2594088417535ef502d8ac4f578b4042e4e15398dc8ef8c73c3e35afd7c258969343893c9d5fbe1eca3adcd3c6670a2b2bfe78dda20fb0876a2cf9d0c6872918cefb44ffe339db42dca82c088c96878ae42ad5e60fd0708521613eb269131d634ebaca4c507bf4443f3ab246387843228442f25f7c0ebfb1d4e3fe4c69e279e157ed88c3ad6415a73c070f782ad1231f61b1d336b7a7cc4e0d3b121335da454673e28bc045fd4e097d0ab6797f3b0c4ad9a0bc9b6e5b3d9ebe22aaa303d5df044e3c4c2a0c1345349fd5aadbc885de940f3360e520af013a25ea115cf38c385d7f17612f8ad7fa33ae6c7e98ecfd7c82bd7d2e25ebb02fa5de02b111a1e5676603627fc635ce9a7c5c4cd5bc1ca30fc7f4c505ac83b731c37bd5d1bed99767a3011ecc8e8eebea0581f60b4405ef7b94ad988758b9d9fec003fcbae02eb65dcca495c86ab3425e3c65b15f1ad9349bde52f421fa60a1fc43436ecd6ed8235564b80bacf7757815e2b42d7a9d3678e4715fef23b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcce01999a7031a11df105f592bfdd035291ecccdf7d29119d2afab34f68ad04b9c1b47c2fce07bc8542e08083bb6c31ca6049497e549ef54f2b7bef4f07c9f6fadd6d2abd6e1279fd9ee6084bffaceb6f1ecc10704495c628322d765c39df53bde31f6341b223c0c4529ab111524a85ef1c30ac3fa4d886e316d39ba4fb193104bf0ed27669fb61a728e5cbc42e8ed2226dacb616c80aff01ddb921e10c183f4b035fa674865b422a3c9ec88f09d2eafcad799b2e8c84e80a20e8314603b229d430e37d03c6e0ffced4f1b40da8d31d4161ec0d36beece6ba4ad287135aaa6bd5db0e720410645c7f64039d65cad2af174d899540da6bff834bdf197d048a2bf2e69c873ad22a8f287be52c8782bf0d5a4b94c0e812f749391a8ebc8c3ceb5d2a3c26b7d1e37dc26578f4de297f48bff4b757f0fcd5634a3248ace6b62beb9ef64b6c1e16c728a4d71d0da31db340b6d9ea16996143cee68845a341b3afea956b72a0bdc981703d5dcbb02a557955f65e4499c2e994c0e8a0d75b6d0c1dd75fb7b7f7cad9b8fa9cd5da7897a80599e4664cd3b4e54a29ac8f98aafe21de41f460488d95a856ca0c707be347fe0a29a78a88793b906909040cfda143ecd5422c68213ce163148372452bade20a1b7256564c198a696fdf7e6dc7607ef4ade79e4e851be691b2002e17c008e74777f399e4a0ebae72253dc3c405f796f56316176435842f2b49b374f6f61fc46f60eb66929b68e0db78c773d3a8d7a48ad83e5bcfab5f4edba9e3c1579b55be6fdc984dd43b481f015b8c9cbae2cd17692de93a1aa380fc6c791b1ff7d62aad32cab61068b749ea31d9c2532ba16dcd7f4ee258ec984c400fcae1abf3fef96889a3279188d722ea837436187dd3b38dd2d4f8dfe87a24dc0f84cc09d41f73d3a1c137b88c16f8a47c285c8074371daeba3826455613bc7715bec4140899e666923d8200e0f94f6fffa96e281a903729e526c473ed318f443349d0304edad8b5ae46f0ece618cabe1cc9fb3fee8c7f56ff07b4b391342f3632783515d5aa129a4b109427b805a7ff54aa2e8e17f6aa8329a15dea10ee26a22b3d1a5a6b3118f153d8749497b5d754775ac2d763647b46eeaa240027596bed6b706d78424a027d2e91f6b42ce8d7eb875a45a7998343395d0b2ca983278c2489fe27f0e78b51102e653447408f0a3d7f1467ac93f1ab0067205e8a2d1b1d50b24d3d8a1b9c8719a743e763966ca5f9b28e79e5a50705f952bbce4b036d446b7f9eb17267a4b97469b2862a82a588fab0d2491fd22c797b1698c58110353224e701f3c7baf419cc3b6ab54def2be422906f23ee3cbd0fe3f9ff56de9b658fcd2594f08484b7a0a6e8f89df235ff735692df540f5b534058698e078354a565c289de27cdc1e8ab9b099df5f56eaae793a9c31191f0c191cf1e1c9a67a304a12e403803548bc7901e03fecf014441105268c8f9559f732a3b4aca7c8b80e342d54af6b10814c1bc9cd95780ea7ac4169d2c832e23dcb1e732e86d5bed37d276e4828532e236e9753afc94cca23a61f13ddcc8e6d56d1aff78c48187ea3792eb78eb667cdf23e896dad67f2225e8a27051df6092c4c9399eb9e3b0ca6109ae17e4531e38d7e64fea7f28d1c86d6ae7d58041159286900a31dccbd9ce7ccb70e751317240b80ac4f17e8adf0c7b700cea2b840972dec78a7e949e53c2321a8a8c25fc50b515f36b107f826d6de276180821550f50355741859ac1d260051d7a1657213db6ac289b57c91269a104ee29a105fef1a3a13e7f01de336ad458c7ab8ab45e2eedf22237c30237431dcdf797e71cc52121567bd15ad9f8afa83fec8ac0743a297249056e9eb501236570c07b36fed24b9712ae79268e16efeb7af86571e3835976d7419ff3799600e56b8ca36ab93d23f0ba53affb7f57ebdba3c16e38ce0c4a4c6c3d2fc1d53ea518c274c94c8af5af97ad1f25e22d1c78b47826ea1a9f4439e429c984e2a15bb96b7633a7417d9bff4668e492e512dd06437a434828e7332487ff2ed0c6d4671ec6724e9482a9d1c7b8eaf76a3772ec61847207e8024bbff89f4b429ba282ba64687c38a7e254b24f766ef3a900c461ddaef95fc785bdeb7b576f8873728ffae1701ad837c78ef929cba56f2044f7864b966c76fa2cc4f8563a3cc73ed12a8c8b4c88d45319336795fac360f7f6eeda0f618c6b268cff35d38b6a3cff1cd74366a67ac654765af2227c41e18395a42c9ab993862db444ef0c7c93150e13d2f7d7b3174611a73635309bf220811b7d902ae0aa2e653530812a6e7567313a8047bef308da58b0ee1bb67355ce454972e462f11851adad2deced5ff4f9d1400db7a834a076f5d27bc867fd0095302fc928385ee4c9063febfe290e662a827b6c662e58da040a2302d5fd444189ce7bffbafe5ddbf2696926cdf159f3db13ec4921e7af8147719822f2ca092186f860dcd0b20d8fc582c51e3ae399489ed46712ac59bea64044ce7c17555049c0b1b2a2c3a100ee97f4febb2c4fec684cc292fefde204c25ece0b21eaf76d582ee80d57964c0d8b8b6829d7e24245b89257fe5f16693f79ab2689d530dfc67c7915e5d90d87939ca762f6f9584981eff64ed50d0fd887f9d8e716401ec467a7d1117f0acb219060e3f291003ca9db7609d78554fd45b1c91159d4acf1f6c28fd277b17944a7445f97ea0d42589bea78fe9166390eb73558c452257c943d7e7deee187a2beeeaaf99f1bfa2635a0eaa13f24f16892f88f747241bd9ea7f15376ffb27e094d95c3339a49f8f1d35edf36760e961cd2ee93f4191daa754a472cda8cef186006b2ab42195610ec59af1bfbb464e91f0ec7bfda9bc93e4741fbc4a986c646add8f6643d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he45ce3a99c9dcaabc58a0664bb95cfb25a7dc62258c633f63ce91d5e3889746f16161360fa2982c2a520674d1a3f13e0c47ac7689ed82da756f8f7766364e987500291db714d402df39b5113a0e527f932d324cd0cfec136ce0e4f545021b012a593bc95541f729be7edd49ade1881dcbc29ff49e0fa4197e4a8d92778f18ada1b378439dc76246a94fd3d192448526acc9412870fb30377f3f7eaf005862e918c49edff32c519dcfa67e52fc70c7c8d78e478461480f85748600db79782cabf580c81c6f88b3f7a0765ab2a96383d46385c9d10c45934c80c0babffd755be4144c181e385e41bd15e94d7767426d34adc4e118718c5f9f66befaa5ce92509ad06f85b755b8f18a5bb683da44f018007e10bf0530a2e8bc5ce7a37234fde3fca97536dc231c5635296a6ee32ae1a750e1435d0674ea7709e25fb1e80fa5d29f258df6707e2ec4c4b3d2dec00a6d40b9808542032c99296cb527d8656e67503baf8a257093d9925bccdf80057108f53910dfd22c0b72958f63afc0e80794273e2d4add2025d9a64336345d2bb25ad594e9c8dba9ee89feff2810a5ae5de71156af8b8db3f3d016ffb69bd048e08071a3835bf53910267212dc0e6d025a39add3393d077b4a7bc2821372662c094d119c583e08e7b68459283f9dc2cb76fc3962701c2ef682eccc02c0b3c0e79524887a85e243526afb7011ab60bfa3d8c4a459bf2608000d749a64fbbfd7a8a6cb615e322868ae4a3d5a9a9b084832d0f137476e2367db494d6243b17ec5ba60a978426a1bb69ece25560ecf96bc189bc3b2b365618162a86375767879c82145764b752b7c8e4c1262b73a01450afd4e501408e6175ccb9d45ba49e493e23fd07905b8d2b3711da110909832061a9d7304c60e2085c0f4dc388d66aceef75f9cee68842d3d69bffaf43c9a6513c7007b2d857dac702601d26adbcc967a8e34084a063ae3e432a1337352eb92fb53526f51f0735dc11b71cc950276b44245bfeec0f534c0ca00401216d60c026dc69370d05ecd7d377c2bcbd05c4ba5e7f23ae40a0c666c79f8d79fb94d36acbab9000f021cedd9e6d384a543ed97822b511c75b8e4fd180fd9c36ddfcf3e9283e72b32add97b7c59bf5cf1df1b945074c53794441e473edfb24bc0df7c3790d105116f6d70dd0cf00b6cd5f3f3918ad457baf50d6aed3da11c81bc85bc667ef83c904249d805ae9719b2bebc64e37ffbc1825cf70ed22f9f7f793a72e5659c4be5d6344393161d1a6941b3162b410eb820a546009a15865c46dbd4b45f61e567eb4f3f5eba900d70803c8a8d49d1afddb9857bfd11de84517392d8c3d9274ae28c1f8145fe6db72f7b4cc09c378c3a7cd1af9d3bb5989a3ae27212eb99300743aa7baba2690bf0e23fcf4d57513ba0488bdd7faa509edcc5186e6bc12e20c2c3c4dc5248b3b64345de0a91bd01e7ecda11dd5f3a10b6b546bcd2fe2e962383e6b6566277ae730ffe2563c21229dfa34c2d3e3c0be936b4c150772f51a70c9fe71d051e17a3b11383eb9b21df9b6627573a4a1b9e0affd943a3b0924b9488049ca813452e3b59504f39ba4331b7c35be5471d2de89bae32b0dce389ee66535933358db0e58068531800e9214598bbc7e4a9e2d5e96d481ff17845894fd5743d51509532476e01d212b9ae77d7bf7ebf115c45408c7f808a73194bcdb441f1ac1f31aa329f1d4d9cc25cb621e2c674489ae786a80f272f80d4a57f9be2549c64052a210e3d09f7bc5c93ec96d628d10ec21e928444ef90d44222e070aff2c8fd9a72db9cbd338b608b86b996cfcd94db48c2719921c782bfa4c1f9c1da94aa20f24975e8784520bd483f34c5cadb0f0b07e09a516afcf5aa3f44fde0d9341bfd46c55e129eed638fc38b3e87603f6c8ae112ca0cbda0432630d5be2cc1e390f98abdb75adcde1533d89bd411bc53bef40d32cf0e60b591a055ef7710561b82328c2143431f89198bfea31fec3b7f9914573c8f38bd2e8c99eac143c7677a503ed504b1eb81259505b9cacd214c21e76925443aa535980032432d30d67706d9fcb5a25cedb87f9a3baaf774bad88b1393b7db12ed7ec312522f9b150acd96f77910321565514a3c0ce866fbcf61015d5a7aa97992add58266d9c3f67e39ddf30dc6c51567b7f2d247d9b5b1b6a292aa4386ef3fb056b74b478896e99b5636693021a04a64bd8cc308fdba1b8ff6a077608186b10c60cd86db10d737ad7231f89997bac2dc4d9513b97a1a684ef8c26ab4df505211174eab0fa0fbe5c136bff133e8033a5bb5c67d8dae748aa75095586e561b8582a9d0b341c0655264b563e8c0628e0a0905e1a347d369467bf9309c2195fef6fd38e888217740854e5c669619e113eb12a3df3e53b5bc50993c12c3600309bf1c0682b2f71e6e5cc536f1ff542335ff5e606b43d2400bdf0d464ba3e3df76ab263adaa29102aa70ee3596a1d23a250cb740f17abd817765dabc2ab1d377cdc935338951d668cb88c79ea7b049aac530f7a5ec5c58d8535731eedfcb771e9545eea710665deb3ddecc502d7625bd1eeaf0ec2960fc62b2b91281d772dcda9a54cff9585caeace1b958c0c148ec75cd5f7f3cdac2449cea1d8af28ccfd03ffb98d1713b316bc9ef6a491b0db485027b9da39420619c5a98487570bf2d4f70d0ec5536d9394a3fd97cf0ea25f7dbf06ac7c51497eab993c76616b6690fdcd30899282ef59c60822dd181abf515f4f8d4102f8b01332672c00e056e909acf978c6908645a4edfe1dc684d8d6ea86af6b4054d5df3c50530c11117bd9d1230aa58797a700fbc137088e2366738272bdcc4abc0f057b6648e106c6223e4674fdfc7f22e99a5ae75b1bb7c102485721451c95b0ec60f5ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha4376b95a7a745a3cc82fd6855ca5c605f1565273421f8e169a163429f0812d77a129b1fcdd09ee8b4b124d9e84c4a528e1adffabfe900ef0ce4bdc97a93b7dd2e5ff254100d19df540f2a829f82fb7e3c50c305dd9865cbbddc1e1adb30c760d153f17ed97aca8d10e671378ce2f35d1c903c1d71390f2c0499336eb5323573efb4e0603607090b032ab7c3b949056d9253b2af99ae267605f5ec87017d0657239dc9980546f5f5aae01b676816f15d3d8a7910897b09c7fb1ceb6a1363aeadad7cd3629c46a6061dba2a6dd7b123bfe62a97287e0a954a70aa7d495e9cac55a14dc325f1425373834a0622085754720bf68f06c0cb090ee93dcc4f356e19438a5e138c4195cedf49c4e2d4dcf6bc43e43f9290225bd2aef16ff836ffb214f59bc6deab7c7a385cb101d79450e6705fd2d2030e484fb251dacc430d657813a6aeb44f5e976137bddc0f30bca53fdc3332da21dd1e18fd3b7b528ee54bba7f301a75c8c7cf3c42ac62a7f06b8800709a28aac6afb86884c58c01afaf347bff36f2bf724d46707ef1e551e91b05c613eddc426a6e006f138289cdb7f491eac8335d2c45bb804a23e582cbecdd077b6966e00c69a11268726599a468a939145fc1e420b12accb77596d91b9a8ad1973ed061593b1f7e969a45642443932fe81b72034191a95519ee3093b59c2b25eacf34e86154eea539757e395eeade18f16ea94a03414db63834a104af0ed1b8d5dc9b71cb3eb96ddb46ea43d00b8add4854535801b78241c6646cd19474b12a4071635e29460ff35723c67e10d8acd939941e8da8b968b2e6dda2d4a79be524052868c7924ce684655a87a05945f8b1e830f810a7701d6cc1c5c77e88ba3fe235866d0fb116daf93ed3ac07b365dd2eb6befa3fa7bd7d8e57c2d5f128b0d2efd8df360fbe14c3426f1ed4102b51aedbca278b5b7ce20f45ceeb7e9efc34397c0579637a1549eaed467ec684bf5a59ab98a5fea626683d7b73831fb4ae7b8d3d43435ed960730aa7f269fc2f3e66334fe1933aeabc399178ab63a012a1b6f0e8fa585c6dfe185dc8758b805cfded5c10aa1393e818e7c31cfc08649f5578ddb1e8dc50221b398705fe4f4aafdc6feb35747bcc0582f31c877fd51e4cebb263bf183120df7e348d0c19ae1c28825b77cb0b4bf7affc0eaa9fc87497e4f0b4a04826d1e61e17643b54869bc2e71c330811aed85a0dc7353ff7df6d4568a000d3ac2dbc315eb34165fa706d42a83e2497bbbe8c800be7d87bfa0c7d5102bf67748beb014dec07a5684075c347b7532c2efea30b821ab9a0883fe1bb8efbcc6f2fa2adda49d9ef0afcad33bb8b100e3ca27d6e75b547417d26512c193385a62aa0f9ba3281cdb3b905eed6d2625db7840bd7d3507a68c58c76469698dbdde98f12e194292f27f94c68263222f8fe95b75ea150e757f1f2a537e89c6356c557461159b4561d5f660364a41af80e29eb19479ac8a14a57e16e9a8822316c9d279c84bfc5d5bd9347530df1e0692eb0f12f3331cf0d3f1cc721dd5e5fce480b8669be47b8edd5b79bab11cc167fe3b7cf79c62a611d0378450223877b2c60c1ea24aa6b825286d938936b46cf3ed6f089305edfbf32fc6f35e2810a7790cebac3ed01455b2e7b8650f0e005e593f181001feeefe04dbecd761ab839ef79f4c821bd51e0771913768d47b313b837fcd9f58831bed0c9e14179d9e59006d6b481fb209af491a1da3f2a96a7a920165d7187ccbb8082fc1a7aba8523ccde1db745782703ba78c4293d5dd4b1ae840cf0dcc5275d053b6eaf5e9897f5483f3cb5e6ebcbd7694fdc6b5adac1d5f6e6a041fb2aecc4a8de3144b8e1a0294ae089a95501eeab865f04878a947a9af154f505af92fa82df2bd43142cb81f0c5d1569bf7aaea9b988291bf28220b097a8314e938b304dd97d99e5de09a6d0e15e6ba076d3de4873a618331c34ef2f3af239ed0150964edecbe39d9dd936f69e10f40f51642f6d5c979ea7ee1f2563beb29fc4b682dfc72a8df1b3b2511de60a4ecf57bb1b2cbe515a223605a8d8fda82088ec9cbdb920b289f184cd0a89dc075b1d8c0630550a82941b9b4cc245c7f4ee004e72e82b4d7488f53216126e31d6af4e3b8ddfd87af76db9a0fbf7f2d476044544ef1dd9666fe931385ced4e704c15e0bdac3474046c0860ca8fe174ffc20b00f4e59660ab7c9ebb1d787fe22541d72b7386ef89621987234f00422aa6bda9185d03827817f5a9806c907ba379ba9dfb2e27d3df5a2fc8e2aa6eb93ba5178e5fd8dbc377f4b116845cd8e4d694f2630a831efb2589a81b9c73c1b0adff74ad5698efee4e72b9f929074ddabe8c7b03a6dad00d078e639374be84b6a69a5e002b5f87c8a98ed2d373e57227c9b2e7d245cf95c35cd60643daac0200726eeaff48039200369bc0ed57c98ad233f5a117dee3cd7b4a1220c27732238e4bfa51b859e10422dc2b776d8b3815c22246bf4497f2c56e514246d452ea1f3b5c596656ac09bc50552f6136e8ffb7cfbb4241429f77b7d6c9d0fecd45dd3a76eab57d0ec089d17ac3ba5498276876ec6150e1d5788d1f0af319cde20b83aebbc970ce369fa7d73b845460e1b8ced74f1323f03a1d91a9f5f972935aa5bdd574fd782d1fe1d2cdc179f384ffd2ef0d5f03dcc069f718370f877bece93fd8527d87af4c9d9d8a3cfdfe166382455f156f74c1e928343ac9f75fadfd96aa30ca90f6ff2314a0cf51fbab31fde0c1bafe353458bbed29d53fd7b8bee282397d3d41d5fdff58f36ab74dca7c888205ae80521f3cc0c269d47fd3b5ce0f731fe9469eaef0a516096fc78f4fbd904c49dc8ba612c01f54e2af3fd096a66e75686bef0ffa54a1fe413e76248f445c9c78394;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he1cdb33ac5b0072fc20333cc4189befbcd5586848e32d7d0d9f70d8ccd903a135d6ab133fbd57505b4b100283633f586e5de3b2ba9baef575061c84ea4ec0f4e8ce2d98c2ed8f5622d7a142ae669ff8c2c513136011c02269c3fa15d2054dfe3be6c6798272f68bc7ecabd55450c407b2c3decbc723e8692deeee29615fd59b8d4d94aa49f9b873340390568cafc0279b1932c7d681635bea4129b3335898f6fa002a54c9ca14ed372d058dd6447807b9d5fb8f8329864c7c09fd07a81419367894ef332d7022b1759947fdf819ca47ec8c764274f3f0a5aee0b2b60b1c0055ac0c477dd099134f0e3b6f6d900fc2e5c6c5b1022bbb2065b69c8735dd0304d3ae562204a3c6be6158cff037092dd4eb6b86fc3d2f091c13926147fbc77a7dcce5c4400420402a3ad9287405c6ca17eeecc2efd40f965d1cebe890bdc3bc16aff7f617f96fbcb0be879ad133e309cefafd5d16fc3c79cdeb35b72e8c6cd22fcfbd7456e9cab13ed36611eda2fa7b81846cb04ae140ee99560553a99494f37acafdf6affa286c6d9cc3d2148ab21f80c4c6ed36e9d501d8b62fe3462483c268425ce7849814a5821ba84039734dc3efe9c7c848b120375e080e4da37460ec7bfbdf048e740a175f3b96398c071a9e0db7887b488aa2cfdcff91deaed7cfabdceae6398f446b836027ae1dce55465fe906dd2489c7feb39f65971d8e4fd5d26540e4f7b225afd6d3d929ca5942c0c292f75b2204478c1ceb73dcb784318237cb0dd7a3b48b31052a31fe8800e99bac22265e4421ea486175c3319a6fad65524ddd7653185b1dcfeb4b1fe14968210e7879524a86c08838b0cc431b5a5464e6e31eb837f5f69858631d28915259f10fa37f448ad24446a96d7c3df2d77e447eeb089e295fbab8dfb241dd94c4f6270a11ec9cef0cf1b60ab8c2cf17d7fa2c6f150f551587301ffab0e8ebb61bcc85a2f3ef83de82e22de52ce4d45085c10b3b88b3901fdebbcc3b156c9c366e1ee05b13c1179ab0bce51e3795c26eda47e29529d74d0979a8fe414cd0afc86dc337369e2da64a35145f09fd6e60b80b9d1a7cb8e3dadd597a811a2d434bbfebb91d47fd29ddcb550d43a24fef37b322b27d5eda8cf98d7b437e73bda5c05c7c72b17ca6157eca85b0c452ff50572da102ea0dd3b3ec42eca62534ddf6f457e22363a122d23570a56ec867b775bdffe9deb868e0e0aec1b29bcc75e69a58bfe580d99e130d7c13dec0cd7fb50fc83cbe92e2cf52029b77f2bb26a6d8a5705bdcb78ee4ec6da96f9db433cd991fe2bf3ddb46cb81898e1041920e2b91d1f295e38b46a2be03ad715ba7a5df9b5ba207427335dc18b1dd0810ffaec675c6d75bb8e0106eb4fd15aa0b8dec676a48d721e4febb6cf604a03220fd6c59af9facd04ccc644981adc6deb6602d23f46ebc3ee152afbb19b66175a0c526c3056016b5f661817dbc3261417775c92a37d4f938c10f20d1fa531c0c6c4588cd9a58729a858064d817dcead3e7a3a0e39764ff7380f17f9cdd93a629687cdd94127b0ec6cbfa5d5ead50a149fb9d0d4070c8641598ad440e3e2e5117bbbc8fbef877cb6753e5fc2f45ee80e873af34812fab01dc6f9eecc2d3c086e9a0808d488efee2cab9636641257328bb4a7b50ee6aacdb5e7e5608a7336ff17b8c08ae1aeb856a84a3fad1fc06f48be8f031ce3b3dde9275dc8460b601e501a4a268d640038f0a81bd6e617522e1524df85e201a1238aebe7bb391e5e256d5625271b2b522c55235ff65d010bff7b7a0cbd6736d8cc3d6cbb5c1bb79dbffc0118f9aa9b702cd800e38b16bed025eb0669a4461395bda93fad84f6c1dead2dbcbe3333292486e49d4d03f8a9d70e84cdcd65d86f56d3067c061b05369a96d9245f589aaa4316a24b136839aadbc5269aefa6b3f9fbee6346386286dd096cdb740d0ceea6f474f79729938d46c7facd91ade142f28348b3155e6369ae7c5d9963a91ff330138cbd98abff588c568703e152e17619215e6bdcd02411ec495d396bd272574dc535f4783db4bd49924762305fdf69593e0ccaf9fe35c2292faeb16e33a4692038000295bc32c2ec0038b12923a94237daf632d4e2b9129e7a7c0f9f690879092bce18353f277dd5f0872fe20457fe23385c0d99ff9e9830dba4a1e78976e00f416d1ae447be4770085b7242e919251464db4f7fa9cff6eeb701f8db0e4f1ce170901c48730c60f7f16f0d131991e41d2b3cc5e7ffb0ee99fa61a3960c13f2e6a55d4e65888501cc3b3fbb8af3b496600287cb89cf819c4f0fcb7c3b71da055ec1f54a67fd1a971f200c1b57fa1f5ebd031776dafa7c56c64b473e96cd4b9777f722dfde4dc0ce50c98a818574d7a1d55561e5ed199d6d187ef6c67bdb517c6952b0d20d1f6a5f3157041d25b217bf315a96f233e608c0f6bb7b6c23986514957e7a664cc42a2e4beaae6bc84c163e9f044ea584097f7c5a4592d44e3ae013e72da4c96120ccb42a5e105da5b4721296ecff5f34fe5388c5e92afcd43b6c1da31bbcef053660d7447f8446ae766889341a91921eaf8d0d089417cc249bb71e8a98ad773183999b570033beb8d3dadf54880e8bfb682793ae5f1a6dae50a017887c88a8fe9a8b03efdd1153df3b8b9eb113ab42c062a3cfc22390dcfe986bb9c8c25bfcce808e5bc9f3de3fe2887cc8e61e6f2fa05d81eb39798b66e7af7bc784660b0e8cd6f8e3d82af8f42cb78de4abbcd17263bcb7c8fc1d0a17d9bba0a11ea4449fafcb2b728ba43135f5a4fbcc82956cfc51ef726c73100b3c29dd52ee078227fbe662b4b7c667aee6d47801f802f5b11145ae397a38893ef8c369bd8b305fc5cba165a990ac84ff5305d8a5056e7e8d958a8f8b413db546c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6159741126c783c80ffc971c3a2bf26a9faf88c3e7f5ab02484f674194bc854ad618fb733e799ef3e04eb6a946b40d701b6d5404430b82edc4771a22be16e9b94646b90c7e700d8b897944d607991d66f8d885ec298bc790443718a9a2e4c6d03e623d15f192eb20b919736841ba706393169a772cf55471655b3c295f7e19498f9c87554c8e4d56ac2639c1a760fb87261a3834df121e51894f11defaf501709e8f2133638ccb510bd5da83e4e1ae6b7d0058be9569ee57f2f441dd22b2e0223dd7e4e7c6eb0ffa1cd1f8f4bd201a969f553d877aceb8ccc1bff93e83be7cce00b22f8b524d03be78c3ef03f4f279aa81f29b5d0f89955de13a1593b3d9935643b7896c95c087d27a67e1bc6494e6c37dc2b73146bab1caf96809f244643d33b18ec08974c8395572f668316e930b7a038ff557174fbf4a87776003bf214a8453e797f66a0db4220a9e954b0587a71dcf2f41db7efbbb1d6618c8acc4116740b6da4625587ceb211120a45617d349ae680e0d293082c0320ca3bbda86da8d3a40ffff909fbe3095796395875e61d739c21e7b814ad2925cd9c4d3153b80f370d564b36eaf36221b42551625bc2f80058f80b14d7bebba61bab5aa9bd3ba282f059039d2c7014dd36c4fb8914c8c11cae311b45082e4db2cc3f76e4ab95c802390301403e243c4f9372af168c3a7c3fbf9053c9b1e871833bcf4c76f018484f7067f7c225c689a3f2470090c0418e02a8586146812cf8f98ef7c217220b1aac0369f07422d1a908149fd946532a5b10a5a2f9d5a86a6e66c3194029f526720f99b58815d9b2abad0a2e978f37ac2ad1326212e8d604dc6babc8b164b982b4e7747619b8cff0e11f4f4e39a7a350a98cc6e780f6146eb5141e65cfbe0696d2523fd255119dbdf31f87175e6af51284cc3e5e513a3caa92e0a235ea5e65047acfdc725f75fc04fd12cd3ce8becf8027c9ab267ff40301186390c413d0e0cf26c133933c5b1b43049714548056bf92202149c88c8bc6357d9024605886f34a223ae4f63911c02e784951cf543186aa30c58d2c75287efb78392dc0a8f1812d9f8a491624d08646f2d0d9970631c2ad8fed5a18f3775126f7ed1cd6eb1460e1724b7786d2b92406ad3af3c56ae0690443ad1b3893cf2a6ec7a6ae4e7beb81f09ad0a57f7820945ebbeb42a0ba4676a325031967ca790ad99060e34aaa34c4285940907fe470773c33a0ae11e35dfc935793420cb1711d21f5b36cc14e7c16c3faaf063f6258a363a5fe11ee9162a99a956d76599d2ffa0e678095ccf288c902ecaee70a31a16ef420b813bf590f7e0fa4ed25c81e4843c9dbf314a1177b393b825113aba6489b5b67895d4cf332bb6d230edac9bc96248a4f52dd9c15fe6b2362786f7b465f5fa473fb28042620a7c9cb1249803648446a721bf983cc93ac800e3d7fb0272aa582d148932ad305930a1c9bfd70894fa407904b8a63901cd805347a7534909da4419aa6b182e956ebaeca9e2a78b7bca4287aca34f85c6f7b74ffb53f2d6a06fe8487f41c28953c7e4d4be2614a4b6eb304c968239a0e80dd8c3116b151773e4d2a5cdd474135b85814b056396fdb89863ebc8fa7b7d910b25261ff14f89edde7d6046cf3191b003530d15211eea5d663bef2180064175c78517c94d1370649351492dd76e1d0444ffa14625eececbed5018ed7f0d3c2f78526fee778fd37dd46f3ea09b98a69f3353d7d2e3f21cd018d4cb4478a699e818e69837d4b7e668660f305e19920b3c85355371a1e498277c98f66cb3715ead51febce2be375694622224fdfa2d40d1fe3b612b53aa11502fbd8fa2e78aaf84975ec2fead0bdbc6cada1a8b7b5b8da58c6494a14bd3d3b3961bd8715a13dbd5b2890e00f933ece25552aad437563e0b2fce1e9d76ecd0fe3fd69ab0deed6e1034b5339c81c50e0d758b162b0c4aa30f2aceeadc0fd0da2c826a7fd2b675d9c6c0cbab436e3983dbae07af984db355ad1c5392e0a06ff7edbb35d953f8a7230f56ddc489631d21ed90c2d5e1e2fb0e40c72f72a4222ff3e9947edd54dc371ebf29f96bfa7770c51a6b81a1edf0439247de58e8e3dfcb7323ea25da743a188ad2a0b5ed57d1c157ccc31db7359fb7d4f78e8ad7a7012f07e505b6293ba2988182124a49d637026aaadd084d9e668dbb96b804b80ce1bb2455fcb293de6415af0aed11fbaf084662a4b23034cc522bc3efd03da8b4614bdb8d1f705cfdfd98536d42c5deca79f62ac6cc449f96fa4fdaed5c8ce78770e948c31e0bc74f9c2902dc833ff62182551d5221b44af4dfc62a2587307eaadb257d44508c3a7fc991d9a70e02f34ee771b668deba313a7a02d5bac6ebe95eafeb8e72112a05ebc8d8a5fc85529ca5d6137d1b82735b79eda44adbf6bda737ee0af10bde7d67e59e3c835b9d7d9982824d358cec624ae18c4e04a00c6266739432773183725c083da053def94685b377da449eebbc24ef0128a39f0397951105a6d0a2e48ef441cca303a415f2c6877e71873e7efc95049dfe762964930c3594f6c9fcc609686a0f8c06dbd4b53de5888a2976cfb7a8625558ce955fdf34b86b3dac35a68c22860d59f57e326406255ec0dca8ba0dfdd3a8e13e56509ee5552621ea217ba5f99c571a9d74720b0634c7ba5389b9c728795cf705508b571c97c6d6d2b06fe7fb0f68cfe8a2cd03877ab942e7fc078c4c8e345bde98bd118475df20129728e5bc32ab5faff575295b13533dd8e644de69d9887ff0c691821e1d6e396c2faa9b940b3417b10ade086d64eb282c95928d7503b91a6a8af53dda15ebc65b6c8841a10775e89f8f420c83a59840b3fb4606a67a898cd371dd105a4277186b03f515d6657a78f3874fcb5f76c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hda390adde308702cb706984aa84b22937af201a140a32c4756bd66e4c9c06490fbc39a3c09a98e0b230f00aab430dbeffae81e9151fbfcfbfca47f19c01ece422876b0a99a7451312bbb704c83fb0ac3554b4371c8c5bc48af391037d09e95bc35a4eebb39b2781aa18f7f295c8cb4d843b60632e3d20890d588a44e2d23f0954cfcccd7d0ccdcb67d2b6bce24bb0f06141e96b64a247b6ec116c041d885b18616f5dc48cf99323d08220db5644e11200b44263cae6db88df344c1f2b655fb28769014f832f80d26b2b8a65a6f94ab528615e1d3e56209713e6b2f164a7bd377fd5512068675d85513b4be8b84010d959677ebe324eb167ca3af6e7a9c0a60ca7253f5d8fbe5ef1b855bb0c8243e773d4740ae6d216e8bb6e8623f9a198aa1a5129b37f841b74db7d73d065017bfe0675d89fb7c70ac915b2ea18c6c48c6d9f6bfdabcd9a48e41d6f10975a3dad425e90fd8f027788e6823057a536b614022b61feffdb62a15b438d437f39158ffb6e3ea36ddea7da03d47259957a1d8f61f064a8f4043b8a0294f022d46e3995a5ec682ed9f5443ea5981eba5908bd05263bade0c23d8596cc0bb0177ecd253a4f8f28e62c33ec2b1b4fb619a903a1fff6d6358a8dc3997201e61c9703d6b040d2d4c1124b0a7ccacf5393b22afcc4f130db6927e75f832d7d3a011f32b7fa08f9bae4875b9249134120d09fefc7b412e4141de58c2237596858ff79d9b60a0f7b446b249b4bfc9f59561ebc6658bd0983a982168a36316ff780eba43926f6aee80f25558eb7dd7c78a2f490df790bd9fb87cff2f1a75958df7ca217c83b0b4f82d0395dad2595eaa3e5df40dbfd4780f2a681bf310e3c43853b19357c09bef172d9131cab095dbd3ff5d59c182d22df91746683f73e0fe0dfd3fd0829edb59610d46e97fbf6b1f806dbbea8a0fbd2f9d02a4d0e95dc1230af03e1917c5e8b3599d83ca605f647c6c34f9a262c9debfed6fdf41034ed4f2d2c03ed21f600900e0c40d2136f721993c5bf4ffb2e26dfe24895e3c2d5da5840e380efb9af3ba97c2353f9b1b5a0e64c2375cbe743f8c237be599290ea08eb648df510668c540fc825f6bacc2a3cb394e3f8a97cceed87368b208b00aac01f2915020594504f7b0f9198c7c2f2ff59c6915934418e17bab009d00fe1b7b4dc7b42731b7d16252a3bd14ecbb12c1f5dcef6ec03eb770c62622edafe1a243058db71cc32b7ea7e27e453c1853abb96ef66c56a353f45122418ce8555cbd20b90649221dd71ff8a6a6d89d1cf6f43e91649ba069e39806e3efd2a9b16e770b4e61de8d5fa5bc4761dc0ac29b9de648bc66d691a75c1d6d4182be837bbcf70532841f18a88ccc8381d6f276082f8d51294d880d8afe3668d5d9aef45ef345e043dbc852f069206092d4d51e18293def80f568b4f14986b2e8249189fb4534acfd7e725767a5476db775abc18be23314863ff4bcc17917f9f6c10c81ec9c2c198e42d11c62f5b9bd40cc843afb05fc2b9ddc18fccff90a6f760fe1d7e6fe836de2013552b70ea669ac0b03b8f39251cac9455009e1bc8a2c1194b7c4e6ad10a7ccd2467b6885be9ba7c1f0983fcab7cec9b2f4f26ea97c9990436d8cb5eb513389b1ed3880d87f756274a58c743901061db88d080b39cd11008184e864467d8e8e3310befc9f3fd95095857baaa03cc6c346ece525ac0fc02f73a7cdbbe1d60097d5c8249d7604af29a8d4f0677c0c94116c24bdf7d575fcda4eacb7d951bee55448b16370646021ff3488eeeda2dddd6bd8b5161569976d99dc8ce81542b98d18d18f4cffb29bec481d026e3ae9cfee0671a8ff896ee116b65f7bfab3fa00aec3c5995354ed762beac88459f243724d0ef6508fb1221ccb87d1bc722217e39fbd9a1c98b43250a14b4b4978f5be67fd3e494cebc4bccba3b4c8fc19c3dc8da3294fa12e2a04437b5a9f50a45f99093ee55e6dd66b6e7d8dd0f97a5d25413e645a73e1074385e87e8778a383970680b946aecbd6530c144b28c79c07b204b7df767fbd052fb9d3d15d0223e344f6bb23c7a49937b54f92ba83bed419f67ec7e6c164f8933a93fbe86d9b875285cb233fad264b474f5254fd708b0d39db80bc48fd06fce73f5d6bcdf56c76f35ab124885797d00016fb137b28e13f7b04d313f309b137f1c895a82d92dcaf7dbf09ad6b83bdc8ded4ba5053f1f758e75166a2b866ccc7503be21b678afd5a992f17ce36c22bc19a41ef974f8adc8778fdad72235949d504fcc2ad3ce0cc5199f0c6a70d253d298ce955aa28ec259218e050a40ab3ac8c7cc5fa970932d011368acb9b1282c4e2b76006be4d5ccfd5224b758971c3cbe5d13956c6bf598941045d4b40d464e3e0d65c4a520384af5cc004c25886ef778e580bc6a04b3bc32c38f29b02937033d2dfa709cb921ecf1dfbbaf88cfd2bf8661da20c66dfbed4ad9828b61a57b109ed62b6dc5bf083b6c3debdfdff4a499754fab21dadacedac4cfb71a7331711c53a5efe97e21c0055c81ade7be8154f159e5886222c72a6f4982e642c07fd12be61d6e89fa106b753a28a67bfb6f5b3d8df11e968c7d2b52e4bb8a20e84e3c708c21e96024fda34193586c4ab31bb23edcb6cec09f6b590d9f8858686689261542a22bdfc7636ed68a816ca0f9878cd4ce0fa5ad779ac1d75274ae366023a1bf72d82c2e6357787bbf7e14a134f511866ed79a252ab58de1f9a22a3ddb8ef20f009ac7f7db8df8a8ad6117cbc41e279455034603160425eb5f8deddf08a811a7368fd710696f31ee36469629d16b78172e915a18710436bc3349969348c4e1d2149bc19150c4cdca7d95d8a501929b788aef275b897d0a1225e2bca8b68404bf2f74bf95b3e18c1a1e8607f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7e65208be59d63392113189515f65675652d9dd86efac7a1ff395b24f5a0754654b2776089d1d570ee4bf8d0242917e8385f6dbabd5989da7b34dd96dde8b5902bc1f05933d89c41db7dc9ee6527676447b2ea807a2abb8a5899a43709bff5baa7a8230c7098a3721b4cd86320f1d9e13c78f669a2fec03492bbeeca7038054ab247c6ddf1795017304f4beb0eb3811e7175703f428e03c4b2fd66ea3037c423d24a6f8812d0a88b72e7c139defe2bbc8aa7674af0fc582473f606166c1628fe20dddadaa7eb0db7d4a37eddf820f4b3ae6ea21bf0ade194bfbf1dc961b5752014fdd21b3632ede049549da81d59ef20df33c6af78d5dbef8ac54a70d803083942a7cefd1cb9dae5dbb2c9dd986eee68225ea7971b2c40a608279b527264ba98b27b1dd5380425c3c8bf65f1d65aefb4d82460b1f821b5a810fc074e972ab1c91e185c0dffe537ca9e26419c4e5f6235d7a0cba29bab33935a46a103e8e3c0760cdefdd2ad458a9bbf7a758f20d25cdb1a7d859cdbb91bbffad7a1071e4b92fea1fda3028eaf1b0935015fc1666161391b21359411b09ab75df95620f2b15cb49099cd9ca79ce675e9c2bf33264ec42a53870abcc89ba10c09eb4662058f91e6ab2bc5264252f80be5a7c1b09068ecb2451754cbc3a8e7c0922ec429c1a85447ff489f600f9e6e3337e7365b8389a5b195d62dcb2cb1a1cd33e9036eae115e15dfac137667e7d212f9cb76738fb3b92d04fd146e86e52f6b0a2ec81480868da4efeb8c7f14a8bb7463902dcacfcad03b29c4ba60556891585e2ef7ac5a585e010e7a4b4a1627408656f19783911ddb7b25be3e7f4229014b7294469a404c8d7cea3bbf55004bff659101206125e13297f5c14c7a91600bf2c83ab2c531228233b29cd1565763978dee5792c1ec547213d068567a6ce0546748e3b36afbd70fcef8978b9a4c0386cabdf09bb1d91db17096a646368dd093984f832813535aeca171072a383849d87e6a4287f9ae19bc1a2aad29df76ea186c7abb0bbed77685363e254a2bdf271adc934105b22211e249cff481cc8be9ce52bcba839fc1671c06003fdae2b965103683eca53c989caaecf397aab6b9bcd4c4000f85fe486104677f2f6b9d02eceedf886e3b5ad35bfe4a2b378d9a7ef8abb599468a2f232dd9d5bdf4732b717f9556f4dfefc5f2714f0f683b029fc060671a3de85ead22df95328698abda6b7d285402061a8917e7b4b68ad40f2f9a860d28e3d33fac159883dd79f5611e806970bd1f2623772e72527bfcc59c8eccb983ed2761c79d7f10323273b381b4fa1659af6a6dfef6bc26ac4e293f87f4046f0c65de5b020887cf7962c05df58a9608ab020c5a3135802f46a14c9894506d2fee5e3ebb15ec569e87186f1c127de520a19c234b2b7d9797a94dd208b44010d8f9f9b0625477ccb81fb49b177372b64168d35bc3ff24c0cd9a06cc861f3c0b308c1070a36767c06e533a1e4af1331d9db3ce188a0f63808e9987993988fec733ebb73dead310d18f2fdd4a871ff863fc7ac2ff6e9ca58dd4b426253bbcd7e427a74e11e26353dc4d577409bf2ae115cbc7fe162c784ed1bd02673333a6d610e186789edd181c8b8b6a1a1c3646e9db05f65a63de642667498d5991b7ab900e7efe771191b83abfe6f99983825ce08767829e077297b2d36112d88d6e4de1b1669053e1948f58749a66e726a2a6db13665c01982a76ad5039b5001231e700a5656c84ad3e32d441099d4ac7d1c9ff4aec5ece32fa50c178f348003d3aa7949be0ed55a887121290482b88936393ffac150e40e9b5e263a633a02c2dd8a8b70e5e82df3c71c7ce95e4bda85ccb397184a87a3dd1608f9d01e31882063adc64d8386ddcfe8bd3f4df5d8f61147e942ccd7bb3c1ec96d3090067952aa5cb59ba4dffbb56e87bf5a6552390003088aec45a5dac963b5a51ddaa196063396c3c547d410e1c7b7f43113afe90064c86e451f832f069e30b4b45de2030463ecda95c32b2ec50cc108e22c07ae875aa9fb5d18a50aa38c45057e62677b5cf7a2b782f7875e975d0c88eda26ab8928f4c686dfa854d5fb87490eac7b0884d0ac4afe42a721df674c709e02c022544a6842dc11e0cfd8438e51ec172237422dd8393e906e0f4925350cda9171179f968ccf70814111eea4d74094bb144f432457ef6c0863ea025c8f26dbbaee7873d080fdbaf664bae3db9c77a02e68a516e5838f370077e981ceb628e9c63f001a083b6643403f4ab1d1c9c7a036f7d06f88cb8705921939d2b4c32173a363f1898329dee379ff3174c28b32f10a6b4eb2340b0224241609d7f53aec59425cf60c369e33313be649f6fe2ad933ccc4c046d7d16e209042c60b5fd3d4870f45df10507892f24a733929d11657cf44c139f2dc4b332e1776f9363363bda79a7914e90331f86690b9fd45f7606060867446b672709a16d973483fd49f10bb3559367a861399bab4cb41b8452665a02627e3fbda86b0c4fdd9c05a8e6221fcfde25a4eda708696be6929e1a274c00620f5be1098f61ad00106139f93f69a29d501ae03fbd3f66c9f3baeee43462a1551a4cd7342a8bdbdbd1e8f63a7e20b41e18675f9ea80ee6cd871d32627bbcec4e704b74c461beb108fa71b156a088de35b052631fad1655a5421c613048d53dc367acdfb55a029657ec1a40018ca6afa8705fd2dd813280cacece297e56ae0d946177cbbf9e16faf89ea2872c176d94fa912029eca906c1fa86c603abdb19cb820bec6adc85f924c88e0c39de289c9298efdbe7332fd618c5d4644e0d9441441838c4f8990f2ec52124c1ef4c3925a2627dbbefb94e15cf0a6f3dedaaf7b37d6941ab456485680e86e8c89378ad0fb5400a03d0c6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4d2d154fbbb12b288433851924b0586b2162505ea59ca2bc57f7b86d384f5ba5134b8e00e7e32b5309f36d5118b6a9b91f9a6a725ffea003deae1c8b26e265531129e19aac0e50e2207c9965dc7b6613b9c8afa42d77fa7dedb624c0d86061fff69600f87345fad254785465627785e85a7938c8389f75f47c5217171c90cf3dd05e9a1ca8151a156618bc77508d22eed90e1fb62ca43958dc41d2e1f070e5a6eb4de676ef9065c49d97853b8f75dc0ac50ee06d53e6142e5ea307058257e3342cf8a7d33ed8252b93b6ab50058d08a9833d26a4807cc4c9e00f3cb103d05e1d278f5ba590e5b578a71b048e270c8accac202c23545a0df32e7f833508d9855ff88a5cc5d6f63d06bf42f4bc81b0576fc5922669d48281d95cf7701a54cb34f3d7d46cbffb1fa54aae69fbdb876ad7829b51aaa9ef245762bad79dccb92758a35a798279f0483898542274d8ce16853156bfcdafb969567b39671c778146c304702a4139b863a3abc63597e27ceac4a0e61428e3e213c881c5b1fadf2179c747428148f5c3de1b2b50dc1f8a7be5f9984801ee8ca7255b78502ca6a50265e5d28c4d2f603c67036f3a7c94cba877679d99ed04cd720be423e288aa72b103b0cbd2c16e1e69512e67313ded489666642d9d3dc77eee9822d83e151e2488062f72f7117628becb3aa5571c202a9ce1f879f9789be15000ca6af262af0dc7237b460c54c6978c2e6252e15132e7bb0dceb2adc786340ca5b6d70704d14134a7521d84c247cb882dc2d4dbf541d0600314126467ed451d721b1a090149d911df1de08930a4a5e859a33653405f1664dd8ada62eaf936879dda6a307ae353e1aa981ef3a55104dc485fda76be53e61cf6ffab7bc5f4da1f994d0212bb9439a2d772d63a321b0f5b3d6b44b4816a558f2ee93bab40eb9fa7424bab996e6f13c5dfa9f1ac6e5101c0b12dab5ec803c23f4c2f1e3c032a699c462c1a1619b6d3b75e406eca8bbca2c094d11b735ebfc3fd50441292e727970e4a52688dc74797a6f1173c6ec94f2ce1aa4f0ef978f2e99e356f2175dc2d6233b212d3ed3b2ebf1bf318cbc68772c11507750fc3f818dc7b48c89fe35c9660c7affc17454c06b2a6792e9106a42694a504d0844ad21205c80abb6f66daf306ab5f0730ec0e32bea0d843b8ed8e36ef31d0b34bfcacd2707cfe83f731354a8f58732b459a3bcc1777e05c366dc07abe1ce8f72cf7a27dc59b83b31343cbc754750cf08d8e96a2ba73b72bc92694c0a697976ac5e2ce1a66f2d349f5e8f7f6fbf52d17a89f46071968b07f4f4335020b2f02b05e2ae37c1bad0b2c0820a1d49cfc032cf43bdee289d20c790fccd1e7e82f25dc7f992752db177dd78c9732a0a5938fa297905ac82efc30efd3cfbbcaa754dcf4722ff33abbccc1bbab3112288cf59333d494db27a5c6f84cff967daaa1318c78285edb4867d83f149e9046358a421d715595c805b1e703fceae7826c46a512933d2d4c0a498148fc284e52af8a55462122d0209cedf1019277e175fcbdb18c1182de025e3dd72dc9836abf4bcf10717c50f081c18046b9966f1605845432b4f466e170e1930f8500c7d3d251e8659da330c042dc330f469a95e53e5ab8cbd9ce538f20c5d7123a7219802bbc037bc2b7a96c324b70b69ed9178a04edff2aa4a134474b47784c0584c36afb14cf688cd57a8266250bda2ea78e00a05dec4211d6a51a467b66e13523fbf9bb4c42a13168e33968cb50429f0ecd90f2dff177cf257d2c55489ccea8f127c70e0a8faa7f235bf9a78bc1a42691c6a1a6cd6b4140b8c1077db4039fc5341be03dbedc0671318a4a778471eba2139d9cfe7dce4900fdaf7e9244a7925380850d8b809689803543af3e2a8365fbe385cf096204720b29563b7d1299e23360c7b0d1579a571ae6f9feb40ac374cc179444527d5912ad5c5cfe12fa56d3157c027034626138f474351b3aa29a08676cd0dd7d0c1f2facc72a3edb9e07488428ec9977cf0c4bf56a89a31baff7353291d8becdd4d10f2dcd70430205776cca352177a7b9a91b0d19b38b84579962b4e1af8523d35a04c2ef0169e82cca2b5d5c80167bae733d36a39017bd44634213a5abc35be648dda6eb6a7a2dcc91fd379ec755ff24671994ee758838088c9c12b9cf254d766585314a83dba0bd762a3569bb060d9c573e5cba0ef0ddea999c8d3f1a58dc4b25b07ffbdb7d3f792acb57139a2fd69f8145e4b0ce2628e9016db184ee7c908f2bbbf9996f5d917eb4ae8772b48bf75bbfe87b15b1168e9a6831b6256b82396eb8c2041b90a8d3c709dcf17d44c976e34099bc01916c7ff3d0951392afbc9d77514efdc8da1ca2479a26e7a94e7067d4be75571e0ed1c22f18edb0b44840d24ccfdfc2659e746138f05942ac29dd3d9d471dc70e4c99e461278df70f7bae247539624d71c3df3370d4331bb193671510fecdec6c73f172963f6c03650c38f09fb514403b60f4f8b91dd22150e65a14bebb348a3fa72e98d61e8c78f81a059c891d27419eba74cd737eb6b9d24f4ef9780c1d0501cd2b3c6f483b986a7f82eaac001803aeac696a5624bb116297683b33345869dd03e28017e367515f6c1ea37d27ff31eb75ed327a2f761ac374b7dcb95d88d8711cb4c7a1100a467ffbbb790f84b1eadfbc9e736f743a4f3580409c70deacc45d04316d3cdf87560ae43646c988e57781dce06d33a746942ea68e9e6264fbfc901047c9e05d61a5c3cd0268fd8813c6cfd379ca29cff7d56b5c95dbbdae5dc5552bc804d70a7828051542ffa99c2843033aff70c471ae20254872c3b4786989b68636a73691f667448c999bd0f1ab8037794a2064d30370c1f04bd3df98e80c3ee8c2d886e3a81de042;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hca5766d97ea277c91511aa191f3a0057084565826e1369b9cb99ed070352218a52c4d76826fd04e07fb59688d226f7db7eb7d16ddbc445eb6db1799460d75a3192f78739682baff86ce4c39f23562c1007f56a0b26c49c4b568a7cd31852c4026a1a9faa4099c2b5f4d4a4b3321280be884ae70a2cc04ffc29d1b32a476f37fd771a507ef0f98144157fe384a4459713cd87223b8a333829e667e799a8562abae6b14fb0528caa6aaccc7b73b5a91f5ab3909efcfe68d63765d5c54d53469276402e3930cccc6f7c1a1d7e54e5d71c46f2e89f667430f3308e8710cca7f34b4d84be2cf67ae18c472df0705616589bab076e0f3cbb6f2e24623cd93467a24d6cfb5d866eba083966c7fbbfcbac5570f945a81c15d812ff66931c16474d87555a45e85cbd3e2a0034e08d623bd37bbe7247d9baba49a9ebe142c9ffc0da48f169d48c53007925afe6ec9a8d83c42448604b841d1e7096528c32fa108b6cbe9c3a57290d1e013700fd49c0c5cb457347f1b2acf97df69e06c61cc92a6dbd76cac302ab4ea454dc96444b3e0759e199eb88a3441b184539a085b61dffb7e2d90bf035dc2addb23e0794ff9f1696cc9cbbde6afbf43e53f90fa6b1ae8b706dc797894b02406c77af98e4622930db06cc653c3a943988821db42c25dbbedf457ff1184dd3d6a3a89a060bce634bb237985a1a136d3e3d921d4baff06b071f44844e51f21605dfe01c95de99658b0fc42a59879d5c4306dcf5018c392571998f5460f6818b3eb6e296bf4e373edbc1b54c946a4c07e8b2e583217ff812d30ca0471d05314ef8b2ac109f14340f1b086a8ce81d940d1daf95a47250ba63e894b2ab16e53f1107386e1ff9f65983393ee85a2e1ac582eb1cbafb90b2da60e239d46c8e76404236cf6670657fe7f531a65b5ab871209147f7340da8efcf93825795de546c3838ffba7517c691191af3b8fd0c63b70fd41054e6e77ec7a4a81e3b0177b71678b857c1941b44e31141f9305f1217f77b7b4ec69bf9b31e1c2d69b21aa4ae6d024ccbe14a706dd3268bc83211f8b3caa262c7cbd721a315d2107ae0470bd69e27982f45d60b895be0d37e73e66dd72fda04449a8aa5a75fdfa8a3ef14ccf6521286d358f8e7e8bfcc0a9022d649b3127510649b79a8412f76373ef44c795ad2e5d14142cb14164bae02660931190933830b4955a52d334d1a426c8c2f5891e13dc0deefa9757da64578218cc74424a4b91de4bcd726923979f8a88835a03f026ab40c0f7f21145b8ddc9a289f90db89ca7641309685db62b1c69d31552536d090851bc660b4cedda2c68d99bce62c704a2065ae2e165e16bf9603fca718a4b0800119b3c0d7989b2e3aeb76f5d447328b5913e3db8eec046352bdb43633efe352f998754a4d0949d2c2849010071c2416c2e0f05dde7405b65944034db104a2e5982a6a65c89a4b92151d00eb3343b1def943cf8aef9f54a343124263d38884acc3746a2893c5e27c147665a6b88c1d64f4eacec8ba58917338ffd3134da1af524371bf6dc2cfd455a10fbd9fbec35f2bfa1609b1ec1ea95fa419966a3ab2e13929b90eb64e0f99f5965229639b619ba64a83e7f0197ea1bffcab88ca99ff305877c28da13ad64866c4fd392cfbca241a116bfcdf8bab9e30626aeb3b3dc27301e9a53bd2391b5037461f97d4e2f30c9cf7428a4084c5f61537ed532c32cbdb059875bbe33aeaf6c546d475dabd8634d994f058b04963079c7ef7d1b33a3fa0c01b24c9c91374ea24e615d224389723e15adaa15c106b284b7dbc992df607fafa20381f8ab583e38c3209a1bd9cfdbe0444036c8a4250c079992a9e6c7c2abbcc4329f69d78b3c640e91cd98ec8205db0af56573c1e6711b20a0cb9383c3c90e4f4b45ce2821de83002879f502bb6a027f55e6085090d52010a5e1430c1ea7e5df4493637f4b8fe911c9cf846c0f403d41d86124a1f0707dcce588064734522eb5086d9e334c092baa7506aec0e69e62e31e193e2004ab8ca6a090562bc377e5c2ffc5367938989c936af548718450e55dbef32244153fa3803b6dba927389981a5f8fb4bbc08cacb30ac804158b47754f93a878c5ebf035c953a3744ded2336017da34a83b75468856097ac90aef56aa6e62ffb034954938657b6919ff4d473629c13be5a6b647e913a7d045c6afd5538f92db0c47d13a4f292e941db8e46ab43eb38e855c60545ffdcbc2ed725c382c4b4366691d7a13dd93d27c81370ecb8664aef4584b83c4f1c663d1edecf90c691b6601002b9151a5e5de585d19c4d8d8199d6d588296ddeb6c67ba2bc0f4bc662ce5d5646137fec132423f5627790fb0ecd4ce866c01cece63e728c15770bfe43a795ccfa82a4f6fd2eb59a5d03854484077bdbcec0b28872d7b3d13d52440ecf5af47f6e8b23cdac2d8bea99567771ded38380ea4b93f4d627a3f1f05186a745ba176c7294e425ab743d066a0dfd102b7ebdef71080718abaf05b546a36f37d33214d97b124063f00e1cbf19ebbdd44b34094bf3ff08a6faf9f99d7aa72ee9902cc6e78a6ab5c6abfdc614f8bffecf9565c73ab529a8a3dd2edfb0b967e35deb1edcffef348bb0750666f217abc58b17819272808d564f0788c6ccd314dd591562bdf34862079128fdd8d0e27636d9270271437d8fd3715d646201b57f08f814350c06bde0fe6ee501d6505aea330c8fab7cc0c22a8bdd6ae2494d646402154777f6c4c70d7101a6bf1f666315aa55404360508fdb41b505012037bab553f9efc8e674a74b5329e81ccd28b963c9bb46622aa1ddcedafff263ff4092d52a583967ead6f50f31a87c2f42e707520a5dda3f9a1a6b59c38a18f4bc957066052fd1ebd113fa60aacc225d316f3cbc9bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3a9330e3fd50791bd6954d1c83b89a0084a2d337f4eda817b50f29bdb3d14ccde74e60b999878fef96ca57fcc9a322cd12eadc66901ed449e3f4a2600a5b07bdadd1067ae49da4d289756045d8d4487a767c7713e8bbcc39882ba3898ade2f6875b73e805b8251f043bb322e4c533c35fb4feaee0ec13d60331f1acd2d8d14123c1997193bdd7a0e39ef4be4e91c8ac68795a2e2aee16848cd19317f5e11b75934afc317354161e793d2b07110944d060a0336c4c1334779918a1f6d942a434d84d3aa19ba666635a4119e5ae65bdbc4f22e2f869c87b9d3115da4e45e60dc29d40afe24693b3e884a86db8eb3f5e2b7ddf595b7d9392ebe7e38205d8c75fdde3fc44b596ddcd47eb8aab4c167c6bda02a32b22d92fe35f333a18ef992fe2dedd5d2677a24af03d1c409b99376275df1ca3c4726ebf2d8f11c0526f067b12941d1273211b99b5e11b1e0a613efd4efb8227727f92cec3c69af68a16140dea4e496cca3cc35b0fcdc85e8578f1709b36ce535533d0b9c32f1a73bf91edd18d95e9946c8ab6f086399f8d5fc1bfe96c53408fb34967bd464d0e3e9f5b35dcb907b51a72c4d2736deedc368d7feb8f2017457301b595a3610d5b827e11e548637b8d2857b6f63a3e1a6e00c7236ed8765954e3257029dac48571f271c3f3b6ff7a1b90e68cbc41a122cf5d1c0167199cc8fc31c1a8c27a2f153a74cfbb0a1ed9e5118924449926b4d46076f0952199287531422f5ecb751c5f866d09a8c9db2ac3c863633aff5ed07d324bc0543148f58b12a2d303e5713eb6956661f1f827aa7aa48c85e692dfb574743d8b3b85842c64ef8a9b712e0d9321f2bc0b208a82b818bd5ec9be07eaf9ac319aaa05aa4450ca6b58c43be3226769ed506f2fc7c05f729918cdb7742b52d16989b813590ee7fcc050df73b65d5960ff42dac6176b8f579f04ac670f97fad6f4aff4cf45eafb94fdb9fa7e29f71c117e7c8a77e0e94c9bb6fb2e54aafc1a8c959af35f8e083e33899267ae6cde08cd2cfd644c9524c711db93264f823f7d25a4f862b8300df75606db088dda7f267cde01862cf7140a3ad51ab543cd2f493e464bb3604a67b7ced8237afff4267f116deac16c882aaabaea946a48a893d958f8a0b4c9b4bac2bfe9d4e33b89dc9b51d34f065f139ea75eef127744098a0d365ad2313a8bd13b45ec3627a60fd537de8214ee506779aa15501f0989bc3ebca7047f2dd28bd31f636c57cf973e709e2c4c45d5c567cbf6f8e7cc7f8d74d1ee1c7687e54f043cd039d43774eee9ecd28112708fd5cbb7faf55c19619e30e35848f99ae272beb3f26339589600f40de3c811e319395ad26e597a3e3d34afa5d6cfe74d026d4d78ba6364f1e6c7773b21297db426bd7a5909cffab819754a3c2250d200cd0636f5dd8dc437d3ef6e8f8e4fae44999e983ee8d9b9e0b43b525d3eaa8b806b433b275a2901bc2cb724d9e86c96c490b55d1825e4b5b995883b5aa2800ab1756455b4c7b82ea833aafb16e694ae7806cf1800088a5c9f1f6e42347697d879ca19f403e71169dd564dae805c72be1ac0318d449f988e6bde557be161494c0bf9190aaef2a76e0d8ad7269ac2512ee8daa9144393b2d55e97c2f2989181d7e418783b6314e4dd7f5f05be2eb9731ec92735879c021d7a15eb089089f040a7b3931998e024303995ff48188fc2e1230c7ca83dd944d42dfe2a983b1e0c8355e64f6c00e60e143389dc03eb19aa62f6f7ce71a44eac1ebb10e4396c373a08a08c300876fb2cc620e54070082ec138c8d249f18b8918cb3ebc61d01c39024fa5898f3605a5a140e2abcb26b638906c7d65b2004ae8acc7dba405d42a1ae6b8c32643f38f1abb8066f365729282650f820b3447186ae694bd3223a85351507f9e413bdf77b0318a41652e73eeb5b20c497a73c4db25237e0b80f9fc5eef999df72ebff8d8e63b6c8efa10961cd813e942a4f76fc63a20526889bb1cdcdcea547408032424672a7aec3565f32ce6e9dfe72fa66dd5171178f4a3a2ce1de29b4ef419ba5799d1976b90ab43656d0c329ae7bc6860faa1024d41fed396a5c009c5ec6d6265a9141b677693205f108c956086df6bc136bb133d98edc2dc2092ff5aa6b464524b3f263cfafae4d1524d9b72884e077534598f04a7997b6dda4df5d425673d254108429b7e7712bdb23e8a7ae28416334654de5d7de24c162c144cd4082084f7d34ca156b7d4bb807fcc483e9d13c458c79f18274e718707125cbb2918417f0ece6376c10de3722d115b37e576e5119e8cee4a000766a111bfce7b2b9f217ae9988b2974c536995c90f1ebbbfcf481eafb47e977de766bcb38a6aadfa981b5223027243b22eb15bd1eef4c055abc967829cca9c26f7802027608d8694844bcaee793ddc5fcbc6e15c102775f5f4f4d0197bd76e3d60b59200e254d88395f6d49387ee0a9dd89e7852b3e71c7e7dde904c7d61c99083114acf1e57c55d3fea26f0cccafac32c60751dec4d437c08b8735f62743541d776a4e402a66c20b6df44bb34b6c87f48af24d2dc4aabf6541c55731a99e4b80fbdd4ebde5dc0e37f67e7c3294ad01756e8b39e686e5150468dcfe6b5fa2184273e4d35fbe6f0d35f759a3ca6ca34a4d6419da3ed87ffb8cb3d8208eaffe547cbc92d85b798281030136569dbd3712c599bb63f880f2b8932b874673e0c31a7ee71ffa9e80c2334894d947c882983c88a080264cda12a30beb1414e5cbef6a7d9b53efe2fd7302a2287db2c14adf07c88bfe1fa2dcc6398e2a47ce039f199d9050b56cea2e11d63c8f392ae4b99c36b07dc6f0d66bc54a42f3364d99237ef4a5ad380e9b03d2baf24aad7059d7819cc263c220409ab3d5a4de39d430ec3bc8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5095ec387e467dea0f20d8cc7ebcc4e70337fac0d6313096f5909fd5d89f50ba624320f3076719310619326c37d5c4fd41c5c371c4284a010110aefd21aa326186bd4e3497a60186eefb01a88bc938f98996c240dab11906b24508d2bd6325090a82f0f76b76598eb8da8e9d0d279ec07da763daa4a2536d7d60a5433171c336db07b6cfd1c4eac037423812c8c50fdca8e3109a69a74d50a369103b71ab8c746d1c864c51ea80b45359c86c46db983cb7853c06b8c599ce64e11c96b9707bcc68c928e0d3e1f8e212682cad4b539bda2addceedf7d338e3d1508ba3d3ec1d951061c78d639d2bbecfdd35b3c307f8bdae919862e0b7c6c71f8b0f83cab14a0d08aaa938b5362cc1da6defff42043b99fca392f2381849fac1b502c3de400b50c78911f2cd1d369373941324b5314098c5b5e81541f323b814dd3b512d5070b5d685346bfa97fb83a6a92c809c33633a836dbd2ac6b03fad6af36367a2061298a4c6bd0ba543b3261f42ae0418ed15527277eb9f22670b5e788fe13ae561a6fee46aff0e6eee9576043469a703810a09deefb3b620ac3efe3aac40f9b8cd03ecd80746f3ec21d3d2c46a3a56e4df719d377d93eef0a77fb22d4432b217494b49d0425a065446f034b26d5b70f561fd4bdbde8ebd1eadf6c0be2e43deba911cf4cfebd27f73127bdf77d43f5e547c5dedafe1347d6fefec0c0000455a5dd18af3d84473cdeb45749f66fc1ff66e35f567bd356322db111e55cf6066cd1d1f6e210029d23f9903d44a1b235253bf874322fecd0af843dfe2b406757c9602826bb53742422d40ea66e6235283bd1c4af939a58b41e7ab44e0da2bf5aad64f9fda4917e54423e2e25d3baa7b00d687912181b7bde741dc2fa5a972ffc57b2c7b64f14c04e9c168d8abedeeead37954ba2a68aac0e7e9c97a8635a1a15b14140396a7190f5ffb7864805d55830b05b3f39ab6aafd483f09d532bb5c55e11e067fa988364e484ec44a8131a2a6853b01e04e1966c55e8c3cb774d781c4140bfcb804a6fc01a3fbeda91635c4ee164ee49fba21fa72b9537cfe5889e0d5cae0b3fa805578f4eec727d68432248d0d3ad69e958c6cb0826e3cdeb6e35af3563ad983d83ccf1c7f801d16a0dbd92ed3f270d4662a0c6571f503503c6a164883de61c99572557b51e5a1434bd2f862fca0d5e08f89030b8e1084484a42a8569e3708f55c001d0b7e9df4dcf597e198e6b184ae54d6fbf17a1183e28a7de474e0308167562f4d020c6076a9c9d4f362f532ba6954cccea944ddcf013ea30709a2e4a13eda182e559cf52dff7f4053c9ddb8d327fcd17b26a61ca2a1cd4ff810ae199a5f53a6f7fcb6c0a7cca2af863abe511e7339f6e3a71a5a07acf6c2c8cc3c9f898346410812d5bc424aa0eaacf8dc797651371674969a97ba098fb8c274cd09986590d5880b920e8aceddfbe8f4d6088a58531218cb035021fffa19242963f240f9fff2b2e4d366438475d5ab42c2d3047d292104ead53df4e9b20dd1242777f5fc73803d15b2e8c587c3a878ac5370a6df35fb4846f7569a0ee177eff8b5a4b0fb8a64875b54fa47ea49311868b449001f53a7e709be7930026ff5b48bb58fb8b3d746df732744296a7eb06ac654fc45ca016f5f9ca3ade07fb7a8a0d0aef0299872b506783aa7f24afce2ea7de44370689fdd1e5251072aaa0d31741194435c231f88a659d53914013efe45b8b49e5424fcaee030ff94d6a9852bc37d5305636d8f763d41d7283d9138cfc57b6f09d4571c17f92275f50027fa7013fc693faffc4fb169a66064c65f097274f4726c6a21f9bab7232e86ed25d7a7c26fe4dd59cc360e245c6386f12cae0c97c98473929082f5b4b542270dd95d89237748fbb19434772ede2d58cac96647af211c19eef14603a5a17c5d3fcff26be4f17526761a9b7bbf9ddbf2e3cc02362b1a028ea9b5416e0c7dc4416fe44c11760ed67048b65d0803cf447a895269b149de616228ff74e636111125b6546fccdd1b48d858f8eae8b0de6d05044107ddac18799df0dc74083287e0a6f1fcdb3e82c117cd4a6686abd6114682c4462607d562d566f8b56824f1bf4403c805f3fa3d2e758ec5f1cd299ddade722d497871251e36f7f990c65d54e96d6c1ebcb395b48c77732c945fcb2b180fc53cf0a27611402d77b1574d144d4c2ad31d1e29c8bbb0c87c632289adef7e0e31a3a566cb67e4e902098f3aa27c9196e46fd3d7ed806eef99f46fc28428947e84aa8f124397b7ee06e46cf8dfef04363393c29dc162ee376c3604773cc39faabd5d7fa876630fb44e68486a9ef82a454621018393dad6caac26b16c0873076bf6b7bf03d1180850b6315b33759557bc412f15a968cb4fd19ea5a6b4c7522d1dbb979ba62c4bfc89c72cb128491b600827df8165ba73176e38b27607a3add7c8c52cd05f3b59eaef21d3d71a266746aed82c35a64d356db8251936abbcecd9752aa91bf306ba2ad6e5d0daa3a0c244de1e08dc9189f98833acf17cfc6b36967c16d944f00ea15dba5083d4acbb3d54c75bd668ca1631dcde7fe06491d7b809b95357e0ef0b87555a0bd53d47fd8b51065184889442346b2c72e8b61ea3a7ab87ec14e80c2385a0afa31b87df60a8e6de0239bf008513a6a9d0c1a71b6b00e675c0db94567a4498ce3c8c3a240ebe019f988b36f37dcbe375c14131fdf859f04279d142cf79ea6cb251c0a024922e5f32bea9245d74f0a888c8addea96bf9262cfc1c88fa0d7b5682cd886902bb5b438a3ec8a43519677292520ffea542f2492db57e89d72ab9f7ba0db22582d11e7accc19df1927b3535967bdaff401ce8338eb3ce11151d1428a1fa386886a4d7d867363322dd2e320c90a2fee50774;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he54f7649631b57286be736f15146a28afbfc0c1e6446b6c118239432e902c03f1893bb14923c390cd86f9a7b5f0b26a1ba6a092e10f45453c89c548051c5ab3ad818c60a596469969e4970cacda06591338bfd0c1b6ba918e901703d737a592569585e35b943c4f4b7cdb4297b615c0d15f2a0458d1298aaab12434514c87230cd49b43d1dbb965ef150673ec7257c5a0c83beac8ca81a9ca2aa111f8496f2588c5f69b6d165d52525915266a85397270ba3f9c66a336f32f7bd8b49c66ad1e901389b5e10bb39f7f3c5aebd385348a9e9f87a38c167c3eca039f1add476ad323f2bc92815783784972662ba35d61faa92cce7bff7c42a11350afd451cd666cf758667ce4a59fcd98cadf6b3916216932422c63826e4b2410e10e1052cce15aa0383ca82d7e5e4cb967e012666272c92d71d3b32e10f0d536240cb6eb8d583592bde53e8d5cc9cb60eb56f190fae6f150a38eacea6f4a46c0d8270d68a4fbf52d7b0aa46ed51b7b4c662d4aa50116db3655b44d6c7c66d8bfe2ada0e72c45d5d1614de141023674d19706e3f0c4e749df0f8b645eeebf44e580ab390e2c4eaf05c394ec052f503f3a1256ff4004bdd5eb6d66a12f63d056112195ba49610c1c5fc92bc432d7e2f99b6f1c1ac69994bcbf7d10c1e77ff0f5d81770b3deee41caf33f40bbd6e3c976ac7494f1aa58653e7d6c482a84ff5e22107b25019a90b2f61bf4765af011b66dcb990967bf7d75b960f75769a0802b0a8ab88dae7ca8c9eb3fd8ec2379eaea89094d7cfc1cebf7f1c54020bd42a19a0f824a42cd55ffc1d519f8627fe242b3b1be619290d9231be8ff381ab1232dc4b196a0a97d4b4d8ebd406729c703862e8a2ffcfc723a358b3e6096c4286b4b82d1532f8c6c3620e02cf5735a343a2ed5f2781705939611144b41db006988cece2036d05365000bc8232a319affcf8ddae01a516fd975c815cf345c15d86f461383a8df8e156905856c7b666624e9bfb2930ce7fc8d69f39a049504639a3f4646423413f78aeadfd22bd6be3eb58d8353bf0284fceef653a74f1d286f9ef16e0af3c3f8253c4e979db6922c14245c01d87a16c59f5a269e8f39e29dec2c335d2ba3764d927716119a6229e7fd807b408605edfe6d8f937cebb826e05e5a1097a231727bcc196ccee693af27c8cf2f38819527252fb3adfe7ab115c2591218c4b69bbeace92e4ba61eeef3d018c5fcfdb7cd7d79cf54b3d7c1464302b733a3b8a579369337b01d2189cca2bcabbdc73bd6a4cca77f0eb97872eca3cc1e353c8192c8590c489382a250e145c927c3d6426c796aeab84e9570bab980f789375bb94e64e27d1ba93f17fd7379e33ba527c4fb736e970f66527448ff010c7f4fdcc4633a77151fc0a1eedc5316b3b7af9ecd0eebe3b4b0e68eae531107988ccbcdd6bbf93ec188056dd9f3cd3acbce329e42cbaef30c7b2d21bae8a88a37de925924e054734fd4ec2d907637036f8b694454348aeeac9794347dda383136968f1d407ba6edf4d2da84c146d0f9d753ed8ad28513b8532f5a73a5bdd2db675fe73d3c5ebddd1e4aba0895f06b0f46655c621e8167ca733d316dcee15672fb0b9257a0f992c57cf590e359e7819834229dcbb5c4f90de4dff8ed5cc94196b06d00c51a863152dbf49758fafde921389752399770a02d173ebb86bba0378d183989688af016630acda5f06ff61b0b4a99839cc2727993547ee6670367c7144f3e66c608b306b748666fc22f593f87fd43fb8ee2f81550c20626a2e2015e1a9b091eb7fa7ed385ed88d0763587bcacc7ca2e328396ffc0384a79b788642df97edc03edaae251ca4078fce194dc174c71dbf0b8059766dc1fe8396ef65e5cfeb177a9c77c0662bd4b8717b37d2e5b154df4a674a4f23ce1a62b6db951c76bf508f43174f6d6d12cbb094fe0a3dfa592994b06ce8f1026ea23ef1e81811995797d130b353d42cc47fb4f2b4155206688f4fe74a1439c8985a0ab892b8e5dc40e5b0892e4b8e57eadd1641888c30992d93f111e1c3bf5d734ded79f626440fda3a70cebe0dc53b1044a1ccee661f0d3026dcc341d5acea87ad94bdd6f824f0956a00c2f7efbdf26232e4b91e354314b10fd91d9aa030aa221941f54816401100d482803553eac6057b8ffa49efb8fabb69c983d6b06cada5d19a5138d9e2c4e9c36c7df85c662ca38542948498a075b1c6006f9ee8cf144198a16f86888bf6b50bd3802633bdfee2238e7f951b8927fde9512bef8d306e79a8ec3450403f4f8789c75cc3a0727f19d86cb369d231da11851455312e9929e23b058d18339a8f247110ec596df27b15ac3cefc1c228f2e37a02716e5ec8b1564dc8b548f1bac3f87bb60d0be12e2168d5973cfe038933e74b044dd80952ee96924542f54fad291e9d283dc9cb782de2d066517d3de0befa9b9bd3ae810d55ed5b538da9773f3e0b9cb0f4725d0aecaa7e6b06403ece1f3a4527e6f9189e7e57cbb83d6eab50872131286e15d984c7c53604bb102b58302f8a61c9c870ac5f2a888338d30337cd39d1ae9f086766045194494c4a1f7524160516ecd94e8eac3934d3462ce8b4f3b944a6918894df807766c6abc9eee06a7e930c3929b305fcc0faad8637317d7df1ae97cd5284b09a581856fc865badbaedcb87997bc5e4827e8fc3f416eb5180ac297c41773e6fb6715b7b5a186cf0e46fd8dd6268edb057ff424118c41ec9294aac643b2d61965e8576df0a963eae6687c2834f79a1261bcb9151cd58d64377d1d80371dd89975c167f317ce9395011a7f6e1e28b3666be494f263b5e27bafc0a0994beaa487171ff9449f08cff1944326eee047725e73f29a6a4ce805d25fd974657eb28b675b43021f150f834890e1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he18c3d3f719aa3b5ba9ac9e3f172944056ff3a3340c5667d918215a37f5ea65a98ab7ec28203dcc0e0cdb5578a6982d98edbf289994ad91f3d65e4bfd0a31eb736f04b5799fdc3742dc01fcafded6dfdd4b596f7079715c19af2feeb5f6b15431800f2e10898900431deac9716f0deb865ca5c3f0a4b926939555c6a16a896e2b62d851c201e4342a11ebf82a09e8facc56a2fa6e94ad9ce94055e6d16695d54fde17a2c647ad222009ae2dde637f3e47416776fbe9e700e2bf8fe8624f56db5a848890ba9920aab14112e53c5c89322b7ee80887a3b5fcd09229af77c242fe515e8e1d5b866383fbb8aafadfa31a5b3c33ef08b109e08f98dce1254f0e1f1a6ade98416b5f74bec5194ed55f395914abbca5c2d9446fc5c085cb672746d883beabdc5c4d7094bacc827a354eb6e4531b22bb35aa1cf882833eee3e2a8bbb66eeef75892eca9fdc012135e5dbb6ae123ae02ea5d4c1e8597e2796ee867475689c5cd669f496a2484bc394c086a879af6f38f417a130b13fdf381965755a66cf5dccb4f589663354e0499c22077c8d3bd288840d85ac7f91a14d0dd904baf0f3185952077844e2c2276c1f5c73b5d417d2221e81c646b93a42b2510b38be05fcd313a2586803f1946de3084a4caff43a9d68c49dc8fbe6b75433816dfc2bc34f4e17d01c147aa025e55a642007778f9bc61fcff3ab2f1f2710b36ac3ae314c79427c56993d6cc1a4f7ede4752ba8ecbf4e055579d8b6b580c9435f5d89fbe65ddfb81b819ec56dc7073dccbbff5d66436e1653e853342f33d0f398b47a3393cd344f13abcae670c08001872e3d764b471998f09bbba13f48bf4d7a3f96c924fad9b628545786db57e1af106dd97b65128b4c8baebe3e31ed3f2b091d8c1911cd673d0bc6eeb2ce993bd475934648a90970159e50fe2de945ec3d0efc572e7c8cd69a3eab4af52c8c74bd1cc973e2bfe96fb81e8f6b430b652cb5af9bfd83274e5908bcc1c5672ba99e3637846825cfe34b87db0792a69ea0b64c19d5e137b8cfbec73b2141022ef9d2801b321854290f8b75344b21a8a6fdb14dbff6bb57dcc9fac7b78bda4504e991aebfe0e3824d8e238f741c79d74aa26004eceb70eb04a6d251a74d16713a4d4f770c5f5ab37ca38c8b46c8dd2da465c3090ed1b7f7bcccf5b9167da7013009785e6310297a4d00cb59f47ef73990ab96fc0cde235d9172edaeff5e745c054e85c2c2a857c3b5309e5da97e23519c2c66e6a9a227cceafede6448064ccfe0d3a905ad445876115652b25281155720f1061baaea54fc04a30afd0a470d8d0dee534be316738fe389204eaedb65fa96057331a33cee5c08db19673e02d45c6317de4a9de712c50fa8cb92e9a05d31c03bc573320b72d7dcfdc5bee343e85efc1c65e679630942c23716007fbd2a59eda1d52ec4ad2c96380bddf825cb56aa02ecca8657d5d9f249bab58484c52a432d9b1a93b1966b3a7560ac1ee924622236950ecf37b3b5b361053ea47732a3276c3e47fdb3096c7242866c5a74f4de6bccdf8bc147108fce9963fff43ab11d50f2009ba48ac0cb4006d869f5d93b8c06144a6a0e66d06cc30944a7cb0dc8c43d045ea59081b9f50b1e3e1b234e22edb62eba8ae835cc952636efb00455e221e11f25d87af115cb35eb22c56767f7e242f637549dbf9cabdc0da6a033acab95642ce79ae7655242ee5603f2cd6f240de2ad92ef2e017f98f29c50af3bf2dd3293d147d838ba8ec84a3deb17ed8b7436f0dfec8be19f9512f429aa5d1c6e9a782f47d2fe4d5ad347134b7deb25e0f7645448c57c5e5986b446a47d605b42a8cdf5ffb09589ebfecc3e24bfc6dee59ac85580df4bb38a3496723a1a62004c49d9d037852a86d7d5c898607e3f890216582a2177bc8795e2e5129b30ae96de11316fbdd6f8d2330457e3a15eb6e10f0371412824cb41eb9ca78d6f9db97597850d6067e15e9584b4e65e4328aec35a54df287645d1255ed6e022ba5a2afe5f9319d5b55f853aa1f21ab5bbacd4c839b615f4f52e7669eb34e496141a8396f414bb2360c59fde8e35b63b6d439ace038b4ee72e03643f307b16b2559ceebd1de3b7da52a0a6a45039eb2937a14f9820f1cf77fd26d9532600b9d011f87a05b452b0f74fd56723492f1ac23859b1895e509ac467abbfa9bd5521bb51964cf7efbe5e34bfd45a9cd5d66cac0f8fc11eba384d7fb8a229e945172d51fe63abca335b77562b86ee887f16296286e43f74077cb1a8e8731f087f3f98674881a1e60c4e4d8402a1ef26a695e4e83515cb46eea4642fb585a1bc858cadd792b8661fb7d420a4ccc3ac28a031886d4e9148363b087e0210e59e703d838f72472af7a2e8e1b3479b598d4223f81c4cde5455e6c417133d5aa457531c21cecc0c24b928416c28603ef2f9762f24b5c9023be71626b115f2c144028a72109d06df67f09c9cbffe6534a2e739df22207f3fda90b50b616211ca59db598249cfcbfe6b472f90b62488448750d63e2e05b93fc2661fdd311e8addfe9d0ba2154d70f51a4f9f7ac5947005631f9223c3cfa17152ab3b8483cc8483eb0814ff87026126240a74f25205e712dfb1e53bea0c14a843fc728d961c91310009a152e5ca6a3adcfd815a35acbfdfb5b2254f190dc6d7bfe04e72c33af74c281c2326268814884bb5ac9642f302fba73b886e7f3de95e7aa338a8df155f2ffda67540918a3cc8c6af672ac8d1618404da079adda83bc88b82249bc2e26733bb3777cbe8fa74325185c41c3e40e562d2a083ce16ccf4067d06b9fb127e0d7bfd47d93cf8de5203c33b5b1512c5f8b07131f40b14e268e9edeaf8b9fefcf3b80b142e43b8b747200e3c824cbe50e15cb0adaa427fdf453ddf9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcdae507a6428613a33fb75b9bcb5866a3b9946a6d02f0aeb9991eb1bcbe92e823de1c35fd660ffef19fa1455c3149578c9754ea7854ee2f05a123a97893874f7fb622d5c9b68bb2f149022e74dfe11889aa9e9d545beeda44d8ec1bc617722534e711a3ce5eeef0541ca237b64fffe10ea375fe67dbf83a59fd8902e90d0d596f315ae2708497f685df90bc84eb435c11734f2a3c32b4e9bfab4930715a5745f71ff993c018d1c8c80e44fff4ba8a5604232c00236607f4ccca05ced78743b1bb12d71528499046862763d00207d9d17303aea60a0906d4824da9cc8691b061c8e68c07da4298c8960f8a2e6ecf1ef79083c3b0212b8aa208399323ca81fabbc2daed3b423799e542fbc9221c0b85fdcb112a0f99c31c5d61ec780fafc9bbbb78dcf41d56080aa06463f6eb10c5e24fd9dd1507202717a8984f8c676f22551393b32a80239990ab22a47a168b7b12ccce0aa2df7c038ba4f9bb62ba91fe9358e0e5e536536dea2f88e23d477c4a6675b965649f517bb786104bbdf2ab944eb72e3eead964a9ce3934a52f024264e205ac683f444cb3503100c320062183793358a88dfd8c62bd610096b3a1c1e1460edee289636ea187aef178f0901c9230c29a36a66cd8b23734b25b3e73ab459150093465f2bca2ef00243ecf5cbfd219d7bf10d044839e9c61c39a64cbf66782b881d34f3398896424aeab459daa4fbbe00131edf882b9b77d07495f66e7651637ca6f509d0caf6fe68b183fa831735ba37adfc178307a8c2596d5e320b20ce5e28d6be87465689b5b30f133b7bda31761bf20faf54c5cfd5645e29b936f72bf0b914e46c37f7684a92af84b0e07fdf6a1d61a1b7a3db6fc13e1ebf51647943ecd98f26bc5e6265a1f52edbf5cb02567461ea26730edc666f1f6f7c7e752ae818bf94db884c3a18f3f136b0c34ddf140314b7e1d43690913faf0bc76d2ba541e7d510aa465661fe3d9f887dd7580520babc427ea495f0e63a71df8b615ea6dc88e213d4dd0c9b1dc7f607478b8a05301609242db9827794b377d22396a40132b5323243c97a06cfde475938c97654ede32c90a33fde72e3a683903353a9468f8b1807e85a4679f332e0a41ac44a8e0a6a51ccb0f76ce5cac0e4172018c76426c2b2462e13c835202518b6e32ba726ace4105c3cc032a04ddcc851880fdf03e464e484c1d9debe06a747a60c786796b29ea0072d7ac08be825dd3f53310faec97842b1f4af3517aba89d2a0a47c1d9bf1f9a2024b4d92f4abf2d0e839274465f07b064f50f57be101b5642ebe9722cb8744a5a754dedf97b29b9253a5d427aa8165618943d2448a397c7ccc8bf760548ee6aea4311094eae07d4f08a1af6e74eb55c44d64872ec78b17e194cb32bc009260e0254acb3a4bec6294443a4f92c2aac590179c5159e1eec471584333a84a2760a8033b05b33650db9682d8b95d4a30f82d1befacd8a91bbbf29d2b6589f3ebfeee7621f50c98b2e2b2a744071ceb4aecab4e2108217d0fbe517d9fe3b8f4e887e4344fa4c2a422c5362ce54849707330fc7d7fae095b2563c9fe7a501ec1fe6b288fb6d65408f82631973a4eab534cf3ac8968bd345eb6eda6f6e5f19945f34b4cec1dc2210b612fc81985566cd4b0de2a6532b2addfbfec5f5efb338b0c2460c1ed43b9e7052ca4a8f36d0831b4b9082afdae3b38829a90d666ba43d8dc5e2184c198d81ffa743e4e76936a20f150fcc566cec24de38df2ec3ff1036e55d7879fd251f7f98f99ae7145c3f10342960d5e11904dad07546bc1f2f16365da34da629ed25473301e059c3aa203393bdf5589dcc61c999d74dc2d3844e14a1ac8491d01c7031695669603943df3af516e07e5019cea8a51c1d72db904cb9c9781c6deb8426f0357277b2b84a8590f4d6f3dfd7c014a7d703aa84335670b9c1de06f271b224d05d86d67e535d29a75e695108ac72bad89a2e9127529fc9f0a239316bb43716c2e5a5f4a9f6abf6f61872d7ec37bebb3cd3cc9edf8b844b81eae71d0a0482f7e1ca5b339181390c188ee386ffe7965ab6c5505af578acacbf65a7b9579cc368a8355390f52e9875cb4bdf2ba02394fed83a7bf8921822185b584cc16fd5f2bbb82f9c460c84eef4cae80568bb7723432eedecffddadafb4bc3d7d84013749eedf62cc15b158a056807f34f1cac2a666f0ea6460f9f3a17fb5d11b6ee022f5360a69bae413b4724923994f491f387fb5cba5d9ea47fa5ca5fbaec3824558f1f4f8f93865535bc6fa9666059e1b11a0d82eae51c2651447053470a599391d32bc22791958f45f298be67746b7ab5d0ebdc311d984fb8a55fbf4941641174c914585e52cad610272abcb5948ad8b0c91f5fd41642dd3c2b5e14926135a7d11625bcb4d48444b9e6d49d0c3c5cb4c4e746c8058a8f3b54f78175f95768deac4f8d39cc3aee3ed103b5026263e367b063cc6c631a55f5c165aec7bc193f4f51276276249dd0156a41d272f5e21e35ffff6c1f29e39943b2df06816c36e6a9992e4f5601c1d43cb98fd0057a91996566a8280699dade7d515c28fb38828e56aaf652ad78e1ed4e0fd755a1762be36f1b7b94c2c2e69465b71c404f7971a30429028ce1c0b58add5f0b18ac8cb6ccf5ec27c5c60e80783f607e345cf1e9c968e3f92215f8d1c7fca4b9cd7829258384070f4e7b7fb3269c5d99c24569f0e1114a12fa6edec8c6370cf6415d243a66b6e3db22bae40b3d3be23f303f436fe3313f194f76e436ba571d34eb6994020dd12c1f3937da9093d968c75a8fd3cc41b3116b486afde893fa92b61b9d75d8d7a93dc6547d622b3b74e906b496e59ddb7058327a6f073e005ba9ea94bd1a0ba882b9e200b6b823e14af2853afb45de803b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4ebc376d7f57d5d9d69d644ed83c215d84460ffc73d0930684c94e121cd83b92a0e355eb66c58a68ddf77801f814ef7c9420819c2795540557c6772f3802416a87a71b2cb5c6db2b2ebcb03402b5b28fb9f190d4274f6e00b43350fd9d5f06c07dc115b5fd16a3151fd34ab3fb48239b9cf595a72db5823346f3c6def76b36d406eb476a5caa22bfedff1948a062ceb2e0c6509360463f4e59ef199886229715d97fe666a098525f28c4380f47a646091a828a2f6202a0a47344a5a11a849dbb40f73e58c115cb1cccb896f58d08874c785609ff082b1d9bea3322b94500e87b02e7009bf9d3d17814c245bfab4ccca612bf63fc76caaf2f081d8800b22e79b8902684aaae2753a42b5dab3ad138ccd45327fe9648fa982fdc2648844d0d584b57907e0f0eb1c94fab917c667ac508a510326f6e60f47e0607edbf19c87a24945954316915292c3be16af39b88d7247d5ecc7bca93e94cb9c286baff5b32c0e8cbe178064c9fd1f3d93c6d8d939b308d52af3bd6fafabe88706d218968a5c5bd21a37991c092ebc7226b159c34942812be29d3189ab3c367e78ddfc9f9f3312bdbd13188ca3cddd519641f87b30e87ef1a2c096c274dc3df50047bbb313ae91672fb09092ac55c4e5b8c15f7fd574ed339230622f1ebcf141abefe3c34a38615bc112fb0396508aa9e10fe49b61b61359a6435ff9d7f1f6f68ced0e1b53b89663e69a2f1798476000a670bdb225f9cf3f26bb50ce3c20849331b9ee57a338c931345d9ef1a54599b8f08418421d0af10addefce21f856f7429f02173a9df3782b01c4267d2ab16da1cc2006a70399b48ab2f2f07fe98515084a6d4e2140c75d18bb85eed582e40f4bd2bd125cbf64d46415a165015cffc8afbe5bc0f20c5d41a0bdc1d7810dfcbefc3fb76e2b34258c01e0f6d4febb50ff31c011841933bf8bc5ac617d65bb5b698ec5c20d6ff7ec6506daa499c74e0116b5fcc55481b421512f3eecbd50e646b736cd771099cbc919572810c03576bdafa2e098440888faf339b67dcd97acee69fd2250e8341d52639f7739fdbb28f5ae373647f681feb3c1fd39970758b458beef5fb53211d69791446cef119cf6c4d007d544f10a346dcba028d1c4d33618142e82de777a0c7230ea73a6d80b49b0f75169335a5320c153fb077702ec4eac36916696707688d87c33f59b8e15b486e8097d3bedf6d1c938f85069cb85d938f8bf4a9ad1943622aa0bb06ff504dc487ea44f31413bd1ea5dd02033962d1728bbab63518ed88281ab2b6a1fcb38ee96835f665be24cc8a70a43628a1214133202665fe399d749f335092701708a66be8a760881c77302ba52600407396cb767c82e0320caccd20c3b2168d680880bcbf9d9e764b188c9c958024a3af131cd6fa5c7d04367c6103da8320ee9575e9fcaa1488f1580e352f0cf43b7409b1ab9881e2b419f66734a1d38b5f3d488d70c4639ce2915eaba3325e77b716060428a57366d6f85186e4e0bcfcec09f9866f9acd4c75bf0789e7c18f2e15e85a6b78794c4b95fc5604452761379b6660bb30fd2eaced20aeb91a3565a4156b3313360131b2cd9db62b8b8dbf19315ea2b1fd3af56657f46ffcd639831497cb52051841c51127d00b03027ef29081fc8e30d7560e69fea9fe25f486d7db42b0fb8cc935548303f7fabdd8488b4569f7f882df8a05a28ba6e76866dbdbc78bea539c85d69750a56594d5394f49f1f418490bfaf04efe4be2718da2c3d5942bfb872285fbdbfb7328b463cac71da67ecbe0260eaf4d84f448246c75dfc4bf13c3d9bea30691d29cd440f694bed5d40fc8f3a4612ca228cd7508b4d491a57ee4130236cb70b368d0eca4b1c9a4c860255e16ecd692861e948de143d49b9fe1c1bf202c8a3f85fcf44ab6ce3f0a528343e89e4ac1ea3c10e6707177fa602a5d9e0d550028b6b34f570b5f19161dca3bb07425bbd65c7c44747de6653aa9e45f435b24014f054039ae1eb11055f3ab009e9487e161fc10454440da406b2f8de35daf5f6b7dd1934c251c9415aa4e3defe11433469ead3a59e9aad8f2880296ee071c6a8c733485405bc1564f4a7756bddbe2bc695f716a170c170269e9754a8b057df6dafbeb8a5244b67d54214c76d6add56d5685b1840a6c1d9ecfd103f8b56c7e0bc596632025eebe312fc30c98860d71b072ff8990b9defaafa923f5c2ae708624c77bb46d929a2e71507fc0a7b131bf83a5069d71d10b01f4395dc87b3c14b2ff51d7246e030bc7615f54533d27f77dd8ee8d14b5b1078dc359ede8b0451824c64929ae88ca10c13337b2da4201ddaee19270368ab0ea25503f6482ddb59e2b5846db932841e5cd4df9b21a07ea4ba8e8d37cf996a24c1b6141ea6776699e40e4e6d77624b06885ce5e98c755e2535865d99e6b3f1a104658c81575b39ffe507fb5b0d5d41ec64db9a2d2cb0729c141bc2536045df81b47ad36055ac0abcf279487dfc69693521adeae5ff7679c30a76fa1f177a3d2157df9c3470314113a6ed9afc9f7bfa6abd24f3eb17d16f192a6f34220ced9d5719e3d6f5d07708eaef97edd765e3c6ca78e626ad5f8f985de90859709e1de44fb429ca36e057c711065bc7cdc826858e831fcbe334a68290d46c79c195bef7d550deb1a70b39b60ff507ec38333ab9ce09f1903a81ea66e4801324aee114d4e463cd50a594dea3feea9c2f688258200670aaa1d5f121d0a058eb396317775f8c69a8b011d51c7b0eb71e8863aeca508645d978772db9f379e6498fb714ddcc2b6af0c9479128377bcd56c66d7fba3cfcf80d663450875240e08e889a5fdc7fb8f583dfd85a3525f8b9cff1a8133355d33bee445dbf76844f0a9392ef3e96421316c108c559edf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h854b36ddb4072d8ca111934a53321f2d4e65f807125287ab6ab9c2126c1a2505c62a81989a4c27dcdba3608dd2031717d7be30e092a341ae9ac527a014a12788034c1cd3ba727a6062edbbc7c292360e8699148b55c2477d7eaf9ace070d57f817598a8f3a8a2d91dedb2a93d06cde6c75f98fa7316800b96f675a070b7a0b5fcee77cb497a112ec85371a91aab352605eb8f798476b7820eaeeb6a1927ff5a812a18c4c1364c8f8ec9e0590704cb09af070d3033c74ac9e4087f4a48edf51d940ef5a209ca6e9b0585d6fc825ffd20b932b38e3ba78936bfa2814dd6fe01569f5e9e027c830c81c1c80db78268530fbc9ffe4694d5f96e15680cec1644c9dcfec23a38baf87119f5197cf1f54cd2108fc931f296388f25e1ad66ee00e4092b3c6b8c21ce4da11c0323bfe4bd2052baccd4a1a9b3c7c622a4d15bf4d7b3a067d96dc1d8e740dccf0ceee976d1ccb97b160cd39b54b9e5c8c8e362026d606a6a457450171ce99712125e4c0cc2a240598aa668b6e4842aa3906b887b8921855f60f0cbf09cf3a59e0585be3be0f0c818c61797f74565c411e068263e5dd1ffce425ba36ebafa49c71c96ca306481009d78f92cb9801ace8cd767463f348ae7fb4db690da8ebb0162344648c016b23335cb6a4163d80c1d175bd8bf93f2e52121540d1589ea022600f514bb3f7780df3621e257eafaf6fdb9cc997909e908bc7dd5e6f0755e1c68190438b8f62ab7ef7517eeafa9735bb07967eb9f1cd07ead43ea0b8827277c3300c275c43f47dec0f52bfb1812a639451e4ab0473d7f6ed1523137268d098b844347e7dd8a61c2d0124aff1b1a60704f34130ea63e83f8b92f2410246ef8798540e890a35096e9665de781d8da78a37ab4bbcbcbc2ce0752c82e7c77f5bce879b2e8c35e73f0ce4d5827e58a9fe7f1d47498f213a396f2768f02b13430ef40cd7296de180009a1fdaae2d80b0d8cb3169c628e98e5091ff1017a508058b1981210c2f307986522625d1e6b24497b0abaac14e703b79f7ca5aa77269e32273e14cbe514cc4e26d61b05a45058ceefe89e0485854ab14a603350643dde85925fca212f78bad5faa7c08bb3bdbf5b283c8a64b73ce7936479b9596ff9ae6c1a4fe56da13f434b923dc882ee8728197deead26e0f4d86207897201cb1f44c38b887402b34f46ca661d9400a09613d1fb021635e0e6a353d0b67dfef041830c77234b6dee6d4187e4e125662122ab022e4afe6b943da0d4a505635ed94a37fac678ecb90d4a109ed791d8c96d7114352b7bfeceba35a053c8c8247bff79207c3c482c731990e953978b98fc0a783ab63187d4a5a87db322b816f0c386d64ee9075ce5c0b5bdc7d62ab1fc98b8f065a8675e47a1aa00cfabd4383a340355bebb8ecd6e5b45f57383fcc3e4c3f3b5ec9449248393071895153e4c414399f219a3813f168c08def8c0e0c91d27cc760b272541c092c998a3f5ffaefa50e0e021a3967206a10cccc121ae9e6f6a78bc51de1bc6b0ffa8e3a15452cc487987ce9fbafe85bcf9937541b4e1dfd3b2c0c0bab952d104f5df0a6d67a340bd0e80c8e3eac437aa8f5b00f39e1c19f735c964e2f4d13981937a3970ce630501686f731b4cfe8d02afcb0d85f25084c5151a7d94a08279ecf2fccd2679bcaf8caaf33198481bc54d4211cbf97022de157c40a0af1bbefb7e57c98a9bc12cf5727e18f99c9a8df9b88d6e93c13a77297820d0671917b3c0390dd562be47449f6ea0ca1459b258008eb10d53e1ef566f0667d74fa168a39e7264b0f04a4f6c3922fb4435f0012f758562204b7b00587b6135604a0d8a34facff0d078d7adcec222d337740ef7ed5da9e48deb99d58cd2db1c373186efad4249ee305bf7539704ee5c7b24ebfc1c9101a4bb38d8c369a50386495bb414dd3ee5ad6ec9b5f24a7c787b69f09833b4a6ef62e914d1fd78ed84fbdc9344b2bcb7629e71bab2a333417e7f374bea8df4385798a8af570ab69ce2b5f21d147a84762232819fa039739afcf1cf37c1a96d533d299e572635e98e6edf3abda67d12e88bc9b9ad8a788a39767f76c4939bb30b30754bc158375c84238a13d172e1637a30f921738c154c6681ae4c3664e9f56a2b075145e86586105d91441b6c45e33a413de1529c004fcffa56da864a21d47baa90c51ad88df1e9b9381fbb11a18fd6a5f47c53cb2bded53a3ec12ac06543f07c2732460be19dd42be104f539cafeeb60c4e11a652f70ddf010d09d63ad8ec1a2a9b49718df19d7a54a3a21f2130bd9487d412da156ff5d1baee90634423c273ddae96f0167d1581361138dea46deb1d81a38fdbcf0eb778176c6dc77f6ca2a04e78532d24dd592b1886e80f810f0f4fe7bfb1ec4e4db9bc20b5301f167de8ae95bd1eead6923b6561cfebba381523ed03f080ea05def2d4c143d1dce794de97fea9c7deb8602617ec45ea3e77e031d2bea1161ea52725765fa962474a7f44eba565fc230c6347af263e1adf03e5dcc01c6606624ff7fe4ed473048ae324db1278fecaf30b5d6d5dc0b8f906f107e0f24618b5b9ac2ca98cf3b9d990eb876e00c3cd49767ecd43eed5b1724774238d9044cea5a1ef9a3945f55ed982e36be6aed21b78abde04da20e9fc261ced6393450177de64329cb3babc0d4383e1dc094467f6049495e8df166c67270c0d490ee98794d6bbfe3894f4f569a15a659f261383902293abebc610afec5d25bc264c047741959beefbb562c31b6d18142f473a4bdf5b5080f6d8ac36b2fccab7723b01edb2a12c470fa4fe7e59d2b3303a1cba254f3628af38375b52c82e25b249b86190629a20d7f0d48b43d93be6441d9c7b9cdd3b85705c4ae5715a75292a2471b6e61afa7126f7f873f120;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcac95eb38981ec6de97b99818bf03d4ff5f3dc4b37811941509648787391c43bb9ce5bdd3cc81fe655ebeb792366979d09ba53f9541966287383a658cc6ddc0ca01584004510250a2d2dc9c795d1d67e9bbc4254225c9e52dc4a80724059a70a3f8200979939de15e8ad24e72567a1069dfccd9dcfdd9c1f4ec2926b57700bf4f9828bda6a1beac8fa9aa50813b83136ad1f41a642e2a453ceec787b6ff5d6aac3dddd5fec60900a68733e33ecaaf8ecba480ee4feef2a6f60410943670fd9f3a81a66a5507a99260e389cb8c1fa19bf7de9c162c57d080a156fad38d29f8d8288cc186a326abf9bb8a59c857968cf3d3a6adc9a011db69b1958749f6a70dc582079c953ceea3aedd3bc6876b49c4bd1e2df9d0c0e6290b4c220e60f53de56903a7fdcb2966afe887d474bd507f330bb906d904d06cb28fa4799a1822ff93ee894a64e8c588ea10e7119fc85a93815672943d202454f28ffa9925f5ce2d874ce4d219b0b545c7f2c74b9e3f7041235066bfec19c028ed1e841faa385a86929beb5797f1b5a1328c94798961aa57b9c012b06fec7f8651c89742e9cd2806278923ab7851b42956307ac81df44f5bf15fd281411db584f2a48fcd79be59b06c1220275f52b72649e82ebe70c1d1bb2b86bf636abe44fbe82be44777ba85a9482496fb478015bbe3d00e7ce6e90f30363d254d3a46b0806b7f55e92ab10e58f8449288ef0a0dd80cd1a5cc59e0c84cce54f13d8a7d90f26326864581be9ca84e587d3e46600b690be13bb3fb9da4d44b3e46e49ee83a46aab5637f7c75d9a13c2beee6daa6b4b7932df3f35bc6d5f431419335413c18e55234b4f00a72cd9accebd100bd4bd1c1f9753615af8ffc6e041f73cb8b0edd5e2f59d75d1e3c97ecfa26bf4fb9e2bac3dafce7c9b1cc9b3d1d1dfc0a39ec91177ce1cc6f48911c94ec01140ee34552ed984fa2508d2eb036c58021ce44c353305e871cbe254547148d1e838c9cfed85805831dc7a6e5ff5821fa50091645d4448acd8ee0ab262f5f48128022d38acb298dd7c6fee5fc9d63dce9a51c6ef5d4df2e3ccb2844fe2ec58703409c3ae808e1504cec33666535d9b8b3228c6bf86b55d04d3d0da915272f1a0a4a50a5d39f498cca68f4445b52a40e0bbb96b002460934ed934a37996d74d99955d0ba53ac0865141a9a42be3e9b025ca18867b607563e2740b7c7a6ffca119e91beb1362437d987cfbdbba8e213c14b85307f09a2d13a3c702fa1887ddc43b8875632a438085ed07d31e990c74a8579cfabe56e475897f84d4dcf86a66e7f202bda7ca0233fb286995d07449c6314f0548434e449d7680c262b4822a7301028c983ddbd1ba55b4775a333078101265bc6a8882d38aeb59d105b0f6d64bebd981f8b772e6ce969f1384322f6c11bcc4e9e24ddb2a8241ab3b84aeb7c3b08f1e59a73ba672c041572896b87f4626c8004a22cc9df8ffb0934406b801fbb00dc93ef23af7fb0172923119e8472450d96fbeea9cce74cd0335f836d959cd698a94385e6a01b3d5c850b89ac753e22dabbbc19eb2f052ef332f2fc1e51976ea8f0a22ebccb17283fc1ee1ec720ffe8ae51d11c1ea83eec1c656b8e48b409932bc4f13d7b0556431864f740725ff4113f2ca4d6e0a45a8ad85a495df559b952217849b03f5df7d4fb7973752438d425a6cc984890abfba82e232a9cac56f1c134801d50911be0daecfc9897af7bcdefc21bf245c740ff3b12bcc17b06aea8c87033c8cf3efc80c15c4dceb5aafc086f9e800d2bd3d9b4cfc97c4afa0d67a85cb9235ec25f359529f09893cb39928a8670400f469c69760da63b0061e75d00eb19f79250096938bfd5285a759ba6986c9f47e1121d1d8cddaad8a6f0edb4acd41899ed0eb3888af90c527fc8f9f4f4db9b86d4fbef3c15be21582238b061cf631dac0746834567419052776f2fa09d06474c1cd960239e011dc67c73371d9cffcb88b4c7194cdaf199b7b535d25e8483e51fcf033728d1e22f07e6caa2047010201d325e810ab03d1107bd81336989abd38ec215156e37b345b50f46db5d4d81c87c80c007c2482251b31a64eda449465a742418011568107bb10b69eac9f7c79837ec7b1299038cfe8ae4374f0c33f7c51ae7585ef31b5aa625fe4eec3d35a22cecfa4844167534c353638e4422cb86606b1313d5dc582e46518b580b2b34925fa7d5b7748a83327a9b584f2551dd2ee5b5e115a1e0fbe643348eb86b4d8e8c5845d551f91fb40f3adbfe1b93d6c145a45b0c622498d434690eca4ced2291576b9249ed7a92448ca8b773dd22c0ef30f22cd31a25d544c7d11ae952628c205a7bfe6dcf7ba9b4930b2affaa5825c03ff26876c40ac653328166d756567c3dc6d6ac2195d8cd9b36134b9d32ee8f845914d001eec525fa592541302e5a5270268024d2320d1316997feecd2577021030d6b5a30b65ec216bf3d622e1ba484fcf675d0486854f0a4d5e9b4865f3c7efd216acd9dcc2f493c9d32f3e3313608a52b040661e30aa44c226324bfc08c11afa461b1a830b21da94f4a7679dc73486db27581fc8900a69738568cd0fc0c1fa7d53a62a4ca7c25a2c950ad554604c55b1649704d2ec76fa208ea28c72574560cbfd9854da0997a3faf6ffe9ec69a9c6b9438c4bd7a1ae132d5e0c5656aeef4b8277dcae9173be14aab9c07e3d9b85042172ecbf3cd6f78dc0e1f0f757068ccf527ad5e01d9c36708572b037f28880f2f42779aa71e37a23d01703129a21050044675496c5409cf503e88605f0c0d7f259a42e224fc3b7915bb79e935960fc9822b87afef3151b0371ed637e45da4c333a2731c385c10357dd697669999bf03a00c9960978d54285ebf49078f31a0b99929e2822c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd5f1bffa89a2ffa717319c2e371995482cdda18945d50df20e02c6e52fa14d449fb5dcc6dd407768e17554f58bda2a29acbb0208ac3391217a785b8e1e1508da89987167a18163ca45b885b43fcc41c00134ce8676a9f77442c7ed86d03f91af51fe931000c0fdf85e14d863c43ba3be7c1d91dc1ed7ffd3c94c3978a7b9e2f96afdfa8c60343266a6b29daaac2cd49b5d03e87bf3dee6e6c39c5526beee69dd97cc7e4f9d0a569cba68fa8ed8158bbb7d011af0774b2aa1dec5b8fc39ae7c6d848701e02b6d4e258820a17765a03d4d63839ad000f5bb827da04e4eaf416c6090598d5400ab6b41a995050d158acd23ff12bd0ef15139bd6d54c57df3542389f0af1d6e3893ec0c54ea54a681e1cdbd24c778e718c069b70c51fe35ecddd0a25a05c2bca751eecdcf00b034de28fedead4e77d5bc944d2ff12f9f90e2f697e811b30860883ed7e243f878e2d2791a863cc36afeeffdfd3483284f745a301e958969f052ef75a67f520679b4c4a1a02ca49328067e08f0c053e3c6971a62b1cb66836588becbb6a856706f857305beb146778b1abc0f36e8640844e7b41988b86e7d8b0129353c67bf91ea882ceda769b8f723738c2a5673878af986ade6d6cbfdcd0da2462cf0a0e5ce6261f19ec662dda93da2621180d322e89cbed54c8bf5b470a538f1b56cb901d7d508012d2cd6fcde47d3a0add89956d7b047cb984d3f633a5c524b76489772bc54f417db2264995d028d1a9885c8318f998b35a5c24df48bdd0b8977dd3d96868f07cbbbbdb668cf74b44fe1109a7e04a214fb79e2b3c0e8334929cb022acd3d10f3ef604526c799f0aaea90f68529608e01b8947bcbe9f99c39c04170fbf15cec097033f3ef251e54dd56c30dd12d5300b96a28c55127146c4c0ea451bd59270453f476b1287085052fb59f3ac4b7d42cf7f60ebe701eb3ca511a63553e97b6f05e3db12b7f3840b68918aad8cebf3e6b6a2d0efd3062ef0a19cf6ff999dd1d3a22b6f1e45f64c06de82a22809ae9e7806cf5224191e12c4e5ce8213f9c24d0b8fcb5a5913e582bdf242fe445adda98c681dae43f1326204449e6e63f95e561995c116c04da323e173869c0f52689381b28ee828809bb7bfca2f6047ef7ae88684c35ecb41e7e9a1b46eba7a0a661ca524d55dd5882daa88cc44a5a74fd588bc68f56c36942f2a5a100f808c7c6fbfac6140e7d2bbb603ecfcda6dda42c2d1e068ef87028e76462158ce479bb886324c41c110a3d701a1e86f1ceeff8ba988394b21f4e0b8a74f62b4e7ce8939a8ddd382a9532b6f8e7f8260670d10f769c4396557ed56a12805f6e51e7838c21dfdf49eb02833f4ebbfe63623c4db887be3dc6348f11a0c97a4322087e7d7387341345752b543b591e21fff2e51268625347e5d6ab01c499e506e38569ac8c31a3b01aeda25be6a6a567dc91f0750a99329a155dac6b62d823eacdacf1809f43ddca291a81d2fb12d9d52fb60f8d11671934f58325822d7b47149f5a5f8cb430b8100343fe0a7136df6a99f8c50a13f11f659dd770003366d7db57aa7eca6c0f7d84639f380f42a0432efe361b1b0bc4a8d7ab67fb19c7e191245bf4f6f6fdaaefdbe89874fd0294b3e992ce114f06847b07d93a691c87fa6a4f345c915803fa13bcac9b480572035aa6f1bfa2033ab60a44b82a57330279ccec581546ecd56635b5e0b6cbb3179910778acb7cac5e1be5673901f6fdb86b8454b064c2c85c136df9e05fdad516ddedccd68e96adda5012830f25f17d6baa2fba00d8bedb01626591ac1aa8f7d6109721b374523f4a6ae1643922c1d1de39bcccd71a970d5856f6a5b73d67b86267c822d948e6f9458d6604d042cca6c90afc57d3fc7b8927d6dc74be6aac7cb4f30fa28cd753f4dec52e492097768a83d2cda5a564f19d37e06c33259a88c3fc3a7b056c0a00c578966c3ca09fcbbddfbfec6f456930f29dac6b09dbb282fa336ef2a16e557d9d84a95906c3d859462769fa03cd376486c57276698d2691e32ed44311aa94cb350b7dc69a4bc170e78aea54e41519c9c75fc70213f0007b0ea6cd60839912e0718673429db2ca567323b171bc6706e470cfcd2654620ca30e965b0f153bc0f3848077b64a4642313e2c5d930745d890a49701a62a44b12070418095c2271237b9aa56fc87ab9373c4769f14be0a48d5efdc17854392d99e4ebec055fb6b8d9aed68d337f0815353274bb979ea0849fc2b1d5fd3559862186e9d93d0c1c4f1bdccbc2a5ac84d059c64bbeb725afaf003d4b8b262d55d9b0f98fe3bdf7d9a4c58e5ceeaf267674bb6249c829b56832480042e27958cecfe2c67730a1ae0c4ba1b2bbfaead909f0ad34183f8e26bd95bd9315361973ee6ef344a6aa2805d4785039e1c3229d5daf4e2b3d07ba0ab674a332dc0923e51ab71e2626f4fc70c6f6add0271968a3a5728fb96004a9a1ddf4aca6ffd511e0d777bbd9a84a720fc00670c4b3a2282c4c2ed96c62be88d83208d13d986dc1457c0e027da81611acd79959f5bfba7af508140450c2588de781f5acbe5385533fc9fb14f007da60d9ac3120190439ccb75245b27722e17ac4ddd478950c396d33d39d39298a1f574a25400beb10a668c5f784b6ebd9ed0f71069715b00a5958904055b5db01461a2f20fd8f6db345f7d78d58a8f81611a4650e8c041f037dd397e8638795c613e050d5e1965cbfce79a0c0da3254d6b848909654ff7332f058db6501604f57973583b7394ffdddb90f22de0cd776f7441a2420691fccac5a905cba101d75118f4c4d0efc26270bf3452c60a32a61a449e377efdfde762f1b80724eaee44a80f09168830424aec47b9398eac6e4f9f5755c581ebbbc94e5cc79ebae422a6c0d669;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc6a30a2493be78180c3a9a15f1009c488ac84e0ae60c2ebf48930b675df979718375e58767053bcf95dbf22febc1205746a85c7ca1cf51028c27b91ca9e9a059fba241747d4d626de3352378afcbc937461de834ae87e290ecd74a5e4e7a71b538f8cfdf3ed735d72564fc8bcf619aa00e7329ea16af2d4564a19acb68ba314e33fb4b49c35d5517efb2d43b0ce02613f1a138b1b56b13c8bd7b946e015dfb2216fd7564a76c39bd803dedfe63bbc73c00d04fe96b40cde655259bc367c852cd3587bf61fbdbb67ba57ad88e5c7384eee220b715d965d03500be894c20ae1e6f16e729868170bbf38bf8d69a00086d0ea5b2a399d8c717c8340d350c6be4db5c3b2904b3efe50c3727d5493831b3bd1c72db1bd62cf3e5fb37daf5a2432b3f250acc6d344182a63580ac09fa2392b2972827b29d0a538962bddf549aef4673f8afb2155325f10ee0fa9d7e3333a92133fdc0c86cd53a0671b7d575cf92c05f09e2609ee77ee0384ec13feecdbffa990fe03e4d3697567f134615aa4e3900ffc16590dd41422608e8f1f92838e5ab11cc96bcf74b89c5f0e0390230caad7e3321194070073838ad36b48c7728cbc7488b9accfd7c8cc20848f89bad8b76df8d5f7b7b0c33805451609b4d367dbd832680f6f707495e3b12ad366119dae29b7c4f254ca9a8490497395ecf3836e79c2fa970eb57915e606699d0ba8c6893d2665fa80fc8a6105be7eee729dbe7d68b784f5ea44447bde88e0ce47e2ac1420961f36cd43df3d7906adab13cfe5a11f440c87e3bfdf9ba8d2d69cf4ad315c536254aba4d66920a280ef5434fe3cc77706219107885ec4fc6efd88217fe44f3d2d2cab4e81ebf610bd4f4a42c477dbcc7cc1b0e3c3e3661eb6d1e2df5e05b5b450ecd9b746381f72b65f45342493a7ccc37ec09e784e423b44aa8dd0ccda7035b1bf64f36da038d0925f12bc513a47d1c123a15ab6222f56226964fd2658a5557faee2f85c19d1ead963c2678dfeb7b13e08b65f69285e441b3bae44ec08561df1a4025e360f5becf70d8e0dcfe0504b233f19a97837e400f71be2415dd675b4a93453242bb4a0437694adf05e61f07d331e0efea29f32abe37facf1cac222378db7667ec92502d1c92b0a8c78c66ce403a36fc2a0a0bcccfbb4805994b6ace802501669c127a9168792f12ed4ec24ad887e1ad22cd0ab89f3b91715c8c044e87cda67862cece4e1eaf5b0b63e4ee212d9253da8fb27522d4ba311c9bd1ecc45c197070faff9d1b270b52d007b31ce04aa3e5411c8ba08f67e2a390e9492e5ef1120dc2607be63c75a33a618e8f87f8bf653ebd6faecf18c09c7be4a96baeeceee11346e12e8e5e7c5db10a64892a711dcda2c428f2d16d9ad2d485aafe0ae605d0df099e3c1f240dde852a5f708ba4308f50e8a97b937c1ee7c8ab682412dfe3615d214b6659ce3506ed0f9d24ff4e699aeece55546ab59abfc880839527d39d19a9ea23d3aca18e22f56337ade89d7121eb2dd89d2ee2b017bea6749bb30c9ce41cce1c9ec9644cddd4aba400ef0d8d6dd55a0e706a9ac0a5e44a34ad754a7f108f8d767b22612089654989c73706d2b8c3c5b3b7fa12a99e39bdd0822b0db5af81f2d47ecc642b7909ec3aacd9650f38285219b1f81152e54858fe52ee3046f483c8d960c09496d31dab4b91fddc1f75838132697c11e8e6299f28af3a1957962514f665205bae155876ab67a92608b3a7556eabdb3e28ecf7e8ccc8b5adc6d826603bfe78a4bae446c55f68c5ff2009cd70212a6aaba8d51ff9adf4a12084f02681048a3c1f77532fc7203caee92d23f856fff66420598dae01462302f9600daa8bdda7d68bc54fa674790882c8e8d5d1630d26e953c480d2b9efd60c49764a7fc109d9ceb78a484c84b6550e3c69b394db88c2c719a74b7c06c158d9dcfd254b369defa11bc6354ae362c728662294d4cb9f460cbb9aa7d65b230cee0c73e15526ec5ee01e4e0976529bdcadcc7f6bb465e11cf78f69a279a7b8dac9147b3ba421cedc8aab7e56043021cf75ab5b9468ac0b0dfa92cdc35217ac204dbc715428b92beeecf34280753f8c4449db1292ccdcb3d04b23747126407bd5998b4426571c86fa2005803dc31ff505dbc08714900c11fb81e6ac8bfc50af8a0a5a70f60bc269a67a67a76509c5cf2c46a6270bb6cf896186e11d3a3cc0a5056f55365f57c268e9a58de3a8fb7b1ca430769bd7972b6b77b1b7528bf62dc4154400bb2606b785a37cd2e0e511e9c19000090ead4187b9776ca2a32cc7c0ce8f9eb4a119ed1b5f5aaa92825b91444a69f3908dd1dd8395cf0fb672dda59376929b50fbe0785d33b06bef3893bb1ab6215d7159dce8bfec7d0fe37ecea30e915f28bd427c3cb8d5a48ab202879d5f26fa71c4a5fa1b6ce1dfb2e93eb7a65ad76967be570b5f73dbb77e0f1cd4992ec56a333731812ef22763e334f77453d3e3c2d4e5cca34c66cb1f2b9a8f37ed51a9e4ae112734d56f670fc864570fcaa188f5eafb405b6ed86dd14e352a35b46e0837365828199bd895d801f321918a088ef0c8d7bc8f83831b67cd4a9d40bc6ec30f4b2d86fad43eee4c199a7c18de60aef6a9f16f8407b7bfc045d248c5af500be2e2c959b1d871bd2ba97c01208db6804022c83fdf58452a592d16766ee6c8a8819d77bfc6c9d0d09aad746e7b667b9c486318274343f736cfe22c85d8b0b97876e9545c771780c69d9fdb389dcf90b59ee751bd4eafc33a10368f57d326cb26a5e6463f89276f9f6a3d6ea613ce7cec6247fdcc3d8a73e327632becb95028e6fc9627cffee03ccc5f73851ac7b8d7da31d58d0e763ae47996fdacb8eaa54533beea9ec03302aa66569472826a4c42be16ec5808df03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha172bd86c97e762248bef9919c8a9fd87a4eb647aaa7c08f1fab3352965308498957785463e483146339717e31a1d94246bd31fac52de686ca937d9c20d70d7c4a579de4268ba83399ce2d14788fb14d9af737d6bf486b25169a45e5aa2018b407515e64cd9f9fd0de9e65453ae6cb1e1743a0df31b07958fd2768ff1f1e66c291ff11867edf0b4ba64ad2fccdf040b3eaae695d32498174e55353bbf33ff6af2de5759b2d39e9591218f8a6e06bdb16085975acd32ceab118a3b2b54f9c2b78b340540bface0292c702727ea8dc6a4aed82efeefa5ae2efb729c002d2589a5bd54cf2c5bee9c25bbb2e67b5babb1c33b0af04ea3c13d06c190e8dc1647d7405e5006833a2065ee3d698e6a424d064a1c031dca715d137f864a5ca276fa2ec3e17fdef41a8a145c553738de9310d61120559ba714048d70465f4b95365066a3155657af19501fcc596e96c228fb5a46481ad33581f412aa20ab2de9e09eb124c20beb59040899e916bd5f8a849d6027b7416506726455747b29368d1b474f3166d8684464197167f561bd3bb78ff9f7a02b916e81f3f5b978dc17d25bab3960ed1c49bf32c750d3a98d54b0a7305eea0859eaaff89bdd7752b3faa3b5485c672a1dc3b8a067629a793972939eeb379a133cbf8f508d91c9f23001857cb8eaa3f031b6fb83dc40dd5fdd9bf7af6842687d973539d391ea206181c5f468432b892418af1416058ef858e94b89979159de5a4aa2116519d764b82a223f82728da219c1f34b9b2c3d5b6723f6cec00402b843f3a110a9d0f3c5500227602566c335037d7c45fbc93008a999f71af755bb04d38cf159822c8a56f6ce2d54db030f5269911f5889fa7cc579b06362ce14ce4f5913554d1ad22a9e5ca97d9c672a946339209d5b098a51226b8f4fba67412404e0e1c17c0318eac7a2e4fa428468b407abca0273ebfd4740c820408ff46a1167e25dd47e85542361e83604afd29e016bdd0ff5cc333d1d95e537d4a938d90682e6728f59168e9899aac27d7ac30ec4b0278c0ed63be3c26b3adc93fa35fa89688093aa986aba59de3eac4c56f261d8f0a7316c4bff44e02b45e0dee3d1d0813b82504087d210522c385da6b9438544b8c3ac5195b0b11b2da29fcc68622b8b67792109d383c1d957244b4d7a7c9fe96dc648c4877b76b02a2fdfd63498af989f0320d5599f95c0c25b05e72f553569d252c2912aa4c63f480a0d0a0cd513d5659a01aae1b788690d94512cb83473d1d312d8d261f6b67c279a2e415b45d3b8bf5d601b6b2c08a8c6beefc5cecc735846dfd1a9a6f6a1c7d0583713c867720794fac3dd3aec4e247c6fb4200361a714ee53d5fb2ea426e8ef033d185b178cd5fee6ee6f7e20021ca4f82959004d8d5b6ad2958215e8c50f0b08a4cd781cb77eb9634ee3a93afac97330a6c3259458be451043c510dcbd7be6ec58c52a62f45708383019c9dfdfe548079c0d24b5e058085fafd597683d00d8ebed694083d86171c7c5f94fd9e31071dd4c5ab89e53571dc33ea174d52d8dd77c02fe7237bd96718309660e3548838eff50b7058104a63510ac90438393917fdf61701f15d9a17d69c9553c31e2d188cf431b60ac60f937b258429efcd50429fc9a44d980f3c2dd6d55cb2e890b8e053e5e9445c7127d745e3fd640a7b0b869bc1f24e657003f6979b8a04b3f7dd7ca9d22d7a12dd0221647f095a3f9d8e25938ea98939a2c86c0eeaff071a59b86927e23ca13f14ab547a407539506ce0d34d75ed73ea5113164a2b4b1928009773294cba04074d7b3088ca0d2dfd73bb200184962464890129957797eaf459714e168a3488fdcc4c2601ae2ec167eb575e9088e1fbbcace3ca2476783788d790066d7a829a2ff82fc8b51b4eb79d8b6fa80eb3333bb970fe250e885881847039145de0930e62315c002096797889662d9ebad60b7a1d15a4d2b7617667e56b2e19311be47470c56cef25940015c5ea36ff684ceb8066cf2e025e7c0d79d80deaf9ff9f46ed0bb3e9355b68e5233b36a15c21379a1b99e39304c65c67687d8f50f4e49dc7fc4d94b3fb0bcedb0a40362df24a02d5a89e664a72e7e1e66260d619ca8f14f7832b8463c27da3f05e89f060c502c80872c7dbe7459bde863af098517b4ca2cef8abfae0a79aa905d5c2ff6eb2ec7a33a0188e434f44b378b995575926ab4a9b61403ef38754bb162364f53ea1b0dba5790f9ce350e65d934883fcbb9c3db54ee374623b7c2cf55c5d3e6ad348bb21305884f0f276a66f4e7915059e48e2e9346982ea2a3463a4eae9520abd0df5e8d0317acd0cf604191517786dd28012505fa4bd152dff6b983381b713ce263faf99f3f73bb2111d6d4eb3e011eda928be3daaee4c7c4e38a273073e0ef3a9cd123b9a62e83321d83b71b87447f1b6bb253548457ff1f64c8df249bd813f1dd32c30d09f5d41d85f557ce61ee6a8e2708f02a71316453b261f2ea0bbe31ae06e20deac0a1bdc89cfe0a4c827edbbde9cc29c509c308536d9c3b9d9d540a5e7248e1ac26b05fee7256df70ac50a1e63e8d68048fbc64e4b2c0f8b974f79d5189762fb51bca2cad64bf4594da5800e346bee2b1a4826b15a10b6fdb53c88bab79e55be8000510bf4523b7086f7a0f597a1000ca2fd949a45291cf9442152f740f54e6006845bf62c554994688be4843b6daf665847ce4adf49d1fc71ccb8087d912b9e104587b79046992a6374e93f10256de0d10c69c6b373bfe8e4461bb4b975324018433d4b8c3acee122f9f046abae6edbbe425e19c1ca0049010aac06f1010efcd10eddb4d9d5cdf0f69532606cb80c43ddfebee4aa45411f24e828d18404541ff9013b75ba6c041754f60ad8bfab2ea0db0fe9fe51b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he3511d700ee35b27a3a0013283cd421229a6bac7b960e8160972ef18c3bb1648c49c489a8b3969d5d55512d362f78a49c26f2500113388cd4d484fdb8abe2250ad4306c45b5c905026e054e48ede72fb07f0ff1cc4d5542a51a3708d04900d11971a170918a17c1adc8a594919b1241955b1fef357a89325c9c35d6804ba9b60525b14c3f1ee337b11069962b7849dea94b557041963c442b6f55e1c989884b1ded478e1c25b4b9174ea91e47646f05d5b430938cb40ddb01aeb3e8db5847c1f74764393e57a890056e617cc2b3186da44917f5688757f996ed1489a1e2154fac009f557bd172c40080d07019691771fbc810a578c909b276d0667e738b389900e46e69046873098b4ea6758c5869e4312097f541a08398a0e69f455da6ee6bd87e431639ba7a1b7608c57f5fb11701203980944d369230ab33560c454b3e321ae54379e9ac10ae59610c4efd40bc6273d3acb69132422ca8861c8304744d99b0b23b8f767952ea4dbacb5ded249e2968bf41089f9878c7c91bce9a69746898ac25f94b0ab7f04668b3d622a6e8fef3971a44af2cb169d6dec4eca1140be4ec58cc07e1f66814ecaa45b6038669af607e187420ed3595fc0099953c35463b86251dffa1a046d4f7260283929e013a68e5535864fc9745877cb8bb634f629dca9ccb5ac5cd810bd0e5112e8a117f7be9bbe2bcc9d65bf8d4283b12854eb2d0f18785ef6b880519bf65d85e6f35713e74079c309934ea8dece1d267d984f98e531c270a622c81f7a46308025a9847fc9fa417b71f1526dc1bf6cbf04c11e52e92bd92007cc315bc07c991d3e555056e33ae64ebd550af2be1b53bbf212a792b8202d6b03ee38a84eca65d258dcfb207c3f812e17f62855b969dc290cbaf149e85f35aaeecf89b1653e0e57cb95501ebae56539acfb542c55e18a6be89e67974864623552a386eb41c22aac0477ba902461585cfade8cddf210d7def5b7f915e43bc13aaa97e03920da61fc08fac498661f4003d0bfe82a2591e3706eb4e4bf6affce74733105f56625be3e9925154a2ed82f3b9388440f34e20310218328876cdaf4ef2da5b82d424103d6469a4199d9a8eb89c0b850ca66db0a5042d77af8f898857f25cc0b353dacbc4566b464f7b89212342e189f99a04da10c42aff69661104a16a0f2d20ac9e0bcfcbf8d76035c391eea9c1cd14653467a09ae39d334c60437e5086c4817dbd8f95fb91a1ddc407d7013e13f24caf938e0586909b537a003a6dafea8dc5aa986f00e026dd7bdf8c699de4211782367b88026a0de34edc3fd900139b9fc8cf49db253624cf4e5d96d770202f7ff5bc6a617f863c5c563de2cb595270b7dfe2ed6b2477e2519b4057bd113c5878621fec21300e2e3d2ca9d97d49f0fccc6468ea2b0d6a7a223b1dffcdb55a8b4d3112f154cbf90cc31433075fe15f103acc400677a48f754e535cda5fcae54faf347f5abea6fc58c40d720cf1584ccfe919ed9f875243ca619168b8231e303f467cb7eb7781d6cd05d80000463061a12148cb651b1f3e898f37646231ec236f53f6656d05ecd892d7f5001928ba039cf857f494b572c83db151a9cbd89a7b90bd31f876c6043888067968a5184b84a9a09c5d6440b9ad169072c44563399cbe8f5acfb88ef466317f09f3ed72d969ed48ad6e18b8430907fa16d13ac05f2709455b0a41fdecafd3351f89c35c0824150762d767ca880a499b33bf0e4d461d7f13f24278326916513265aad8cf0b882896d02ddbfe400aa44c2f09b24a65f1b7ad76d384c3cfa4cd739a4da0fa0c7124fdc0dfe583457f6520f16195d824cc8e55c2a436617cfaa3fa4b09a7281e25d0fbf32c53a97e702d3aee2648fe7c722e81bc591213be468b1ae4158a97ad38f96d8c5d31970d2b4d501bc9b80b2ec8855ab77474f9f92f34f6b51be44e99a278d3a0a12c74ba77249b2ff7f8e11dfbcacc378fac6ccf54bd1018f2e137c0b7ff067841f4b130ee8cd8c7a8addf0bac6dab0bda40dd624be16ac79116f739fb2bd14a5613a4e2b440611d13d93d6ab486adb88394b8f011b1274dee10165ab91593fa7c9b826e72f264babea9e96e5da9ab43386e0dadaaf29b7f97fa791994d7574310a303e2a61884a8860a7e9dd976aa27dd9696be48af79acc8eaeff227f59bd044a0ca8d5e5721138ea67c301efb81b1b3d41cfe3b2f0e1bd58d01cca55058ec040595e011d7b50c4497483a47c92cdd8e8805c7b28bfac210e8477f7a41a6c739b5caf12dff2f768625e5e2931e6134309968f47a1634dd4ad74b22705e98c5ddcdac072f7b22f65edd5e09b59aadb1c4dbf8d0897c3eeb1afed72c714015909d8cd8c3d81a94c436f57cb14f0e5d4786649b79425bd2a79784aa14e52da616aa5fffef7f1ac57386c4304452f05f95c28c11ffe10459fdd3d2f16906becb0d4a520c0e9e6bb627fd8327bab37389ed305085221e062411400c8e8bab7c1b85bc35ac4165fe4ff75bdcf4252070e4d706db0348937776a46663a956bbb6528470fc466616acf0c7deaabe8f5a78a478abfe6b29ec12fc6f369683d795bbb53ee2d1b569495bd05eafe4904416690bfb81a6544b56694694c3c9dd77a079a2699c2c9f5565daee5e2250754816cf5b1139347ada478f5abaf210c7328f4bec66b13f4228d689aa0bce13a23412de10be7ead2f7115b715779ccbba4a0cfaaa75992543e2b4fbaa4e6883bb98f8466b59d3f5cc7bb1d46f029900a2b14bf90577705d91f30831c8fb921c6badab30f01c0d54852d13ef36bd4602285a35d7595098aa30bc245b6ece22525d4ce83a5f0f1d58b48b36249b786a59805336ea12e3092f0b23f1c02adcb76b504afaf7cac465b29e55c0c841a3c35ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h638f4929e2567b3402029c75e416e0fc4db64e7cfc46c4dff234f4270ee064ae241ea0c4193450942a6c924ae5f48a57b7169e82b936037340ec299a78b6654acdb9a46992549ce2d06fb56a41af0653207f711f30cf98cc4045c2d6d08b641fc1e6e32d0cb2f5fc70d569c3c4e583b2c1d7a062670344fefaf4213faad511d912f473c9c0d1c1f043f0c48cc4dfa9e362bc9094f18591b99c309ae231df34302a7f104676f9ec3ce6384c0743e298c791eabc814d4a670e4499b62ce046993ddd3c60c3e7178705d663252eabc2f88dcd44725d707ff14d4fcd360f4141415eee11ed4bf33f4ab463ff830e43b35ec0e7be962c5cc32811ed47191b5799a12837a66ba71964b970f3370d85c5aa7b8bf01b7c75befd7775416cc539ff0dade5a031ec56fddc6108deb1194a12491f6c0603956ee2ac9ffb2dc87dfdd31d7d86cfdbd10d64ccfff1276ff28b547b3d2dd7f20952385e307e4385821ad9ee149d41f691c1851bf785444670502ffe7e50222cc4d21828b02a246110750ff408acd8040cee7b6da5609bc80988f69f61e25fadb46bf89049da96d43065ea2cb956d196a83e2f47a0bbe18d6b1e05a0544caf60fa5f9d943b36850f099d414ee47b1e0515a93043d13bd688d1054118e8096ebd481fe03ca51da171c83e9124b79d269c55b63aca35b2a98e7c1a694724cf19233b51bf54a048af0fc45d4db9156b3197b0c7d9a792e8a7c9569cdccc9e97625aa4d3837bb28462ebf7371451daa93675c92be8a1d7afb3f08bc7e0a23ceb10eb21f84441e1e9e504a8e6338442afc8d2e50efa4d1ab8a909e183b972200a77608a276cce316fbb964f49d18944881e65a6cd9838ec1b0298d1af623b50737acf8ae84746e2f44dcffccdbe9e2090757c44a57d281b9072a8a8ee0658274b65de2c743ed7c7168d17dd7a3d9cd77a425f80f02cc4dd31dbf600f7dd5f8adb4af7f28947a16edf5ca3886a7296f683a9700567b401959d7ec66681ad24463beedcc17d580f8abfc809d3d4e3b80d92c7ff8a61e914dcb33c97f5b0e87c1bddaa8dc902383d144dd9f0032a77bd35e19df9b074ec0f45823091c67131bb40f93f209599162e38512608c8668529a729c2840ef9cebcc52fd06ab7ea9e37486d4ba33fc36cfcd2338fc3224800c517603f9270006e3071ddb40ad0d89083be33b40f9ae50945781586f4fa17dfd9fa7299af50efbfb5bcba386e1144969c0d131fe91a1dfaedd501c11356bfef52c1fb81df6b3e450035423eef36b4857a9106f881f7bc15d982bcd5b5a6a9af6ddbd2da9522aefbce7f58650043c3a391a38564d702f4e60812ab530177a6a49328180626a8845d8b6fc1364740e95857294ed0a64277b593d182de425190dd6e075b2b509320aadbfe09f47b87d8f15c1362e923a23396b836873e6029731f2a161031a7bc65592725959a456b269f50a6d79327af926bce6208d880406192e3f1433547b2dea0cee63e7d65708dbeb02e422136156449ad1bf1ad016e4614a3d50738a746ceb8a3dfbcbcd6dfee8a1e84d39e925222e02f102f554e30078add87bb08a2808b0554b333dda8abd8689728e8e344a62abb21cce7fdc508282fd79658a237d6c7167b41f0f6960838a96ee97c00069adef3b381c12a89f929bf53b3ec932aee9564b821d347691db866063ba6dab06072aba20d584c383a1539533c26b86c29470d217d2d84b2a2dd549543f4307b45615fed416465a042b79cd0016df6d996b85aa8b8b598a4f0b2cc9ea27aca894bbbbd821de10e7e91c08a3d0344be05d5ffc9c3ee5e75789d1a09a134f1f80673e9c3a1ae20d2ff9b82408fd77ae22da3e980e5c4f32942dfc671de54b1c4c5f37fa7cd684db0a31deb697e793ecfbd99f087e09b7b204c51f7c9646d3e39a4912c5c8f08c2963c63c16bee9ab5bac83d74d6d02b2c069342a87d4a16e8806018b2ed377ae1f44e0bd2603363303c84b2dfb359a11317aaa3573527ae365aa1189388df14a7f60411f8ecdc032828ecdc6aecb27c8097ac903a9b026cee86e024a4f4cacaf587e0c32b6e4f3e5a21a557186a0ba91c59b554c217454bdac1e07648124809905d5f592ac798763324cb3453dfe0e2b5c1d4f8a2bb22c09e7eaf7143559a30293fbca954b23cf1e34d9922290b1adef7aff2e629ca0fc7d23fe9599218cfa7de697239b8e3a6d6986a1c079230ef9be6bb326f5c10f9abdf8c27ebaabf7d7d869377285b6245b7ad4b75a89e0a05ddbb21d9734559c5d5028ac06bbe93b50507eaeb90924ac0c07dfbacc5d966bc5a7e50365ac09428563ef078b2d91dd8fb7bf37de44b307e1e8ec8ece8422aa97f08c58ee85de10eca49241ed62ae244967c964d547641f1147863de16f1e5b7c4f4e16e6fd4a62c7901faea4bfe0de20352616b0905d78a006b5d053ac8a0da7cf1cb14e69f62c8cbab2b9b1304f7ae408ec7e33b867650f3581b7055d481ad927a2a55f4274f4416fa08889d5a25cf801e4cca737d104d17a872c468193df155028fac662c26aab48eb924df9789f14e2bfdbfe0ea0762847450db5282489aea15faa7c9a0548463bfc07287ff95b0fc93f30f88c0f4336bd4defbd94fd8209dc3451971760fe8fac8e5551f87303918c6c77af0193845da811064fcdee3901e9e3bcd272b8d926fd61366a457b6c58193dadd5a02150882b63b3bd8d4b49fc52cb85ba511e3512031abbf6aa86b6ebfb5a5b0aa4e342ec596213b44c6010f341abe615695bee59939343e5e6e4ce7aca4e7a5fe995b6ee93a8a77e60c5a4f351274d84862e1a3ec411665500ac1f3e4af5e0a27791c0c31af74996a56b0676fb884248d4fa064ff77bfff2006d300aca9265887a6aabdf8a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf1f546b6e55fb6416a14342a814cc57fb6d441d284b763f9e04206a6c822bd0c5cda5e6dcd43b8da1070b6b18576e7e0e1fe678870572386a9573d0de1af1157fdae4b404d7d14d763e6e746f8d3194500b80e2afd45cb393361f90c100829eb4b9f3e1f585ca8f1dca33490d0550e4b64e04c51ef435fc707754396a6a99078df33241a2efa28dd674adc72ab38f8be1a1479e33b5b6a998415abc80831df59e53cee99eddea442489a21faaa1e9c47afb5400c353cbf32a3cc7457607e4055292f7a0512e5e192730ce2dd00d040111f501a1b48cfd0026541bda7430480a27096248d6843622a29bcbd28361cdbdc7e480f938c7ea7ef7a4275a4d87e81fdcf89f41028266f695d1f433c39bdceec09fc19021fe8fd4f7da1998131b9b82719820ed4cf0aaeb2b8084cf9359e5771864f3ea81207f992d8f541d45d73a281134e0d5623e86ea53df77889e06887d13dfc67f395e012b79c2dbaa31a12fa7d4343ee90f456b36159ef2efe614e5fc52dde1a97e121dea7d9b10a699ece89c3e1d3979a1cb03b879df55404e456d6d5436eacc694b121d301176c6f076c89cfb098a067971ad6d7ce55b7e747f9e9a52bab73b3a2b600a69980337a94a13a64c1adc23be2b7efec92dab7ce42990cce12240c5e28aa7375fddcdb43fcc2adcc8e3421de0fbdb76c1aac066f7e4812f888118193472db2fb9441f87497e6f36603e9606f0e38a76abf2fb8320e4f01f874d2d6da5a28e22263e9e3e343682e64cb0e7c67262f87e8541ab22db09e8dcde4b538d46c18f4df60122b794b40756e5b3c229f1c324dd9f71f5315d3c6c840c78fd2458f266bd8e88c4aa6100a6ea2e0732b30a7ff5b69aaf644abee5f16ce069b37304f982f1a18bb1b0f62356801225198a09d158ce89dfddb45db04d9599dd51e1b9fc6361b3437313ca73357a8a93d98263831f2f715035f8787087dac6a7bd118f4601a8184549769d3082ae7b55ba47a0097ce5e4af4dbe8b0a662bf8bb9e2fe7786e4256f1e8f1dcbfad7ab32ae9ee493dac839db10926dd79da9489e1d06f34208913f74f85138ee1a30edceb0f7380269282d319a2b927487f30afe195d8058a9d976c6a7926e10a87174ba157bbd91e1f6634c04c6bd5babca2c485b3cf6aff95a3f68473f07032807db00bce3f64695f7ac0f1a608bd15adf192ef701deaeb6556c294f388391041bf56a6cf48399c28261d740dc3915714cece2c0119ce8a161767ce17899a0c2a553c729eac6c7ef1ed2e5db2ddea685f28535d7253ea11687fe0318b6f611c913863450022788a70c0ee4cd6977f0854882825342bd1138bcaba199b35b5322890a339c5cf2c950dfc05d023cf283e6c69d932f544823ff0191c980c711f10fd47081af3c98a96865a5b0ce093e44798b60206b146256d4d9d633c954e6446c7b2fc7f2474a29f0aa566d0293e718f014f910fcc4b29e481066ca465a34df1d2848fc2549edae7762262bd1d78fecc1607978edd4b28e1a40b9332dfa41a5469f3d3009d208445fb35eaa7c62070a983dfe6f7594adca4349ba19a7a5e8a2257e6434591c406e76c52b0abd7e5da9f2c00ba1a2191c9762636c59d17e6673e4c234f5ddd308681b596140e9758334ad80b13101c0fa4b6ee8b44525dd8d1c096ce743b35529611a06038829751d635c40415fd3cd3a8ebf2c52faceff176a0428f945418c2224a3c751b3b0d1d9b16cbfbca9e20ce93cfc2687244adc90fa9b8640b25d6d9a4e83f760e2fbae2a86d9134dc42591c58734c72df587f4feaf7707c54c983a3952bad6fe0f8b8814838663d3e5c6fa32e39f0d6c4448ffba7ba5a899190eeb7516561e85c1d51443f8376250b5628cc2b1b4e7148fc1b28976d4cbcaf3cf2da23917cc6ce80e695be4d864dbe7626f07c720a21da85124fd4a1f325e072ce1f1639b7d1c5d7e36c6e16857a2d42b59cdcf294c828dc0934647744a82fddf21b7488012e408f8a9755c309faa79f47707518fb65c15ef66c8c66f00c9fd42f5dc9f6ff26ddc6ace57d2209c656b8f59c9903267944ab9819265cc2120943e65459a75e51d5d93c447b9fbc4d2d6c4d640e16d8f8f317fc9493ad2060974f6756d8ee1e25030134619e4a4f42cefcd2a115f96e7f4830c9e95b4910c119126b48b2db2709937959d24008873157c32a03f35c299b0514fb348edf5bbf7df6c601beb0888f961302e738c8003aa3de9b54ec39a23b0ea54f301d1f99d21d68a9a1dfab0db6d6b6e09607ba5782972ff5552328aff1b48dd325fc85fad8906d0f023c84d2b2f9a907427ceb218e61edd29640a62f6de8b716a04a4e396fd40457c362a5a8d36b9e08f82c0f284e5729364e3ef369fde6314709c44cc6e8dffdf4f834ac2bd4157b41b75da2dced50c95f6520d0342fbfe8091a980556178599c8f01b70dd019c3492ec3997eb969b1e30a54fdf869c53540018834f583357742fc1d3aee629faeceeb63823ba1017fb6f959f2ab953b8143ab0506a427ce303297f8686558568149606e6d90084916d8636fcb7ad6b96e3f9d2a614db0a31378285f75f995acffbb2ae3e51f04d399268c80d5d01d53254c83f5708b9e8d33f4090c13447e70bd8fae3ef28cb2df3d49c711701714c871496d94c37f1e42a70e599ba086768dfad469cebbbb1861bec68cc82b9470802b160f245cb905fe3719387b7d2bd599744f884dacc1ed6646e0a67f87de7aa828bf71ecbe5f478d6a3f7ff7943db7fba17371d2e7920037258e3672f4b1d3ee28104aab82509bb63ee3db6589d05b8ad6cd35f1319b8df158ed568d9776516b9ab35bac0713bd1ea27f0814f7d4f80930540607265970328f03b60e99ac3153e19f99f76400b9f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hae499f9550422a6732776eeda66c3f4486d60a2243ea118d4bd9b6f07501a72fdf7c74cb3665e431a944bf88e5bd8b7e8a5a02ee59f013f82e2664e3d499ef6602a32907a2acc63eb986cef492fa896fdd44689cdd07d1f4a99f71895a07a50b4a4b38ee417b216ec54087211b7f11de81dde808c476bf17b3d0edce9de33dcee05030cbb40717c32d5d2be17bf50a14cd9718755f3f4b8acb4da8606d737ccd962ac1fb8184091a70703e5cd5629212bad83bfeac102c7c5652f5487489e77de996183cb6f5790acdfed8e129de47a93c22ba77db43b3e2d1a3fb0ee7139e85e70a939021564bdb2ad1f54412f7999895ba9fb9f4e625eb9f31e7cc32422d64376ffed8a519a1f624415dab81b34f7c485068a1003ded1469f147cff91c8410f6b26805233f31fc779a0918a998ba43c2aad3dc44fdb97b25226d21c647789135d7f54e151aa19ad0a810a5af4613514e43b5451b8edae2549e18ec8ef96143fd36d0c144901f0c494171f819178a6c331f112e3426600e9e1b56397b759c2872eaf0dad7277384902bdee81d2e99cff65ac5d896422047d2702de0b06c497cf3cb1cf5df9a4df0eeaa91ebb3b3a1f9351b811877849bcd312fee424a4e12c08e6b5f958d6314c0837a7cedb4abcd7a3c4a9e8f96cc293dcb95a823ab04e29448ebe472ba408dd105aff3536287f1ed22eae92bc44f6e635e9086e4e2b5385a3e8b60d92707d1eecd13d07957ebda65c34a9494881836e559e966e36f60f5f8eb9c12132db2f321ffe95750165a5bd0c4df20dc6d8fe698622c5d5d40c2249a86c79b944e51fc40c584f8a1cde29f8e393495c52f1bc640174f4687054498f7772de705210e3706e3da5cddff4f03e866b3a5d2ac79795d7378030bb942313c33e092bd7333a2711d8d30b0fb1cde39fdcb0ebd1fd436ab9b3aafc08710e844900282754ac7b41418cf11869c012cec4f5d01f30a9f6decd6c021589a92d0e2eca4ffd3e3391e059bcd2dca1f6ded47783fcb9142d36b1318de8d558760b0b337e6a8c3014fdbe005b67c780af29817c41373c869badf430fa65cbcfa2dbee12efc89cf712556de092d1234a1aa3aae387d6f26774f7d7451b85a2fa835d676b92c223036ce411c3f686ed9d0c71b845acc5fe7344905627ec56d271debbe53385581b1f2d057df4f42ab4e03fd4ad8a9c588415135b5ae4f1f0888791f8a7e51b83ba3a1716a0470f6f867126d61b1da16874763ce85c0a74561010c3cef42d73a0f5764219ca64c8c347403cdfaf9ce860639419d9f3fd6086df40c88e84092336686a23348681793f6e41430ec4b07919c32db9d439eff23575866a2ddfb5a964d14946bde7b582351d025b09771071d54945ed89760bf683c307e57d7e4c6f06efc57aa873ac28404362f066d385227c22fa464913ac092d8d478bf384c967656abb9a633efb566c10a4953ab3c6cca7faf43cf3e6dc0ccc1b976f6b544ec4a154fbfdcf85e7c6e78c22b55d7a640232423cf57044a1d703cdde1741f9e903e14d2f175b703c77ae8ff8259e41f3351146c306cf7d666c81db3bfa2680ad9c7a08f6e0a11d3c008e736b38f34e999c31685c2e8fb777626b7586a5fc9aa93aedec7a758b8dc19c1a541d9f756094f86bd030a4fdbbe9c1e93eabd929172de81d870fc1986bd645caea2a57ed752626726401ca3be78b2aedb29f02a856802efba210d21aa9b9046608f4cf8cc860acddb1a8b629454e11d995c5aac0bcd7a2f1d5f75c3a038640d3c196fac74447b917fe3225f8da3148b44c6c987fd1f1438b7ea411b1bc02226b795479bffc44c38e7c2b461f25698dbbebff8c153d12293dc5d254e7897df12a8ca24d0845bad2f238792a2fde5a1e6d324a8a18ac2f68da61e3e44b00e78de3302b0b47efb186fdabb6e4a3e6e9059eedb4917218c4b226f9dfa3bd5e478d61834454bb0029a99731d14464939e80f6d9c2302853a3175e1bc10310c18c7bda163ce78fc3bb544cb1f7d47246ff6db34aa1035d91274cdb6ab1986ce79835c13c087e7dabccbdb12625d4f380978913a5d26216ba597dc08b32e9fdc4ddf5588c7d83c2520a670fe52b890f13f78e53f13e2e93be813dd041a33b7fbf6ee5dc4cb8cb5e4f1057c2554227e3b8f998af244a7a2d2a20a84584f1c1cfdd6bb1db8bddca9a7e30fa62a2b6f6416c64b8b1378c744d51b86018e3bd4ae279dceeb0f2f65592ea397e4316a42390f59036a9ca44e6d8346e116cabca4947877818ed87fcf1a47b501d8589b1cd313bbed3edce919e0f833addbf29cc41870b99fa3273d1d77750510efe6734cde9d80b3ec88324cd54afbf0ec2594441b47fd3c42808de61ab224c6237e2390e3a67eaf5de26f9a8254433e2faa56b172a05c23ea59149fc121ca98508f48404fb0d68d911bf86924bd574cde4bb332594a2fa7ee0eeb9bdedd157aede7dcc559f887761c228855df0f3c6522d5b2d41c3f29f43073305101b1909b8fa3833811040c29c026d25926ed59c25a36cb5628691769c0efc12be6849cd12ee71a0effd8007379fac9441d593309cafa9c06d3b2245315e30d4c31ce329398c02eca79bd03388efc503b1d12d4a798c22ae85a206c8bb3dc527c8cc44020017e4790e909cb275673e38f8c869ca793c4e1e6cc4264e2f2d95b89645549b9c6a5c15231b1141574e4ffa626278065e83926c58d30866d95ad83960fd22b6381f8c661a1c49eb16114f048742298fd2e18cae42d307021550e46eb9766fa621ac631c08377d1d325714e0aadb6ce892e1216c1eefb8b2984a4a3a948856db9b78da0aea65f204da86210f39bfc7e72f26663772f2a93afd31676cd9412d658a0fcbc969ea973b5e095e61891d547;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h564da2bdf0dbd44a39ac69a4bdd9e9318dd459491182350d927930472b877c612a257fb874f4f590e390203d56925f46c4cf6011035d4f95a7cf661f97ed53f9b903c323ac641f6fe96738ccafbbd4676ec87f6ce00c63362bfaeb261eaab1be7d25d087f4393fbda4c46f0f6bd1a26ec0171d03f512a1b9b72fb8f27f8e5fe934714168080f3997999c586d1791840c87e61254994b6975226d41d5ca49ddc9ae8e012b5ca6cd666af55c7156232eca327255807eb99b965d9bd103ab6683e6cd476dc9a9899d404cc9d6688c41c7c07cb8dd51f9e3b291bbb40238e6869d93a21e29f21a79fbb296ea7b584440e619c5622527f0886b7b4abb265aea279bc4519ceae3d6d099e6c940c14b433456b6fdfc239833885a54f14b99bb62b55dd78748f9b6e808c41f23bdf42310ab27b2de5ed3de711f3c7f2843a2e758d5d4dc3fae6d75836e5bc597b7ff0b3dd6eb0ff92777e35d1d06a91407f2bb442a73c0b51152d8d47da76b5bc03f3ff87a51cf5a7c00482d071c7a78ea700454725bb8a0d74b858897fcafe7a5a14668384dac7de93cc5ec18838be99e58e2a6750e9177cbdd20c6e1688e374030c8d2eb6f5a9e6647a75a649f26986cb86e2f91c8ffcb97efc141779e5dc36a191bf9bdad992235c627ecadd6e9ec494a4f16912cd9204513dd1db35eab4aa5777a232ea7452672b0e65f9da2b19b1e702fceec478d709e90122b53d559d71318597af25762fdcba9ac5ba97b702ee56ee2db54760292f1a51c68c9cbceb8effe1b0f846f2939ec379ac55165d10613a568531913556dfcc140a656023c4771785323b90ab55228ca93a855a205288cac90354b47b0692237c7dfb18d4e928578efdec1d90fc018859cc3b0e77e24ee8336c599319ec4ee3e5a71e6f193933bcc1f1ecaec57a17a5a0491fee268b350996ebe9e8f6820150e31e6bd467c5ca1cf1ac33e823b902f7bb6e2992b5f3ff2d17859524ef269240faf32d290989b3ffb65056680ea01fb14c0a7ae2ed94842f9ec03886684037d3375498f5730e50cd7f33fc84470d846233f83223fd3d2582afd810c258913c4912de58a26182749334dfbb5e2ab353abf4d972e9ea2cd652304cc4fc425edc0c7b98e6015b50cdfdda7f568e8696099e55fd853953aa73d3f2827bf287043ebb10628bdd3b1c3ba3c66ee23c407d40989649946412f02f150d9ea348a47e8e65ef7e5e75a9cee8633f9948afe2dd3d6f84b22f67f247632b3d004c600819bbcb4e87b084c60a301b17c3b7e8440314454b6e6bf7cc639d752bb70023bcc38f20c30071548145a8e894ddcb08d1a5c985f71b76dfa46792af6086941e64aaaf4315190452e015c1d6a48913fe02bcdbfa4b1a1e101027bde4387b2ad4bc2b432bf7ae7af9ddeba8065eb5e695dc03ee79bfe9b4560399da83ee0ab13e0c4de2e03213638162d1be291ed0d6c014ea1a1f63f82746857980005aa7d664d6dec7afa4cc11bf20f2b755182f37b5370ee15a6296ef97c1b413905cb731af5abb604ca520b8edc0a756212704fa638626c8da97aa1d1068cc9a31188de04c799fcd22fab81035859f8efd7842a33c34f404db38a7ae94acf6d908530f3e5e9255406bf3c472876720e3a799e8923b0100dea9fb75e89527567d4278aad1c259e930a90ab5fa18b8859131cefbde762661c47afb982b51f73110f1f346d4b198325187628ab1144933d3f98771cef8f1be67afd918641ccc46cc0eefb06cc5558ce4ae111daf8f7dea33f1c85608f4e7f44f7d5595959078efef4bc4415e1ef4274f8f37f023bb748b8319e05f1039335f59536e2bd8beb3436b5bc9223608d0178762f3534803065accba0027251cb979438bdaee1853a5c02d1b4e4c7cbdee61a1ccfda09bc28db2058a5dc353a74e4dc846d423dcbc0d91308a893ddb2a14066dd1d335f571a08bf1a1453c71da6354eeb55fc8af26e30195757c6d4bf14fbda97fae6cacbc60cba2f3fb6b3c58c1a1d3ed3109641f4ca2e2d97b4a1da41de072ea39a016ff959a32eb468f3c74ad04dd8757dd246dbe61bc76dfb2a22e56c35d206d5216cfe6542309fff0ab84b9dd7f60154432c9d5f8506ca931a7c3d93fe3f401e61f7131d3cdd92402a62a728724d09c37ec94399737f7091ded1108a1a08c249eaf1798ba894fea022ad3acf6361bf7951d4fa49b02b9c16e301bf98a09ca68c54d7f79142656a5312499e89ff066e6742e68635d21cd74720d1c85cd79d8f69b134c088d974bd698c9094f7878a35fe8442eec3013860a0a01345e1b538d88ef01051faba07da11c3a77a57a5329bbdcf3913f1b9c4208d9f3e3c5409b68130332e00af8aee76cf92c783e1737c3bd98af527e19dbb5c4849ecaa33e0a6df9c3c7480da8ea9ee485cfbaaf8d242ac6576ea589d98990693f94479abc49cda57aac9ea36a5c2576cd18a4e8d52d3a8f3d749b69be05e5c311c29efb34406c6f8e2e4f7dd95c1f86bebdea4fd31c93996db9c42836f84f34a75e4ecf859ef984e0e84dda14da5c5259491f4622f4936a901f6956d87cdbf93b76bbd2940cd4e67a1a68d1e72c2d0ac52c0cd2ee858ffdc476b0bee9197d977fd21e05df1378b05d18329d10beadf6576847f3d74dbca43a171f94a52d96e8b4d273a068258e046969693bf0423d3c22b4d9024c87ad2eef4a2c1434f2a4502ba764f7212f3dd2d3ae79ba4d05db08fc9bb3f02814cd1afb73dd0b9a15f90f547f726ac2e053649cdb1874edb539370bc2e163e3dbdbb21aabb64c91a222230ffb4550422b61840b039c6a6ecb513941d1b3508adec6e3e01864441dd63c527f3b749f51abc6ff39d93646f2c62ac80c09de1bc5ef5b3ac7334420aa37cc19694a3253;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6e626b1280bc18412910d0b41fe050a0ea6a132eb2a2f95d46dce74c7d7c3f754740cfe506355a577827f6465578d94785ab3727785ee88dfbecdfb6efa72db11eca515ece3060dc923ab5362380d3d307dae31f524b4e1f7ced95f350263863ad58fd9f29cf8024e75a5022be81ddfea6553eccbccc955a5090a2abd652303822644b331da9756d277e5acf4b3c63a79c321781116e2aa2a506a297e9814eb03a3aa9d57b37b654dac6941299fffe0c2bf545f1da5228bbdbd9d5846c2ee19ef899c4410a0c43521290c8090b6009f6ce38aa7ac1bed7a170f1a53dcb466a844e04b7dc00fff7a1ac29cbfe9a1768388df1aca87059be4558ea2cbe94d8724ebf2b4e46b39cbfd9ec205edf1b318f63e462f4ca95ce67a8c4a7289ee8d9d59defcf0c09351e56fcbecded29fc79a0fc3b2fd707765f7ec7bb9d3c6a265662cb4120393d12601a0b3cab0888eef7db7c8330adb3f5275d14e3cf7293c305ab4b2f92e283e2cdc43e26c30c7e9eb04723e081c03ddc513498e150de5712e9dd6f5ea8cb6d0f675a56e2a1c808c756911e5013a363b783d3a7d2e13f022e2aa76f1a2ff9d2b6eb138e53dc738a49719bb7932e54790c75e09828eab920852dd20fedd2a346e67325b8856de1b844cbe81672ccf24468140a327a9b2dd03ee190e40e81aaa56d648a08a5495735be889ed4e08e442b43b5af39a104f372680f27ccef94f86303a6e947ac37ab976e655cb2d0ba7df06f44c9db37dc7a28d76fc37b758897bb6a19865a94a7628f323a9392aaa250dca776e14ddb3cd129e8c2d027d8eca9b14af2a9998ca258666e313358d6ced876b0559db974e69ecd8b6217b5065e06a3625a60268886f75139bcc1a9203e3b29744becd254e3b632d5dbe34a59c145e9313845a1ab8c8733761dfb5d0a3601b5184bb9df899951a0a5ee6f3f00fce10690dd3708006d64cf1ac18a63a80ec272be2331ba8aa2f6ec08f5d860395e578c6364de9dd72470a7bbba314c593723eeeecfafaacb713d13a4473f6a3a373d82513993b6b5812d00aebfac7e6631c9bb9af546269ce3579f3db2b6966f7389fd97d5385cca0c871a07040b3f162dd6f91018b4baac677d92f102c8dbe47c5adbcae394d5cefc431654578d94605d88af593378aecb0be228ad9a82e0e2967b3d2de444a7e5c89897ad3541df3a48b49ce14219ce942bbe65f5ac1335a4059b6638b27190185c22cdcaad30e217306701da3f3c2bbd6e3051e7959b81d23a945e79e73f41b853479b46bde2d62dacfff4da6dcd1d43f5a27094d221d3c8eea1863f640dbe5f34d23258318b9483bc0df2c1babe6b49f4b4727f591ff50b7fa7f4fb806e5eb6bbf168e38398396274927aa4f4ad354a1e0e04efc5f23bd91bef2cdc4f9b6504e007e4aee888ab581183ef420b780b7a5d54af73cd50e762cd5063af91f9576af9d6e1ff452dd02782392113f679dba2c130ed84b3fe058b65bc340192394ec99b95ce4cedf1ada45f3d812e65a263c5e3e3ba7a71b3f9089ad7bb03c3a09046f754a5498021eae0cc059be6a6845445894b4bb9883c1be5d5051c0a04f26d6d3e4fb10e37575cfc7437071a2be3b8f0394392d23db7332e38b8be5d47a3911df905cba698647021df32b60e2cbc40b6d1dc470f552db9d2012227eb22899061c8e8605f508c5aa4427fde9a7fbaef2cdb578ea824da3b73376cf67f86548aafb35dc8c75ba9b3da59506828762b3594013373626d4de406f0ca11c875e3d702102b916d9e2c3f01eca417e752177c1ffee7edc58166d2427b5376983c96eb37891c4654d9d41f1ae6b46167867a7b69dcc4ba73877ae34dd22202fc70739d70530600ab7395c15baaa134b0179dc0fe7b47216905f62dc1f1f0c9e2e852a5ae1b14ffe4f401a0158fd0ac0eed50b1e1d30b2c2746034c356501b87cfd2b5aa163baad6400f23929ff9f255f68a9bf964d5c6a9bd98ffc88aebcb4437832c209835db9b497e0b4a43c79c3990d835ce3361d57b64d8e99b7ae6c1ed091c8ae816ba7dfc20b7fc5aad29cb270fbbeb5f36b6455cb2b45d4b626f32a2b8d2ea60d38890b0172237592a674a9cd8382ceb1f8d0a94ea641e79d2b202510f18d20d198ec1e72f1dfa04a4bc0c647ccead6415420d286778b284c0983caf07f8be81fbd6bcf63fb19965dd82f364643f84ae3a7cbc40655ce93ef596a5d41714ff7507a7b1263d72cd32a4f2473a97b46730b366cb2d355e3a118cfe2315abfb3a9ba5fcff5ec34194bcbdae4fcb43447d2133521216d84b2cf694e7bd385a5c72c2c75d34e201af3ffbc4fd394ae69738202684166683ac06f218b01e327865c23addd4e6bf21af98db9f5cd99a16c2ed827d12f9a0fe4519a00238e96b7b69122c3d929627cce4626e1f0148efd32a3f98ac72091f2ec802c1e43565b31d5653fdc9655850f33c0c98139744f0c8feae8446b4c43e9b7d62cf4b04cd38667359b29990a68f95da9f6c5d77c03c808fa9bae02d59014c1e47cce35976fc5645ce1007a0cebc950266b724c94ae1100e98f2bdbecf8ed103baea0c7bf986abf0df230684b54475aab67b1675668833f24523e7c9514b0b0e1d6f60eaea579b9be9ed45d37711d25d9f94542d7f87ca2b6841b1f66fb3f648fb7eb4c1b56d288eb036423746f64b9a22a792af4c18b375b7006a1d2ece9a63d1d0765b7ce7513c17d230089f5df27ef8a4bb863b824fe9f790e01950432258818df2241a059619283a5b7fb0a2ce9547ab06cbfc8d091a58efbcd17e5ceffa785ada6e961e0a195109e00c1470abb6eec299fc10088a4f37cfca4e6e0ddd5c3b14a9f2ca7108ef4b08ba1bb16a56a5ecbc2f1ef78b89b5a5ae749c97eb859374e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he3c2f72ce0027c4a1f7fe9c274f4db8be85d6a010e984fb62dafaf62e5b368e110cd6e1552c867ceee4144b9d19716c202512d47b2143f17f71ddf086310f7c0770c54f293bf1e938d7f8fda9c6ced777a96278649cabe55d963a9b1fd9f7688863f628f63652f619f400bbe3e1dd238463ce654f21849385d2a90ef047c015241aecf5746f1b74bb4e058abaadba56e1631e5c9cda6a45aceb97e3813d99cc41ae98faafe372df51c5794c24143cd2fc66ab2cad9783aa7d6ff9f9b95134d8bfee0c9fff39fba8d0810998941ea8dc76db666f52ef4fbb2558fd43dca46639296ea453a263c8882eb199abb7b41f621647cb64e1cc77709e54238f75c41f04874ba807cda02264612fb73d706a726a9eaef498e4c4b4de64e133a42eb85e6825b94fbda86862895229d8e4f466ffdf4f3250825b8cffb82bacd5a7566cdcd944ae55569b4dc758a982e875e2ba2bbde63617e63346737b76c0661c5b017cf3d750a659c625ca0622f774dda44565e43e096d750a807cfd26395c0c4a000e0f20324019a4b2849e771940fa6deb0059da7710a7aafb9e599869672f8fda186f59d9d3770778c312989cb5bd42599639a48ce30ec759c115272f7b18df024f0d00758de8b47a02a022f446e1a410fd82c49d62e79f63a37e2df8080bbd9ef0e67e69a0f5371093afee374754363b724bee4a729dc56b6157979c8f0d068a4b6ccb9fe3625b979ed1505ed21adde08be1fbd8cca10cc9f38ae5f76da3502dcdd3220cf1c0acf2148d32bf55dd28686f6b18ec62cd7c758808b69ce79f9fb032f22e6cc8023c3e680408771635e89c3f7b54db68a804a56d88d2ab2fe717742d533174c529a662560b9c8bb886201b50fd72542a1c396a035313134dcc390489d76be4bff2c4e2ba05ac4ffedeff8eb766e43085a07208eb1a5aaef6d9c4b099b05fa1c36565b35fff18e511bccc414e59a032ea564996dfe3a104bda072bc4b8a24a4c944014e8597b4d2e9bf77a14f707da20d335daa21d17d25c4b4582b3567bf388d01a24d6ea5a7e8473f45e81f5e6f21f8d3219ecf388d598a2c7c15deee314b68184c0edffdb12991d9345abad9391333573d5b1ac588efcb4570e81f0450c3aa4760b4df5f9be2b6f0c18cd599692398099033bf6737bcb61a667b1a2acab712a814ae896bd5a0b759d35ab596954ae3ef0995c580f37da0f084f0dbbc8bfb01548a19c5505cd2503c52fc44dfb856038ec576d6ff5c756ce8573df6689e75c0a1601bd9fd0811dab2b9da9cbcc2ae9ce7f314971298b3af13c0c4a69d883dff4a1fc51abefed4e3590506864b29107bffcd3aed016f780f2cf81c72bb9a5626dfdc361f319b3e4a73226dde0c1f188131ff765fc8a87b230ce3a5d802e1d82f15bfc8a48c5c2c44c8aaf6e06cc1e6645844b2bfe8d8ae850a5f3b467cbfed86b8947bc4d9669ab6f43849979bd34a5ebab83673584da79edfa8f245229f8d84cafae3ad9f19e34e27498cd71b0151298e8db6677a09a5a25d6ff862119ce4b7c1f60bb928dedb2f1130e1fceaa5f2531c823eccec6f89717801d00d710fbcb905d04d1a30ae27e889beae83af9fc0b9c40c2185c9e95e8a8a352bf57ebbfe0c0dad1ddb54f467d644986fa9867e61becf6eed02b4ba79b5742a13e2bc4264d3e46d398eacb9b9d0d1f3e44a68429471048580f3c6f26cb0d07bc4ed91e3466c76ad163f854f59d21e5c82a1531f6e054326daab3af3b164ee622e8d9d9db35aefd58471b94f442e58dc5c450c66c1c50a334b878a790030605d21e578b1ae5a47190d11eb4e9a340b5e0085f54d6259efa5353c9dd7b6cc1f1340032a33c0d485ef8a43b04736931d97168df9b762153729b2e19e381ffae2f67f2a4a8527d4754041b1700119fe65c39b03fa622575126b659ca645c86c2700e35496bfa4593ca5357235844e445fe302e8649eb31654e529f26be8783fec638c4f64a1632dea4d3d076d9b7984c2d0860d7c5113e8eff1c0f64d615c16343dec01a1eed1425f7c4b1a62c9b1520ff035adb5e8593ca64eb09f93f008090d764a84b255ffb66200d3c65dc899de95d682fffaee0fcfa941127c4d14bbe7adaa0fc5634e327d5180b93180a2f8365f14f4573136c6577e88aa28faa58144ad62ddee53add986397816925c849ad5c1731d2474759d6f1a6791a13be1b4151e0abcd43d51b21a8d6870abd74cf52d5ebcd49040bca201480f1578fd56041c85c3bd4520f0e194dbafc1ab6f9aabad42009968d2f2871066cb7e1ec839c13095a8b1add453752edd95acfb929f900d893f04a299fed920215b61243e06917846d1370976fbbe1e7934103bd9ed81d10a51b5eaf09a3481ad521ec33a42b4241c8e692190b96c8ca5d7ecb7d9dded8e060dfa1134d10660df5f24ab2d82905edf3fe2ad19f5260a6efda8e0df198d0382302adda7bf9cddd5eb11438bea55c25ac37be70846e2fe0f4ed859ef1455908791e4d00d78302395142bf372013d5693699cdd357668f1abeaad22c97486c7a0af203daefb96bbbe64bfb44ad88db7479a229fb203655f003cf7f1df078fdabb03cc7128bf1278303dceb16e44cec525325ef1e024333cdcb635ae18c9ead621a758f8e4855b6d0b47e8c94c1b005ad57df47fb45d1c33056099888228c152705918d10c6a069558bf61f4a37a8f9cba745329c121ce8e3f91093300d0dca4c5ef82a62a9f356ec8e12e46e10b933952a05f333247f40ae8475d4d6e1fe561500097ca3e0a0919a287abd57746f5b1ed6ce74abe5727745d032af673ef04b59d9ba1337d3fba9a6c0635a8abc90cbd5503c757aede381c294ae4152f94ebacd38b91e79fdd48d6996afe978b6511535029d5385ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb90340bdf8d39eb9b4af4c72615e8eb90d790962a949e1645a9f97d8b271826e554f7d54fdf4dfdcdbe41044361aeafb01141ead8c586fb9040f140db1799a6c1a7f6fe0165dc3aa8c99ada908dfa96a2d133f9078d95e9057d39af30e7ec12e752799f926b9dbae7e52f94efe79e1cb03c64a1c1646c3e9f0e8a59fb3e5bf065d25136a1d9979a0403249ea82d5cc521dd7d926f94520b83d7f8078c62374ca91484de0d538be745d8debd49b67c2e523c434056eb48bb1f4f9e42015ffba2ff1a94bfad1b435843502beedcf377b4cd07bff8027cceeee3096d1448116048c117557556c6c4f6de615de0d21e8b875e01f4da138a6a3d4b5b137793fda218ec1d8af13b4a7ba0ea0f0393da01a1331d154b20a4d582fd84752e6a5bf78de1d69e5f1cf4c6d38d63fc1344796d1040a8cf7e15079f0400709858dc774a69e4603500c0c5cbcf14df7abca37ed210a32b8afb06620bb52b9476ee5e5ce63bea729dad4ebab5a13aa903cb0ec4df002a3c25d954f8de4fa68f397c3f561746afd62c2f9490374ea209624d1bd7d236d4d168e00603115daa7cc703c72cb221acb3e295c0d506b7ae5dd406c266c5bc3e8aa1512e7dcadbc4b83ba6f1b6016e08d6e58ebe07f18bb267220cedca4c4b9399a3f7194252aec0346788b187bf3e89b4ffac86861b287292fcef15ddaa7f263a9cfc87bd116fe85e957bf7e97dfb6bf96b35d2235bfea9cb3b27ac87ceca0411f8dd38ae4eb83c2df0fa7512344f68eeeae2f6063e72523da90f3057d5bc03d485b8faeda26501bd0fd472133ac1a5b851060383d6eaa53cf4e24ec7a9d28e841de920b163f6f36003111b728aac252987aa2fc8a3c7f1d2da3e389a42261eb4299505349af2829d8b673f6ce61446d29fc6522d3a963a758e1b04883b439fe8d68d393eb6db9d35492df294775482fc456244640d98be547f691a7b62c8d5391d3be3ab7244cc928115abc2d1ec4c1b018339a809c1bd9e459f6cc63cecc6d157baa023a530a680f4b0698c6fa55fa2d63ddb63d4c3de54aedc2f241fea5800b1224d503d2bcb65df2dce5bcf863538f2513c4d1456da0172da544730b5b271e363b8e83da8cbcb80abbc7c343c89b7e5162a87387d7aba9a50f70bf427c897c09aae3807123bc63d7ba6b7666e69f0476aadaf44e2073db1090fe816d49d41a6e47733e044c9d56fe9b448819efe4f1cab822bc7631e594fe248435b32b4116ec763c0fa08c41721cdc832e071c0acf6a7dca9a6a5ded72855bd038defa52f5403ab8e7bb9710b2fcdf24d03c895f902532c8e1f7a604bf704851e564ab7a8e845a0efc041f86eb3cb6a53d5e87b97955f81369f99a4aff0069d1014ee3b48a937ee20fa895c83b0b34faea90ab9b994db23200ee540c2504db3d5f8158ed93ccd9713aa14e2e21a70f71b675a527a0b9c1de8d40e4c6e37486ccd72260aee677626367ddad905735787f8a077d13b9a25e6adcb878f6e0be1c61858c27fff14bcbd93a23a9dbe8fcfbd2f9a51bf29f105c85299e83f08b8391bc95e5ce676ebb1ff5bbea58882429392a521dd038162653bee0be0425ed8222ea21c3912b8c3c3713fdaa1d838bd2fe2c3739f0445ef1d5cec8ef333987d10eb5f4cdbd557431e7c2760d8e6299f3d662e45cd616d8181ec9c75ff938d0514881c83a479809c18716440360cbe253115d61bad96902c1be68890f387f739b6cf9df9c38af9682d4d1ab709715cbca493190fc5ba8e87777ffd2bdf087fd0be6ae44bcfc46cc0baaccf585a63edcb140afa536d81fb7b1126f8c61fe8a6d749fe37cb8147d2919b8529c81667ace2e224d78d91af3819fa90ded56a05f409a1309aa3145f4bc97b51fdfa358cc34586690a8297e67718061ccdca2cc4e04fb4d21a945f18fc32834951a3948336bc2ddae8d0d3da766b52337778aa10f798eff3098343dab4fe25c119f4bf79ed55cf269958ad0cbe60ae31668c4cacdb895d2535f18611f2671cec2c9259a361fd3dc67ab35eb8191fa37bd85dcdb1bb39246d2cdbf67b57dc7e9b731224b7da1ef95239ce87d164fd1d3645943610001dad1258f217e7bce7027ce316f1cbb04452522f01cb9e6a8923d5969b40d5e558422f7da7506cdd611fdaff4643dbd9c4dfe462197762c0a2e068126ac6ba68f5608dce4ced28737d469c44d7753abd8bc37e4e75691e3d9c13aae8c8f8f27d4ae22873c2912825265f36272d04279d7be9ce187d237f11c0856e3b0f4fda4ee93136712ea098a165aceca94d3d5ffc79bbcadc528517d5fa81bbac4fa82cc0060a4aa71055cfddb3b457d4079dbb4fe11cc2db5eae297dc506fd56650ae086feb0ee8207a624047cb12453b6722e6db099621b48abfe036840bff858735a81c826f008a8d8207889bf91dfc8e0f6b33c2982b16bfd940e57192aef1fad232810aa1c0be71e15067d87410527253c238a00faed49f09a87e5d3aa0d99211e6b98db80caf068884a58bb5c208620004d167acebaa957a2af39357a4056a5aa3368598f7d733a8f49c3457d05d5c7c4afa12406299fc290332841f73912937c8fd5c0d7e3955d335ac8629ab4bb3024518f19bd04d18840390668476f9ce7d58a412c9eff1f0a9608c6236983e3ca9432fa7e058762f21e88c1a5fc3a10a7b22c12245dd5be91d423b6af0f3c5f8c0db9bf1e2719e0a559db519b54d64437ec1ace41f3d3ab4b2e6d0c22e283f647ca758c074df2f502c7eba5b2163c984e30ffe87713606fa68e6bb1bab92892c71e458bea4443d046b8288e1058a0ef8686bab89cc31c5fba5df424d0a2b6d739e38712d111cafe540d5b852c476c181f220142ebb48870d45259903e759d4ea2b767399e666a270625f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h83c4f1a7a4cf6a2a540b1fa2cf24380bc3856c91cdd86e92d86b727b7989206500c81108d592bf65c17045033af5e7d4b6930b2e1b460d4ad0d5d4e85f2de1100caa145f0db0732980a494a9905cff49e7ec2dc97ae8d7f5d3d564d04fecf436ccba3a56e0f741973096f2fb302d870e3fcef4082b8574c823bbe7476a6e765f206cefd70c3bbe010a9e57417782f1e6808e98f6e3f6bd533ca96f80483524e146614ff5875a5bb64bd8a8c869ef48d3450795db271969c6a9870c8b599b6f4c193c7ca8ce1644d40a18e090c58722eb81b4e3738a5d50c1d41331545434e0486fa752e13bfd6292209085de413145fa8f0628ec9c0e09fb25e8fc6cedec6b30d6bbf40e6277c23bf4e77b2fb538c458146183f77c11c490050ca35751f66fa316c2ed9814d4e6dc9503705fc76bb0c38d4c8c9b456710eac67215300ccb1f0ae9c6dc08f12bd925f8c40d6ebd766ce35bf69a1f474682fc1dab432e09be337577e34c05abfc71ab238a4dccddb6267bf5cc15c8f2c4a9009f12d6bff9d548b09f01d95a9e0e3a6f4a0936d84a416a778f0c2dff5b53e163ba2397ea05793014d534aface8c083ff45e4cf6ceb37c7c6fb3b406d7a0aed0a4018663e652346aa74a19ad086c5822becd2e8ce1d6f9d20645fd08ad34d680e84b5b2fc370431a72a8142ae5e1850f17bf529f296d3717f9420d0c6d30ecf278e4206156f47e3823f35ae60fc4ca2de7ea3c9abde3a571c7343843724c023b749776230f413f4af2d45bf1a20a63a5825dd177959a82b3add49aa39559c86c933145a28408c9b72b157dd91b322102782894c46ba14b49e92bd3f4bff5758ef38f6c343a887b556173e52f273a6fc1424c4048c806955e1e7955ff128a65e4639f10668de7b46b7f2a1d038f9d3efcfe232c32f90eb0c8b76e02f9fcf95b939977981c7c46c51a44767e175568b39e8f119c016a557e6782b55d2ab49fc30d54cc3a40a16afef8efe83c6a51183972b85f7edd4ec7ca17a8696b01c5f6734876d234f86cf2d5a9e02550a11766b75f8cbd2b377499cabf118bc551947669e7337a6c8a6a14d925de1fea95f9e0bcb84142c07387b7a47cfdc948d7a9327a2dd49a9866ebb741244f5edb0f910e79f2eb6ff7db35275f857631502b505cee78c31b93b6147010999dddb74bc2149bb838f5a296811bebc227dae91c37aa514b6a7ad86aaf2d83258aa4b5948a9d6657bc1fba9bc734ac6dde7c1bb9a3dc05de242e55e15d71fa5fe294ec7e6a590aaf98b5a6fd0cc18a645c762c2951eea993b6ee8515d5fff7f27e6b8429714ede62da955c4c4220f5b6e866e75237dcc516621f4d97cf80c17322d8e7efaa1fd8fc16187bbb7433652075719da53ce0bf8ad6260fcce1025b10c5eba360c00d118e85113167fb245e28339f9e733bf8314b6eeb5d1cb6fbdc82d2aa0fef7115a83826a9a3401fe233fcc4d81cb981c2b42151ca7cb2af339208b479fd0fad376ff1b438e14c27ef2f6ffbea9de65ea725ab388edbd4934faf91a4bb0f2106a34644fa18ba384c5f6300af151df8a4472ebc8fe1d411ad61683755876db0bfab228bdade00f095a23574b25b6e1f7aead91d729f85eac25a0c83226512212dacff3b2efac14761bf493f194e11d7d01fcc50005aeda39bccacd8d30bbb801ce3d50936fbaa2b80588b25ddbba396d36fa06531f0fedffb58d85f18112bc416019c7e337ada418d458f11e4479ebe1653f9966a2e96ae87535188b69d48dbb0332c904de497a9046c81447512d5b47089db5fde41208c41eedc7338a528b7063e7b0faa93b970c1643938af89627ef821dbab9743ee006a49ba6da026ef6862049412437a0a18aaf254499acd28bf18bbbed6877fd54589cde500c0dfbabcb98eb82bf69e8c60a372c7ebaad2a460ce47f57999a9ad351ce920caa85d23d01678d38e3ce68e7eac568dceec048108b23ea3a203511a83a03ff6ddeb00db9bea28e9acb72395cd24a1697306cfee3bafe687cb7a9c250b09d6c81e0e28717099c5dca0100a24b19c5974e4e436f19fce535c9874ee3e5c5fe93da3703e64907b9984f02b0c68fd74754590466785a46bf3c5686c157778f47c383e0c801190098dd6ef099e834e9d66f4bf277c30b353dc713dde1225d26678318b313b7f14be2dfa4bf1d7dd756b7a8196c5d9172536f200024f9b804cefe7e70791077e8e84dad1b0a9dc3f8c9f5ae4151027a872e1212377c4c241823fd987a50b168197e91601a1680b6ab6978e5f9fbe5e07455dad8472e8b18845c88ed997f5dac4684be3a4a8079e97eb97436df908c4dfc2ebfcd046611168d16f253fc5764dbde67885c55f3487ea4c4ed5bff54e952ab7b201a04193bba71dd8e4d0b4d03470830d4285caf5d2fb953e54c0a098a759a4e2c6e276d0c7aded58f0039e01fc051ee2f873387587d27e40d883252ccf4e5a68d9cab199dad7dc416c447c51d95d5d7f224f21eb47211c399f2775786cf353f9281e80b22b2cff68580a4fb0570ba0ff925e7031a6b3f63f1f65a6560f832c3e96bdaf125901b63245b94451f30389f9f217f38e5fbe3e61a5ac0cbd0641dab17abe0812e96c8aaaff257966cca39e2c9d2b64bef7b59987fa2ff151aac8bd27656e582bbbab8b220a53c6fba5fc8bf3b669b94542469a63b9fd8a87979c8ce5798683b17dc191e2f05b2a34b87d507d8721f7cf7aa309d68a839b3674f29b2fc6730f4b6f4ca32d4616b9649450cf1fab26709c6bff1100b779227d1cd475de3249958667b9a3b8380d93f74796642ffcdf40b5761b960cdafe7e08bab92bae3db45d105cd9f06b337de7263a18bf1c1a7989b7c990970390838fbcb8dfe8b77554a04586f5788b554930;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h43c1cad07fd868e2180b39ebf73cf6530cf9ea308afecd02af7c23b7d13fe2a8545ea6effb5b16c3db58dbe2d19935658af440e1caeb87ce2fc027293bbd155184c0912915b2b514030f24d39fb1543762dbc7f156374cd1047488eec3315da2c6a16c7d65e44b58040f10a31cf9b511be272eb7707ca45ebdaf95202c452049e8270a5d781a86dc8b3acc028e34614d16e4dac1d35ee62de6cb8833ebce74dbe7dc7c8c7fb6ca9769f8e30b7b8e99278bc514bef626faf86eb7321b79e6e0a4c9f8e31d39b0546a81b7e22ada400e39bf0b8edd292f3a422ceb27f6050c9d6b9844a67c909733cff00cba636974dfd7e2976b20398b0ce8414957042f7d4ded3a4a558ea9c495f5c0971d7a485efc77fbe3d638fed748c7081f8c06780d093e25940e1b0f855de0497e287b7e9cf42aa3f43fa0bdef52b566283a291b2fc14689b31fed27d5cbd150d0632869b8ded930d32016f047544d83bc54cb039ec4ef30bdcfe9f42b3564f3829c9a39df6015487e6fec0567c18ff9844caa803c38ccd596598d68689c9472c772c122b4fb61d1ef6582b09e2b13a74cb7dfa091b6282fe0ddb6f65566aae2ff55faea62a0a34f97dbbb7e3ecf4dd41d67c02169c8254aab5ff93f87b7ea7758b15f1f0c3598ebcd90911cf58991b21f0ba521c1b08cf5e9120cd002248a5b5954f05d8a00e40e0fb7b6a141f736db0e6c549470c05d1ad39c2d64146abf117b5ac8938db837c2536a3d1eb61e1827542d5aca5a7902599819b53333384b8ea7211c96ca14a767ee789b7044313ad40f04704e65007275d4785fde6a5beb703b09e8261f24aca32ac03cb5fed85a4452b4bffa21f21e464288e699bbbd179c155d66d73e8c61618e6919fa3fe61d1f52a513cf4fee2b7d1399d2aa2b56d1e59bcb58b2d24667f30206a3ebc9e1ebd97d1484e8b03b8863be1ee40fb80641a69fb504358f5f46b6f849d3376982ee664d40cb53b04ff4bd20a827ed4031b9e8e0001fd235b6c97e7fe5d25d7b11edbe8547653ec284363951d6030f3ef50b7f25aecb12c7b59ac5036a95fa07a4ed29bd469b4d075bb46d634e5cbbfe95a2a5bb3149734ab4304f04919cc00ae21f7948c4d170ce0de1d4596fe3fb8c7372b24d1f56e655147cf26ce78766078f85eccbb75a6868ca17003f4667353851c116eb8973486cfd3bf7d4e267b3e08672a20c35fbd69d909637c125e921775122f335edf8cf4beaa7adb0e51c2fb62450dbf8924e7112bdccbd5189eda1e046a12cb9add0f6bb48ff9a99ff84da7b2c88489b0daf61c21c21375b1e31b540df341e212b800ff66ddbe88a5a54713ed53b4a81251138b79bc9ef5641079c7b92209cffff972db4b05806f3c546adb577b919cbb10e5339447026e360e9569df91307ba9e9d7aa6623690a5198c66e3bff3b83fd0730c0982cc8a3c9c644a1885a6cc9fa26296e6fcda0b96366c66ad09e94cc3e6deb0a387b746b623c7b89906f880ed2aa355eeedab868f93e2c4309f498d4d6319ce00ec2b8e4f17c4af8b93248672be621402852af0303c4ae582ea03bad0fc5009799355f8fd9cfacf9e403ad8dec4403cdab572d3c1bb96bfe5de9c01d9a79ea883224e19cd8a0050f77921d257587b5cedf217ebb9c6bbd35f7e40f5425de37f2c6feed7e81292396744155b7b0db9ea7e7847ae6317933646abe1fef6acf31a3b449620bfda6d62966216b66d25a2ae04e6630b481c6f33be04b35950a383949249d74410ffd07df64c8271181d7783c530de58d526b677343892ef71e26fdb73edafafcaa60bdb787e4f95e6ac04d2b7d5fdbaee36fe12937a836e81d0b206d78ed9d390b712a169fea386694ccf8050aa20f0908aecbb07b0135e9fc6ad5d9aa5bf69b6ec7f6768548eb702462253564f7342caebb10e46d1b5fb3ca8c842149bc6a5ba3668a6a35e1094336e4d99daa19e12f3217941aad355a289727c5ae8daf23924ee307e408e2b17849c909c4053018b882cd1daa6be9a2cf9875e11584ca182ab5940ae7f0665da7609d0f0101fb5f5266c66c1212a390ce5e3aadba922128ee626a2a0c22040fabe7fde1640ea69d63d3929bcfd563ba2373791202c0d085a192de8085df0bbe67c8b61479259bb79b128f78005962abb97cd5c5e77c50fe07556c5259d6a67afdc6f8e8889938f996ecf21c680a41020b56d41e3c4b804c62b7758be7d6e53e6ad27d0abc95a04b649f04ab67dcc5dc7c89d278a4e6c1d3c3d8d35964f0886e4839d622ddc31fe2d6defb1847b6f2c53d7f899339c8f969238de95139306e244225365c2ebd377293d441703d5f39fde1a43f548640a0f3bc2788ce06b57db246da631d35cc50b23dd15e75c81e9e7061d181afff306675682019d5f3d8212b01dc354a1f51dda872f143d5b16cabe176658371f8aaa96f84cddf81fccd3e3d596aedf208d558c52752e16aa5bc5d907d1f394e0978e1453d717c6d5efe9cd40dd0f17bd7943e6e9817be92619160a12984a13fb6919002d7006db059d23d1a9d16b806422617c4a62e338cf1450bea6d407c0501fc4061cb2d228a8f29296dc69e83fd7f0967419001bdca06cd130fc61eb7f8b0073d59f467c4177b9571b041bba34493e053fc6a25f7fa08c21af6ed1809296d91c0e523e19ff5fb1e21ddc2c3d2c609e05a063037cc87f5d501062528d23464c30af10a3771a4ceaad8f03bb77a6c592e7fc4f6df0de01e87df952d2d01504450907cbac8faf79450ce10e42f78c61bba17a77b75fe32e0ef10aebb6dc329c6f68c7f34a82e4edf03e80d18ea9ad6d8b339e7f3743086d33699f9c83e8a39bfc4370ec95f5e248606715c8601d05127fd2465d356226213193d52276eb1a95dc2965;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd42215a1e94d3a5d6bd578566a115a502500862c4dbcd6d158f79c25f013b4e205a85d74be7033120b94f94ee6b35ec8873195b3e879e857496a085e02a6fb5cd5f5ca46dc0daedaf088d3eacdeb5fd85f665561eb1922f35d9eff2f9a5e17da8d7c5220aa74a66790ef52a8c28048e2c4e4c6cd0149441a07f1f7d4034da88c79a3dab3abb8092fe518e006a997412a70f95dbc58d2555482c8a3b4d01972286a77f2e6f7660d06e5921c9c9fc94c797852e46dc365f9983095c5e65fb569b5fe32a698a77743c20cd0c760cf889bde509599d241184135c68680440e15210581f369cfffa78a303e99066f970f3cea85d1e39de5581425e0b382340ef2fefa95594aaa0cb7c45f9123851bc219c8ad91eaa0e9e7a4b3972fd9b50270542ea01e30e37b8c1d39fd60ad0ce0136fc7477d2043cd9ab83ecc7d53b3ddb7bf1625a7d690fe6c58029f5f0f50205b23cd989bdf788ca0014f1074745dff29f90d24d9eef64c8444fd3168404efaf235a66269d3b2e0b89902cc94961707e9448deb9d3debeca81904333e61e3727c6d30ae1799732dbf444a8c65e49720ff89377226ec9ba9490aff9385809b60b5553737f3b5476544750552a68fecf197cdf00406569ce7c881595f68130d3f3ac139e3235afe64198011fd959bd9f91705e426a344c700ad90542ce333562e401e8f9fb2e1ef3ae65c9cc686f35549f9f54c879f809a0f81007c0443f619659e4f2892523316e0b9d859125b29f1b7554f80a64205c3984fc5c85bf5ee571e35058ce8ac6547ec5e7f23dcda48926d73168d63fc42b1b67901bae5cac9dab8e6637e3600c6ad757b70ad81cadbefe49e925c96568c21e98165babf99a53eefe8ab7d01aeafa47ceebd789c2e15daf1ba919aa71eefecece8973d40de2cafadda31543c0ec7ada5039944eea1977c525bb91d264995cc709dcfe17d884f66a74254363e4c8f1b6c86e4dc3f17dae6dea80c3621de539acde6c7045d3c65eae6f116934eabd35f490775d108cb881f7f9defea42bef067c7505daf2bee2e5f7b51bc6526b1fd5c5284faad77622a3171f833936aa6ab25f4ac877a9fbab04b22e45aee7a635d1f7c8e665a183d250073c58c425b00a373da6b4e16edb3de72e3a96c09fb2aae0029be8786633869079dbf2155cdc6f28df38fdff476171b507a14054c2a4d51d5f2dd9ffa5af2b8bb817559b69563b8ed1af32932efbd9878fb3b650c558de90f1b96aad67950320f29cc1c5eba0bf092b06db16a992e636b80e966eba2124b9a84e720edb385ae1b9b91db1111e83c23134b569e4735fb8271123ed8c09e7de8ecfc4258f852dad7f211c2334d5910e075d5af7d168cb112df1c3189f7fe3bc4c52f6c1b7d13023bcdf15d83f0907a33058506895bb5b89d2ba8f20516892828cdba0c75988767a8392da6ee76c72d9ec778a3f9d3c23edfb18963cf18410045eb48dded72c2cc2529a701d308c1814013b3893fd6c89266d19bc47dd589eb81acc95a2b90c55e3d0faf196cc0e94b8a7b4ed1dac845063f64ea4a3e6580113b7801e7f10dcb8a6d9abb36ccf4d7adb841b6fb5c0d6c5f2b98c558b2d2b293f9f1705873076510049e3dc91efef83d6a85e09981421797b3f041aa98880bdb30a79ed917789fe72a8e4f314537be918d5d73991f0ed970406621c083d2dae5a0a82e1d620eca33217a686c9f8a67740e76eaf2af9349b46ef5a2ad1d63af9c4075395d019636438ca4a70071348776418fec3d062a7d4206b5a039689704e0015c3925f621d7781e1f788316e774b6b9757af2c66ce76f12b2ac315e562a045a40148e366ce999fb1eb956272053e57e4d0b3cdba51a6add84607a4d5fd1cd9f9fa9bc151802ab740f67d6dec37ee2d309f7cbc48d8aecf7497223fe34f740b2d3339aac30ffcc45339d501579d8027c14d39e965a56036ffbade02113ed3109cff45b559491a3058475d683f9e54358e321c84ca5549a647eff07191606fca86c3ad8a0dfcb63b6f92840b92a0556418e4ff8aaa4b1cfe398f90ce73db871e382c995298bbb1e0abdc9658256973541b6bb9beaa8383641694baee2b1914491f2c08036a50a8fd1a073471e396a0821861f95941bea5ab99d085451fd0bbd4fde5f07159eb851efd9db51e9cad0dc01ea167369c2672ddf5c7deb4ff76b7db90ea2aead76e09e3fa4563d1816b6eddba3a23a2a03d18722d6263a73d0d70f0fdc400360d5758052489a4c02a65adbd9220b65de608edc589a387aa8f5854a472020b00d8d9ed93966f87459d87f53ac7820a8d0901c8436b0846f7e0fa607ed9fc75281b36bc9edc2524a85a18310bd1f0e831c593430c2a6df2736d0343ead183279b4b6e06337b7d4e1924bbd7e3bb3ee67ca600f27c8f2f22eadc86ce7b4daf77754ad512942f71e0e4cd1c66b52c27e2c50e0d96647b56a1f2dd7f404228e9b92e3c5075c9508705fab5dafaf5cab79793995f2ef6bfe72cd51463f3c1c967c31e473e9cb01813d9b207d6c49e9b5ebf3ca9b1ed3634e6166d8aa53c37c95fe863e73829d81cd7b55d25bed875d2facd931f2c83b6a8656e17d65357a6d9453a23e5a176f4272bd2585f41c152b39982b4724f4204b6778b9036a5ee841055c8ce25a540c6613c670cfc3a6b06a15ff1e2201749c8c8b8ec0a21e994e2eb00d7e324270fe49cb71c9f1a2caeb9f576a7164488d431faa1271f120f508fb5d7d5578b9b3d0fe8c685f53d57806f4d300fd11c3cb8da911ea5139cc396c355eeb89351732d8016e57b31b90c51f02c2888bb535c6f22f0220fdea6d2b9b0ac53fb33fed066d53b62925c36d63f2d2875043d4d4af36f612f4f3f1ae0ea95abf8f908ba898293b311853fe81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5d52c31cc94c83a5a09602e67a99fad84f8e2c2bbe63de3956cee4661606f1bcf6d0314bb0305f4c41cc9356dfce7a862a5af896506081bb745a6361d7e3ca917fb9fcb145b32d736210728052e22314130cfe2db43e36213fe785b1015f726b8711ddcb86092459bd43e02d09970b4f4013bb1dd70991d6e8c30729968b34edb82d01795be2708566df8ba9bf4920b00e51716bafe36b3d6b3590338285bfd8afb1ce7da43548b3eaa6f42ab5de996764aaa40acbb1427cc8e7b09fab79732c27e7c1a533ce8a48757fc5dce4e7ba0b769abc194fc7b80f34b2f1ced7a53b5323432cf641677ff1500ddb2442f3bf141a7324e2884534b391b6ee0484db33d3c3d2fb8ba6def1e830796da157098193c8f81e56a4208bc781e4d221b53101869b1f3294e9c22369cba7ee22450a996825712a47f58e2dd702c5d91c7e673168510d97f7c0a98d4d8ccb651caa30eb6767c4c711213e5734b7d5e4926963a25aff3a14272b5e003ef11f69004f7253a9afe5ca8ab53f2bc1237ce231e35eedd1e5d1e062da416822c98f014bd16139a46227e558afae48a05d78e86a47758bda809c001439859861b7aa7abb09a89d8912f98050c058953d90ea04726ff69ef9bd82db32eba5ab26f9a3397745e3e54ae3b54d51ef4f5b5bdbbbf7c2b1a8cf9052f9719efa38eba11e33c72345e6c9e02e018625804fe07a24d4b27965f1984cab23bc4a4d630cccd3a78ea62bfe84a0dcdc3a411d7e60e80550d00bdb8b2628bede36701d76c958a86f57cb506934647000c46cf46e7217053e5c743069949a69374bc7d815c355a9e6f932511de8cb68b8e3ae25005b7f079ff8352dccb9a553c8a3ab9c8c691c51e4f296bac68f0336911b589c5508c88584e5c8bf7629bed8423a635f288c06ff09f7e6823976ba4accac3941e8e0def9fb5930e9e4bdb65719761e99f4855c1a696ab8ef1b4e2eb1a49bb744e4c49df404b9fbad3814e2332ced523ae7d13d1f2f3108736b4044b307f98bc2cc8a0477b3f2df289efd148c42d08ee2823944977d74edcc15b1e6e81eb9ead9751a829e919b7c120e30122c69ea6c6bcb9be8c6a9985bb3d57ce6131caed884983d9e7c84a3a462a392318ce2416df15de63fe7bf7022dc3a677f23d83afe14c82b48317984b036246dfee9ef41181bc602b6b679bc9ce4aa980898a1ed153b7b2e6d6677296c388f02512f37715aa281be67446d3ae5610d0fc0d4fc73489beb22a78afd5f7b849c2717939c93fd3b726e4354756156b3e94e9b8560f2dc19533eaeee9e17a6e6cc346f97573b1d9baf80e76be3a04b8855002c9cebfd492270a811c58bc6fad8214bf907f1bf93dd6ac86cd1f9edffd4eaa4166b2da329670ca1b9b3eef13cefd6749eb71c0460d97f2421c53df488a33f8f77bfbc68c7d6faa24665a0405e84f0531eff831360aec6bd92686ca1b5a8db9fb22d27992e65b230e8d9c8e202a547af2bef3bb15c9ff5aaa1ce008017212a57f26e3dde6185a0e54e83a0b542ba0b3e6130bb62a219e0c3bc91fc659d4fd86e109a698fa9207885bfc5a29de1e5700839546cf6f4697e34b7c1719ce25ada60029281beec24e00c557072847a8df98e5a1990de1af82a4184877df9305b1031668a0d2904177113c6ff46993f5c00411ef159a9dc5527c5c6510910ebfc6bad8e3a0c480fe60e28fc94033db42f55f3ff17c788e8d4327df7dc37bad1ac6935dae5ccde6e29ce0abb2401d8fd2d6253b6063db90b1884d11a10e2c0baba791b2375846214a9356f3a2d1240aef49df65e88b95d7060d1d71b88cf53545e8e0bb6dedaf546469a9820dd814455b690c2e2d6e69aa769992f81de1d265ea226f7a4646b0a3b98e4a3dbf1270df82f00e1a0d9d33319fd936415067fa9b2b400bd801c0338185de59c09910e35cb058715989fb7a61181792bf963cb78bc8098647e0004365d77bd4187580479183c90f18fd4bbaaa0fb1bcbba2c78c1dad26047f1fa1f57cddb9c0eb95aa60188ace8e27531b7652e4aa74e93cb4c03cad9cc51720b935af2d386267c6793bc5e5472715bdad526ac6c5e97e69e29f647be891791cabc05f9dfcca7770c98509788cf34e50403f59fc26fab5cd71edcba54d2cc20090e811899ff9120870744e9986507dfb5a46626e1ac58a908b7ac64a36b3685befd567014143d75c966ddd3a2dca86f80b71a7be96358e1703deb3330ddc91a225c23a304edc34c360d593b35fdf66fc459c4702f77c584828d998ef9d2a580c13a060c59ce7f3c1a9b0ac30beefcb27fcbd9b464ca5b69268b577641f1cdd0ca6e84c21d399b40b67e83c1b1654d605458c1d1a2d77b2550ad01770d1ac302006e52c06bec2556f35d4f93bae09eeb5f6934cf8324cd05d42f6832ddf10dfaadfae06c594fae7ec43f96ac34d26a8e01e88a0c57975170c513604e2179369dc0f37491ce8ee48d7ec233b32413fa84dc3ff991bc4d27c2ac869a7d60c7de1a7c2a257e8b2f44266576efa23b3e60b7c3566e68bd9f2b1cf015584ed878321697f3be31be9231f7d27402cab95aebab575024395adbc8bfd14b892cc204f660081e945deeea744a7f1761e2a12473c7d04d7c22ed73554587711da58206a2519a856298e133c89d66e46a77f6f4e8f30b623c0954d6c8db1c1ff2510015c3f208acd001e7fd1ddc76adb23e9a89debfe99c49e9b54822621d49810760c83a0f14056ae5892dc251aee76d9a753024d05299518fc6bd2287d526b1316103cedae8e60e112c98317aea2a040428e0ee93b9a2bbbab470726ee1ca49376b1510a6d0375bc62120d34d0236dec468aa5592f5a3cc86af87d7898ca205e317c3a51e8dd11a596aa49c52d86640ab29af16bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2440e20aafb8386904843f93ea52d92ce64e40fa21d9ab9642548e68d617f3372682696850244b2a46e181be45e69992c11e40c464b187ec7e0db78e6e65ebb9da55bac69fc76d2fe6b99a162daab055dbb0445396fb77e59348b2e219f4c77a768c12a0f9ef544aca42547adff05e225c5943c3277acf889ed6742880069b6369a20cb90a5f1ee4b35d3f47a64d8190a013684f7c27c67665ad55be2fea57619fdc492097b460bc2b4133412cc451797869f3ebc68cec05aecd234c01f6817a32dd130669b7fb9a875fcdd10bd462921cbd0c3ad781cd6b3aa05a6d37178f0ca35d55470f85cf4a606e4cc445b9a46c0039d3926f91758fd84990c2a63763ed84287d3a141c37d24a65379b03ea5c2fdff45f32d4d757e4427f7de28cf0a64d2df6106abf8409ec466ba023b9550edda1ae3fea518ae5786ed2e872b43bfaa5cfaf0f61af1f602953bd6f8319d343db32110238c3cd4eacc062251485c85cfdad4e02ea6e1af0068d6b5ff53cb2f463f49a5bab7506d57feebfa7dd49e03381ade5e4084eaca9e23bf10e1cb6d48598e44027f16c372e174fb763aa26b43f9253b9a5275617d57db801d1e569ebddf6093e13f4ea609aecb54a4eee50ee20f4ee81e141a72d8d9df1a4fa93bee277fe7b82c044319e64dbebe577649ea5e49c66c8235d693af5bf904f27ebce4f7547aeadacdc0b0f48f39df4fbdbbae1db8ed5569b1a5f6ca5473825b15cff8442bc002959bb2df74b0ee95af863e9118783f99dd3ce9d81dbda0e4219008dc680a6e3c88c67a091435c929d5796c31d54d5f3849c5011f3dfa920613a04558893a816461aeb995043006c28070b42549bb92a2e6ee0f19382420ecf2df88368ad3fefd8a428d45a7b258116cc5bac14566794dfc2594ef135db6a53ab2447131079aba0e85b43038acf538eadcc4648cfd23c721a0701f24263873eb0423674236d54cbf5d6fbbc38738cb89091d2cf13357f2c32e4fc143575cd8d18b703b57ba960e9f35d4950a6f573c9142dadb001fe532940923c556058aa0ae1ab82a9b51d8ab5859bd21bbbe77f784a8ce4c261837bcb9e0b301f6428430f70682726b662b3ed5c4cfd6d89f84d48948f13e18516af80942d170037f1c6703e9e610b623491d3951f964b9363a98fb24855b6d279ea6ec37ce50318ce14796147de541fb5b1366340005a614a46bd382f9f5abefe7c4d2ce9d4e9da1f1608aa5b6b7120998a1af1d3e8b6b576c813e4882db5f1f3e2f6c042a135b2fcc856ec4f05223f3f1775c0910eb153b7a5c153ef83d56a9ab74bade2633484a7ff106932beeee6e5d12bb35df91a8199750443b40dde9a63d7d4c3392491fbf2a6ea01ee7b149e3063840bee9f6fbaeb103380b03198923e6464ece48361edd356217fdddd41253c37450a4c79c625b8eb77c008c05f7b63629c8607c07ac3fc19a2db8c1af35230edee1e019fb929727b7b18755a084fac19aa00533cf35f2914b88823beddc9090607283b75910b1975c54de6bc5d7d18b23bcd71902f4fc36cf35895b60f5826e9dce0710c3700bb185b5a97889d116946804f31ec03c54989eaf1e182ee6a45a9a921af1459416c367b814c445f7c1a4123699e4a594f60f14475e3d8e1c1bc78b35a2fffe72e77928d23fd018be30c41122c13e504ee19a5d1fc9eebc1babe68b0fe313d8fa2958832ae3ff1d31aa52cc82399665cf2e7dbee62ffd4f1e3da39bc5b89196b0544a74d3d385cd444785b63e44e809345e753b24b3f3790ae16f752c21189975aa00f260db2d66973f83908074ddcc4670e95ca0f36c79dd628fe645d62575b050ea6eeb275f18b7fcbf28a11a9f3c8c46b8f7a5c31d9b9d6d6be09a08a9dfab559e6e2249772e030356b867194d071495b448e9282e14bf818666fb2d59206fd768631990c97f871bfec62dad41f5c4288ae6d9d1adb1d3a6849f45b2baac943678931b69e909a72c85731e2a0e4f8e1281c4776686680fd6a6ad59fd8553999a53cce407519c7f340cabca6036e9e7de3a566016ad8b9e4a4bf37594bd338a604032be2ebee0f3c35f1053dacf95326f141fc4391889436c6e144075c8212a4d8d313d1df73bce28b21acd6fd89dd1bcc4d3eeda13061cb020143b4826c8cd4a133bd12a4b095aff0e46134f7e0d69a15bcbd39de1ac016c2091cb491b8a509df73e20ea79e3ebd4d2d1303715f53c3ebb77efd0fb8beb879835b033ba3ce4400fdeeebb682b3eedece74235b7544a781fba662995af66e2187c3b412a1a5a74b974b00d13c0411d1a43733b4be33361949db62206e5b25394708500077fe7c93eaeb468a331921e4aab349875ac094ed818fd8e6267d283caec7b70b41c5075f7f5e4d882269cbc3d8f4eab7578384f38db692e7169d0fd4e7cdcb7cd97dc41f65bab10cc962c1f2d8cd8215a14af28386f6ec9b1205a013a463916ad8e56d0672c06f8ed298bad869825076735c682f4bccae98121736ec84453d5e429cad712ddcf2015f301835880eab8e4cb624718a9fe24825c925159b10040c5b2e3367846dce947766f08ab836c31f7dd96b2c9101f797b1eb11c77f531582b2c912f35f3912839988d59b644a90e1750b4d99d38dce8a00d8a5360814520f3c64890a372c2a80102c962f575fc913e0718dcce5867bdf123047e885e92c5fba3880bad15351ececf7406cfa20568185f6a76a393949345616e0316a8aeaa3a0d4599d625a16228fe3bf2409abbc2fbd6867da34ff3d537bd27d55b361c2269f64555b732166559a2706cd3a4731662329b879425fecf70b2819a1796c94f0cf6224163f2eafc6a835176ffdca53627256ad337a0ef8bce166a4c43579877b77e99383d57417f6e982873b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha2c64242ccbd7f18d019d82d7d53efb7cdd49df248be3891cbea61fca1ba2d39061455117a3bceb95a2a1f628a6f58ec8da92f01115cf6c55063dedfc2f483bed8b08cc478b8455ce6bbe4d49c889546397652cae0813b6497509674e630f398850ff5ce6c87df3c227f0fe4310d0687f12c5835ec8c0c5510d680d662407ae337ca54bfadab7101cddc382698b84eaeecd22347d6980640c5aaa58a5849a880a3a7c83656f9f07aecd40b2fd3fd80002f4160fb881a3f9b9f5d6c0eecb7ec60574f827b6921c6f68f302a9ac8dcd2cb008246f091d5296bcb5e6e050bb6be6431546050ef3a40ee3fc64e28d159a5324e920cdd9e76230c878131adc2f06c2d7cb733c907b0b67ec8b03db4bebea860ad196c0bc6628c2d51c45ab9485bfa24ba29dc5a074ccada231fef034f167866560ed1192c9b0eb4673f59db9930fc983c56eef1482bcb9b6c119b512db25b58fdd92fc2301aa7fbc9a57e17b5238633c2e1d24a2eae8531da48a238ee88a70403554166ebdb6082cca91fbfdb6b39b58859565b08c7e3b2d0880c379e67c88a47fb72a6a63a9b5610423e2d99d44b365f7498307ca2285062de601b06249b62ed71d9aa9694e57431737e0b32789b5fe371c825ea0630dd0946143f0590660f6a19f0f77cca570fe119f70c7273191255df979b9e09f821ed07b70d4d075ec811864a7e6543a10af39432a8b066b79761e94febea8531deb68e4c0773504df4c70a48c31c214c74d3d2e719c3cf2caf3f2957507ddb498f5155ba9ad52251001defeb596571bf522710b234e7868dd0dfda2fd91093534f65b70d1b1c1dbaffd5d270272c7721ae30c10d06544083246c1b55b53c38778729bc0364b878f7f2b809fdfa725deb3aacee20e29bd95fbdc72d8447b3232afbbe9e7f8fd45335027c3f917ddf3f9e43d4a110f4e0c51c21e9f1baa9351e9e35f3e9d9a80ee46577a02e904757756d528297d374c58bbd030a8337f3a05ba35e0516f9ab320f8a7625653bfec40408cbb09975d48d68e7ad5884694844096d6591ea93fe4477ec92d46221c93cf8ca5d91ec86eddbdf275f4fb879497c38428ac772799c750729c7f9942d193f5df82fab1bb172f996fb3c5df471381422dcd19b2303ad8b159c415f65c5bbe46e8f5cbbd7bd317d8492508b5ab13ca80936761f30c315d38fa1ea187f6aebb2fb240beddad87bafe0ff423492c33f905dc9a2b158404885b537f8347788a2acc0aa4686a55be292e4734e63b50bf24d78dffcc5d26aee24a5a7eee1a79ed74f16d2bc4ce169b838746be6a3415f8c9b3b06ce29076618e39d540f1acc01933fe7917fb0662e8241b2ff45ebb30197e4d002631377d5bdd747989d04087d91e6d3c3518c5d6883bfef3e67f53e7b0bdcd6e13d287980123d2c7fb09139437c232d5a8edccd963c94fa31745a93afe9b41cdca3917542bf509a3d65359aa792df278b16e385cb9d8d67d1379202d040336799c7fe7e205909d20ab1901402a9c3781e3cccc6da7800b06bee1a7cbe7f6adfb6e5f8d04a01d86801e3c6e7fb811b3147fc3b3f516af8e64967fbd0859359e7f8c86326beee7ed746954f768282fe909f2fccc2227ffa86af9289c2d60d1c919fb19985b20468befc621d1ddc438b4847f9164144cee791c8b8d1bf00de10e9936013c516893ad0cc30106c223fb1adfcd5ebc5fe9219622b304e264a39f914b8981cffcd191a7c3771eb52e64c9f8200000b7c5a72278b938dd34bea87def6001312d2b642a265b8e5b93f29ebb96fa8dec8d887054e2aeae752855496fae69d131e0f1491f5fb68325e2f6b050f7516efcca91073b68df7376308770774c5a471269cc028a41d83101655330187a7ae464c8615c24484b0211c7467c009202244c1a8a51e168b62ee9aee86c3035727c1c1632fdd6e42e6d274039867507af924d8fd051be723ce1aed67556c1485307137f95b669c3893b15a5da622113d577b256456a079f3418e42f0c737100bc84116e534560dd79282e20aca2ccb10a28bd4ddeaac12dd3956fffeea654f24f5b3309e87629f7c75b7e81e382914ddc358cb772520e2d125b6f457e1d168d3f6e9a85ac5b3d8900c2eefea9ea4bdb3407c0d9f5349896114e3dd768b6d4bfd07a6a86b62173388691ba9fb80037a252f8c6750afcdd5c657ef8a81a95a8a7a837d8bd7a4161e767407d36aaf120cf484c95e4221cc2ea22fc25b91199304cb3c9223e093c699fceb5a4fedae3b87bf9e87d0407f63de69b6f259a30dcae6999eb570b990dbf15933b1b6efceb2cd217d6c743d6a8ee45f1401da537e12d32cbed3c724500416a4921c2c3f5907e1b3a59465fdffec179f9e31bfb49365532399e323198193ceaa8579079bfc6225fc0265882dd9661d4d9d2dc563e04afd9af0d205c649c601249eb1b0c853072e5fcdeac3f7ad250ae3bef6c3cdad591898a1bab27e92fcc4a255964cff8ebe1f72f357e605c6ef894ddc17eeaa42d90c1c028e210959e8f3b3e447313979d98d6f0003493dba73c1233056a8a3dd3712aae6ce0194434c8440fcc622bc88f8e923ea9ec9bd471b87a2e04e28b0a90b750ae268cd61b63ef08788103a07161dff23eff839c05ae1b0ac6c7b8a3c95ff81f72e89db1bc6b1c6bf098e10cab3b1f17572e9b6bd22afb3c620b7ab10a987b7a219f86af5b3217c316028c6257e0c372279c2603f4201786919c4c02cc411b8fa76f29d0f704cddd6afa9e3314579dc5247d09201d14f2702e5ca11c17202f115f362cb4d666c398ef0fb1d12d358517efb80112870a75c4918c3c8516c37cfad4d4bc183420c7c8650320568c8b65182e926673152350f8bc566aa7f5b082cfb7cd90767043f3a351633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb1d3c47fcee9a0ff55fc688ca883d218828cda1be1054304efc9892570930746246b598934a8726b382a10874b6c74eceb2759997d63cb2db42d6c0e20370954deadfb1afe058cc4c836aee8df5ca1db73f9fba6ccff260e7e9002027258b17713a06ddad186f17756e80b571a92b02ca2cec5385f4d84533ac28bbbce16957bb9cf6802cb68e986c9566607c10d8d0ee1270c54f50901277c05edce8566679d8587bb806c097711f65f8211ed4a41ebc1cc40b9697e306bbd8d1ab2a92efac28a6c76b332f73844ea44391d5cab9e0dd693a792e88c91cfad674a78c948514155c759ef4205b235bffdc4019532a0fdb8ea32f4649df7f4003ab219446e79b23683d84b5f6c369d9633560635b8290fd8dcc1f7c16ce9fabeecce25ad0eda89ab627368253392f9955402a9afa246798ef3d6493cf00ce7b8d551aa49edfd996b6ddfa8cd3242f88710ba619af8c3b5cdc76d190529d951565b0445f4c041706b26cc685b13d574de7287325300d928a17e46554051cc9c5b6929de80e8d5393d605a2229a4dbf421a64829f818ebb6d9b34603ae6ed6b4a6d109eef36e506afba09c7fe30f46b9e085428363e574b20dfcacca15bc972f0b2989bc22f9791749618246d2e0c74fc3f230fc2b1eb65c5e4e98854f1ddd694238645e0d96750b9b7062e6c49b7da593559fb97f144e3bfe5de8351e1ac810f127064e8612f40dcf0fbaaa3df4a5205e162ae2a7bb61a4ab03eb033ae87e6a153e357c2ec6e551b207638359bea97c3d16f010ad7590dc596115c79609e5ed62ee944d326762cd6044382ebbd4d4a96b98ea14731b44224b35df895506fa847e394775a7a6506fd4acc2839e2595c59f91146e6fb34717ef75ff27d68e6a42618a43220296f64b020c41d93ad552df6f6d1409a100379c273bbebc6009526d6c642ba754ddd3e6328a05c23273e9587ba76f198349037134e89f867af5173090b3dff75fc11eb16c9395afa9a45540c16b314957019d9a4713ff6e19707d987ebd90bfb1a79cbbbe5df959d6ab563b8958fae1a64e048bd7520a53bbb897c317365f5e2a8d4d2698c6e665a63e09a93a12ccfd62474e19462b14ae50d4d91fcc9202f58328c0d2286398c73abe6a9b893503d1f8887dd5ebe760f339a1fe8ff2c4170f62483aa462c840a569988329338a293be31df1024d3ba1e7c012d28d86ce33583844c0ef64fffece1755b9947dd199463b1418250903e4d4cd879a90d64f978457ac717203b87eb8f13f4c57dfa7dab3a9a74e8941424dfc49c75ef7e890077be4790458aa12cffd0deb78d5b6e6eacc540a27fd2c60971e1e54e16e9dad3304aa904b9bc0cdd78b6b215902c670f8686e74e14a7f7a5595f0699a3ec3415ea37b807523efd09b1c249f48413ec88fa4394f829eafee75c38b1ab4e6875cf52a8f2708e52444b8b57cc764ab5b50b7e4595171dd8d885b2fcaf796714e1ba8f75831b5aa4e198d1f3c28abac5bbbc9b39735a77eea93c5e47d3bde1841f38388f248281d71def6fc721a69e2d08e837575bd18eb25ce24a68b544fd67b71ed6bdf4c85f12afff191630977135d4cc186f63543b457fcf40afb9fd57a6259881e1bfd6951b78ec1d7af1101bc30a7d90756546dd6301bd3308d396be49b3f970adb9484d287ee2660dba892aeb87eb3b09a40af59834511960814620d9ee5cddb6e9fd490e118849a64d7adcbfbf1cb6feac68b09c265a1f9132076b7c5c79bb8e3e452b11ac4b020809c654a9b6add66cf3445b6e3eb38efb1819eac4f1033c974e14d89dfc0153a43340b31232697298f12ce5cb758d6934fd362c11f8c9420d937300edd86b5c386de5fde69bcffc4e2ec8aeae3bb0049ac22126755d4c2a45d0f8b7906431dda0f48d2f23263b543d9792ba59e78771b28e2333e627f3f9c76de0ea5f79be0a250a14b6ee82e85d018bd0a1cd642c2679977a6d67c09defcf9506b9a2afe4b5d77d6b92b65a5f76aeb4f637e6387ad684d11cf5e9a1bd3ee719fb85d64e8ee4c26dbd645cc3c39ddfe916525e4fc6be2dc18fa713f390a02df7ef04688ebc6e8942e56e4c06f1364b053bd6c12f6310da062750c388b925dd0ef728eda99bd0237633d59676d7ebb975b76c022f88f0cea8f9600f87238a142267f599bc46c32c92e8614dccf3b653f5a9f211fef1ef01adeb85c4481cc55155ea57f1786dd7b0aa1db0ae959101fb3391675504a4ab08da3a3a2f324e472f41500236504f45c4ffdd54bb9c177b4752beaa64d849d58422756e476d989afbc7fe78e4519fdad7e97e97e994bccd520bffe87945eeb28fc2b71a5efc15c8cfa2b4178b6d1d4dbfc9eaaef4c814433e64c2336d80d58913faf8d4a44c8119448affb9c3b93a2b993228a1cc4c66f907ee6a870e380a82315a02bd7bf021e60245337e58c29d39ae57d2d7a07e13485fed051faf826a2b0f512400fb0b6dcbd61f867deade9e71ce43ab422f225e127d928e11e0a1c768c51f921a7335c9697c381263a53fe4dc510501849dd2b088d3a1b6b61be5d4f0fb93f337260366deb49bb5878311ba26649d4b65f64c027b52d0820b9d93063c2dc819e6f56c11d52458888bf3796b13edd0e6c3f01deafe08c1d4bf378700a4958c4df9693ff3ab2d2fe0d4809e9a26e2bf69ac22867b73b7e5cab01b3262ddd3a9b0b2ea9210a2b36d6f880a45e79870e6fd92bf8c17aa156b890e807f69e1a2f96a2421b56bbab380175ba88dd48fa142cb451bacf6e3be7af99e0e4bd5545e73c34f408eda649ba8d70740c78809c75eedc97ada2c10b9df79df948ea09e26c5b9177dd211e474b52404dfb5a471a866f6b5144267e531a4bf34454de27aba2fc16c799526697d7c70f63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb8efe56ab25a0dccb924ae086bfc095f47aaca56ef2acbfcfdff2be9a252a1174ba27150b27f2cfcf10b09b990c428c7d384a96353611fbf409802465949041d4b52ae80f909a9f0dc7913e5100d4d63f389067931246900257e437c5d2de40bc4715b4f27c24edb39f979fd0b0158038f342e31bf4790aa57886cd39c1041c85f6583d8d21ac73ac45ab5085881295ef313281ea0161131226554260e407e324a41e5076d8de13a6d643895cea7fc3fbff80bc818cf52f69a9f0dc31e56c951088b79ca21ea0361362ce1043b76ca330c618183ce6516a147bead1a1bd58d37b2251ec820ece2caecc7fec5933af3d4f9fb4bf42fcd4c09b3cb8f3d778192e07eec880def8ac6b8f0c7dd22a4f668821c4dc460f03f6e5288653cbf262fd9f271364dd90c3a8164310cd67ee1b9d292f87a2e10ef5f62303ed0b8d8582a3d0814d260fa47ccc3bbe1c2617691ef92f65eb9d49137eb8a5e9192b0e36a82d5a93a699ab90b3f23b0e197273548534eb27783dd386c9ac42a6a3ba58cb21ee673a2c3caa5d1ecba4f6e18159883212dfc82b56d03c1559692116217137d2f389b64f1984de2e0abb00f394ee8ab2822117a33024d1ed8ceeee1bdb06f6609242b0f69d3dab6c669cdca840e834ce69ed9dbf116179743ca0743a7fe25dc5536c749f17477e0e7cb5c4211e60fbeb8108a389b239f756235816bfa2aa09afd0bb96f33f54c05e4b94b345cbbde92058be5ba26cfd1cca234aadd2c7727637e760218f30d7f629646c0d6efb06fee546736ccecdc8f8630f233c5fdedacf6122e8c9235c3550177f488ece7d02790cd2d56397dade8b39b792b3a93d3957c13cba2e907af93878dc44c8c5fcfb9829a6162a162babd6fda396add2ebcfbfbfcbeae67469be2530ba29eea40b96c0685d9a3dad5703953e9c211b27d16dad1a9f544a84a11fea2a8340a39d62328396ba5419bc5dc7892054fc50e83cd27fb6cda8feb430fe382bfa1f4617176de28715164698a8b1bf0275db57ca8e14fe34c6d8dabcaa987a68959dce3908b75f9d881e0886119eecde4f3da4a27ca2691bd2c08ba2dafdaf0335d83d69eda0cedcdb786ec1e468baa035832c48c4ba67937e8eb776c390c87789c8277512b5602902e8dab226d8b7d249896b4768878f1fde55ccf9b05b24fdb560e951c696897fb1496004780d953cb1336d7939377bf4215df3069fae6323a6c2d5a3b6da6f529a45e126562ac51acd3b4331be66279c944dc057334fcf4dd7661f76dbcbdbe2873ffbf6913580d040f6270519893f9c4b155a2c2e4cd417f64778e8dc75a91dcb5d9935f4fc7d6367d34624068e05b1d0029e46bb11fc67016e4f5698baa6fd8ab9af09983d03fa2e45265a7c2734e8f5e0248a0a9a7f064b424a8af1fec593ea518d02a10be0d1b104d2992e4396d763806744fba6d0328ad9953b239c44c1c6c2928509b00432bc92dd556c8ca42eb1f65827d8e835103e645063f8292d5179d9cfe0ad1edc1f9ba611d1a4abb5d0bf3bc6348335425724de0a87c0b4274812855d03084fee38856b538fde189599176f145121a9a70241360dfaef35c7654b22cbebfe34249cd481708326b3ef7f8d3651a7dc4e045dfb758b21cbbe11feb160b29596d957105919879f1a28f1a50c171072f4dd81cda64cb76e757786fc1a67a75b9c50847f265be9fa6959ba74e606e0549f0743af459ef6658aff34b7f7b1120b0324075da824f3c0c60bdfd93bf0b0fd1b01aa85f07bb9b020890543f0ba081ba01dad7a534d56470b4163400c5a54f8e4f590821a5553a829f6d4aeaa1cc8e8270b3e5d6ff4148d089760423a66991f10c09c0bdf22de43b8e94157e0be65d4abf3bf8fc1c069bd81cb07b02ef06bc8445eda88d5219eb2d587022c4540c886486ab4b4a50dd6cded61bf056eab909059e01aa7f6da575203432480682f3971a249de1bc35b87ed6a1ed157b07488be381d53ecfc7de846523528e3766e52c4e7242d2f73fbcf4f5509bb0a98647fa7533a62323426ecbdce99bbf648f99404cc8ff996ae4cd17bb4a79950606d2f47edccae3ed95e08445031ac07e70b0290623671f5731e0016c0974c8418cbe03e8b9e216e14ee762bd7a62c23dbad10a6bb690750d15b24f327ba7964a599082359b895b69f3fbddf7e59ac10cfdd27ea6451499957dccffc3dcdf20f6ac062469774ad67bf577e6d2881b3fefe13a07b150c1d11f9866dbbb73e9298d46de93cdfa7b29cfcbc1179b3dc0a80e5b73629f281bdf887c58b9e5325ae32318ce8f5b98e00afec9ffcca4ab222a21d3da6480307d7b59c90b060f0c3f37a28764df473d3d659897f3101f4c246a2040caaa3beeb5ffa9e6a7a6a11aad1faa0e6a15f07a04ac598e0c7d9872a141f2e6e389f90d6d984a748e6f9ade3d51fe0a43893b8edca27e595be59ef2b58f77157f62ef08507c9dcd5d7d2d61c8d0574bd3c3389bca969d198b290c6de0188ba2cfcf7e79fd62f0aa1552046e47da84b1c235899c31390ea94115efc8ae936d3f65eb3e4cd829d621480e96424c60116654402a3ffc69fdda4542e0cfa94c3eeb66623428a840189a44489db52207b04cbb363fe8aa54fcd26375dc975f598e9d0bbae4bfb27c9daecdfcbf31b05b1655281eeeb56e919d5737889d93c9e3f86830d2d8955e61c29a92f2063c4f7628e7aa23cd9f6804dd391c3b46da37976da85f5867171c58af1592c27bccc846fe0755d28eb213b9223e55588e615c8950f3b304d44604c3453eec2df0f7363d1b8eb8ff8b61d66f99638a6c2b027813f49a085e256db9b1fd1737fb5be1cefabb74ec3c70ee6d735c63a1f3c72734936a50acf92d64f43f7b47b237ff67553caa811;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h52c2bae48511dfd50eacdf5ac46a63f871028540b8e289ef5a45e2084f338daa5a2e42ceb0678f6535ce8a82b32d4e1af085b1210ea6696ffacd6d3625c3718a9b4ae62ac729ec8f46fe9244e9b0dd29f6306ec897f9d9b76bea226ab40303dbda339ea81eb3ffc146731961cf7d5c9f981b2ba8f5bb6dd836bc249756489fb5dc8eabd3380e5897eff75a8b3443b35d43632790240d5b65a5d59b10cdd0d54b8d36c96b10b5ae22fbe95956479268725c1cd5f326b9d1682438ec96c4e361fd89963ec98ecfeda70863b70f6d8666db88081d9f2be1c49fcf4c8b697f7e34ae238212d0438abec3e7e3bc961ba12b7858101f7ebacc1df215fc41c2a5987838996f5df71deeb548a9b9e556febb48758b9d088a29338813f3b8a039dd6233085470787fdf1d170a9418f257e6ee15e8e7fe2c621fea668ddab91b7478b78503112372826d3f414b0db2cd3b4e16670cb7913d249118703462800cf33b9ef5f068680ea85908bac32d378033b14f95ed5fc9a6d6b6ad004230b9c3eba9ce3b0f146b0ae09c9f1a74e9d8af36949c1c375bd9778337a365462c142f80d56d0397d493b42f55fc98c6a381eb2414ab8b8f8c6cccc8df6adeb476f55dfe17542c0a54d36a46fdfbb43a217b509dc6006d60f702b6164dde3c4eeecbad52e5be89066d3932e1d27d734d5af907b2a414a82f4f60b5d201bce6bbc53353d2e554bc7e4ddbc62d9c1147c4552f9c89523496b780a025cd97281c8d357a9da7b5775d75058d883bc791fc33b52a5774050290f01c3c06d1a6e6f9e4b9964733b00d3dee6e05df887e11484665823f1066dd4fb77fb30dd37a761c7e380879c214841e565061bdd379acb53a0add0bba0530615ab74c19e3aa4e4acf6935b02971a8d3d63972d6552294c52ebb85cf8852219e22cc264901849b35a60aeb9b38e88ea9701a430330e7c0d85720f0624aa81a84e39ce225b5c8ec3c05b4036111b28a7ae08d86d8764dfd544fd75d4aa00abcaae7c3e5117f0a2e0ed9027976ed3b5482981bb5e4d47767c871fb8b3182e93e148f0da72021d868bd2c1dcfd4918935a7fd9216d32c112c16441e1aaae865a84de20b274554d51d59ff3b51d6e950875301dc4faa75bc667b4b49a2976796907c707c697c2b7115ac0a2f3e6ebc93a864381504451cefa3006659226a2a4fbd5ff47a527733bfa451df41233672f6ab0678e525e1edcebbcba87ba3462674f59b57cb6ca18ca782f479431fee72e8fe41eea42d071692f195da1512f9f82360f61afa8d22749a6066fc92c7dcff7bbaa5681040dd377bae42082f3e02d2481195bc7e1f4811b06b2c7ebe898ccd5855f4c325e180b8eb1c6705e5c361e37c5ee759db69a98093bb64c964e46e69a677852c71557b386e886794836d39522b169ad81fc0e861c1782d0088005a70606117cbdd4a352134744b6f6895d5d85e1b05818abfe928ee1c3d1aeccf8b143ef34973e81994dc1e567cba66cb8565f6b89512ea9b92fb76c2b06cda6a4146676df1efb526a567d89e82c5100da18e533d552620dc66986fc063fbae680d93b1041ab933f87a043a7861f001c16ce34bd43171c51f37fdbf6e3bd207d2ea326e74c4d02766ff80aa38b37de73799a5b4f38542b3370c4db9ff97d17c4a08f5f9dbf7c55a00b1f3300b0469291292cffe6f815f2c4db570068c6b4cab63d62057d31dacda1db8aeb05d80387aba794fe349bed519d2c0468ad4384dd7122518689cd537d24efa9ffd17014ceb3b5485e3f4c590589409f9654c20d3fa070d93f4c757540046f2e84dfa0f1e0f0fa55ffa7caf4e48850be94d0049292d7c18268c08b8ffebf5c678ada49f84bed96a91ae58bdd5e0041c20fddfaf500aea20ddc5cbdfa664c46c4613653b8135f3d349a8fc6814f4b9533866fbc739e443c0c0434423b157223c5c81241c73a53ed73fb592c68b31a370b124d7969f9bacf5d07eb677d48e16058b3d5d3c4ce16cf52de010ddf22609ba3727c4f0a87503a451ec5f2d10bfaf020f19e2557b4445d8e05566e114ad4bfcc60340b3bb82b3d909133c0ff4f00fa1f3a7fdca67e4e4a152a102fbf890f9965549f63bb05644b5adf0d7840eb83c1b780dc6d839b8e541b7692e694869d636538b3dcc596d35a25307ce84d09a28522e6affcb75b08b56052ad31cdd3b014d3a829ec0976d18ffb40bb6e8d8e2d3be1ecfc74e0d4006f4e99223ae6b33f4ed8cb9d62173cef842ec34e8f57ec4a4e4c9ae104d76f25bdfe57e036896f77c1d3834506f544ff3e0ab64e1ff946a8f22030d5aa258c9db9848d08440ffde1d79d3b8e077c7c081b318259bebd075931c0faa848d75fba4c5e8b1d39ee4b7683703430759a249faedc107e2f1c1e85192470d602ac34e0d573b672b1f7a769df1c6a361d8ba165e829bea272e00078f76fd195dab6eade433adc523d30f82217758021e2a22b25d4723ae9b6e7f15255ec247261a7f1040f0db62bbbda029852d416d48aba4c6f722415bebeef809c08026d82b848e9aa0a066c8755127e6f9b4af809ead641220ea547866cb026c86f913ea54dc8115c0ab6cabb129c92602563a990a51780a921e156320b370e9833ae56f09189fd1dba444993fa4ab5a222e4245afc4fbee74cb7e70eb924d89d298e3cae859d005ece84705efd8c3b230e910384a699cd526c80647875f5f2ea5e24efc1293044e2b4d8e072bd4edaeb7981eb878c50d162c850a70e25227787ce449b7f355d23c836a603d9079b98d50cf26dff973acf73ae4d7b90953ee1e4dfb619c84be68818584bde470099d9be3988b6bf222fd5994598a4a4c39d17e0445415e9d50f422744f2a68f815519ffde215fbc1f940a70526ae3b4c6c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb531bc4080477060b453d3b9fbafe9012b00aa840f5f4d0651dbea6c1bb19b9bb08e4635f1906f8be59f1d34c79de5ec6b872a743169ad7ba2a332d66ff917341eba0885ef53ce57fe03d2e83e00d10b5b27647a475c98f1c6ce8a01b4c2f01635f4634f2955a77b65dd394674aec78aad4cb63118fa1692712ce8c49c5b63416f91b4d02261220163f7026dbe7cbd0bb0acf9948c49380f0f0bcf4790b2972e80533859147084cc97be604e5c48a1d0936009e0529022df464adfc1395834bcd67aaca9cb1a9b0e79525d54dcfc8b700e0d618230f8621eef538faf137a0b9b4fc73bbcd177e9d0df5cc26c6d91738e4b570dd730338dfe5e886f1389e0e33f06b0564f9c696673e04d3795d7fc1b8c01dfa52076f50a130d5cffc3d0de2a80fe462a46fac64833f259136784322a1c9fdbb4d62762ea0118a800d8d88fc0059c2060e42c426face58de22e1a37f4404da428867ef673e2525a64169f10d6b9722c528d7b3e4149cc02da3c54576bdb319bb12447759b35780fc5d3d5bfcf61f24ad8f6c53aade139de1f44e49c7fa78df627228402678e54947c1f7f5e2b5c8977b4bda3f2de9dbaa3578072f90c4454918044789d88d373f4a8753fc7c7f6f30a65cc49e78b1393c104aeff4ee11a8ff985530e739a433fa7b7373dbf3faa97d4d43ad50d94adff3c5c0a484341b92112f55f122c09e92257efc09097a104ccd8c59be99b54f502e9036f71ef0eccf7e158d5c69f215e96eb543fa3f921fb81dcaa411b937c158b300481062b8dab5f3d74d6828daa6cd5775b9c9a6784f0c4e85f1e9f67095235f59736f5c03bdc13e6d496dc97684fca7dde218bf6e5090fa4dc3e6a09da2b8028c5ddead1f5b1deb22abd23ddd4aea5821b9ea28d96bdc6df7e09eabada48c923e52858571358149bb0582dff7933a55b0e13ec51f3ff84f635e1e1ec61bc7314f29d66dcdc5d137187b1ca95c487bf998a0a5f8ddfaccd11d1ba93979a3bb3b1bc1a5679775f52a3b3023b6a060892929c1f62d30fd5d78018262e26ede7b9b8bde128f9d30fcf9c7c8ac84ce3a2b0f0083607018f9295b31a7d4fe9f2c346df4ea30e574b2a2740356f9874e3a4b42f6a30e327f210554f038250244d547cfb03ec314bce34823889661c2d873c506e2fccc03696d4f7186e90fa34eb367313f344ba11d94057497ff577ad93bc59db119c28f636095cf3c0d76ec3509bee86bfe93cea76a183be417f601eda050be9d92a4d8d49b41e790b537a9d7e5802d2c68e6f88fca529c2e20fce9a1f3003dd2a4749981de4821607335a4cf1977d8163ae450eb72bb6db1b136ebf0b78693cce736cf4bd20588ac6c377cfd1f45cc214c56e9e64918dbab70df55867d4757e869b999ed0d312071376ca9347f070e6ffd595333170382c56241ce644021728870c9b27a6bafe1b822e32683d5bc570f580806031263509d99daa00c779b416ad662e442f945ed86b5233b3eb712a2dd357e92bf5f0b3a3c423491fa6e14110c89cc938c73ea1bc7c1d09051c3a782970a21d4dd1fe68ce2e0f0db66fe43bc62ad2e7846d6baa9b70537c0721e350e144903d93c6aca51cfd109fc2dee67fe1749f5a24585184b58d611bed605ee87789eb51a796e3f1dc74ac5f1763db11ea25b9cf323ea03523dea4984a2cc3dd8b83be69337aa1553fecafa946927104576828facd1f21f6a01207a752053c781577f39fb14b1f78cde0620dd4fc4c820ee2de529c12ea74eca689148d77dfde7fe00eb696b3a26dee704448302512de3500a1675ab2bcd9e6751fac18970f742e1d87524bf754d2810600717f1e2ee05d134b48cc780f87e5895791ad27d51f514e6eb8a4873818c8e0cdf9f7cc5941897011986a0df5787ce4114095763e70dd8e9c6fdf22858ba0d455f17a7130ae14314788a682e87cdbe81fb6ff6d8e9ea51cefd5698257e1dbeb0d01c811fe93557a1bcc68ff40f1af50bd2c83728992f5fa1f5dde6808185af4d35d7b3bc56f255bd98c70c3fca474a9269420827eeb84e9652d76cd91895ae70279ef968d9d887d2b6735ab51d54aba1412a761546be12f3bf0c9101546c92a07c7f3112d77aa82b52fdf762750d81e850aa63e4b4bae1d6b47253256a5e8b7ac466126793d47070d1b12d73a88a231f4eed7d1498b815f99b4268100f2ce6a9d6262c53917eaaa901cb214373f065b4bdb1fc677801f9b2c4f2f4827462f163b24ed9a5da64dcfcb8f57bb9cbd42a72734d96a2f67513e72d3126864bd414e742a9601e81f7831597c491e3b582e885a670ec935aad2be989698d2166239fb2498378779aa228c7af2ee9512893ee9083ad320cd1274c0183394b09a3ae9a3c8234d9b36040a5d152f78e9dea44ea69adabbd564ce95c92208e6ff2eaee14d94bdfea694cb1efa18016f86889ddd7f2bb997e80cf1108d5193ce247d016614786e5aa241d3af724c2c193855ca4cf643c3b066c88ce7665e7c7d57af07799aa34de6839c9b5c3b6b01bb621ed74768613ab1eedde611df5253c740afddb80ba765245051c93b78fa06872def9a2df28c526730501baa6ad5a81b453ea90ba15dc2038e0bc7f7feb4e7b472325666a19176854072ae2b9aa3662c087ad45c9edac23d4703a3c5115650f13ebdde0fc5eed7328b55290a4535f089625d5a561438a2de87b4f3e5bd1444e4a1d0bed60a2cf9eb43090c78c776ef6dbe77762dd2d37a302e36ddf3e31e3bcf916f6cc35ddd20edc9023031630ea2bf84c380d0f5e1ee036a3721f55954445f29e9f7776daa37a9919a1cf9037a536bbb202ad8a72d511069c95eaf66880785d9c585a186d2a1d4e4c09f6765db8a8280b2e93f6675222a19de729aa741efd0064d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h36975894161b86e251cd7ee64bbddb62c794a68b9d3902f10966853b13d31ca2090a416e97c29eedd06607940ee28b96f55de51ae4aa9c9f03b0c3e62b3402cf5eb7e2ebca6fa66e24aaded72d629a64ed7bd43f6a19980602fa41141e39dec7dd31448f50568cc028fbe85553680cd9ddca0809ca8095d2584e3b333ca89e4534caa6d9468aba2c3852286448c33be2112d69f6a5fa5c5cd87026f9fb31d122138940de87bf9e67681b4b4d1bbe94aa63a64057e9392d0387a9f51db82cf85ebc99bdc4c712571efce83aac4db2bcb78bb133a3578c687327bfd6e03491fa0e3a31580e6d7383343e9b95865388c25c07e4a29712f8d2036ba05cd9aafbd5d9ac75ccbffca7ee87aac8a823a2bc848db4522aaf9f46b821a4b77beee3fa96a39ca4836ed50d4a926c95b21d399b27e62b787ae00e9401ecb030b0e58afeb5be0f9b3339520b1f9b0930475d933e5c18ac95297a22cb8ad78a724febda5057a77eb441396230e1ac15ccc547987abf9b5a404f9cdbfba572b89692a542a144ab3a6d539053be77c55e75f9738a363e8d50910b1ffa0e8e1a0affc5c758eb9f81a644c68d250c0f7946e1103fb852ca88a51456d2cfdfbe6dd851a6e28e603789077e3a6ff2a7f69249c4e0f4309d52b8146ed787c3549a1e3f17a977130d36805678af10de2433a6df8573614e4203f7e196fc27b6a42bb69e9debe9e6618e29bbfd712fe721d68fbc391531b0f02fc77135ecb33ad7530517d23c5c4dbb4df9c251b4a3c837ed978e62917a98e1532133b282aec1f520d14d877106e84bcf653200d245dd39c1038928ce35cd18864c1a78efe2197e58cdc169cebca955079d1a4bad1ea9e1e0a2790c2c0942eca8b22ed7ebef5f774d679a47254b3c49b82c00e119ab6ede125e87205dce7b8929f2afe8e800f68376cf89eac08ce0742424be5be8a9083d1dc3520fec7e462d98a08b2f665f519371a415fc03889bba132180757983939950e0d0ff2bb2584c8790325d69ca3ff870c9999ed1cec7595378575b6f37cb0b86fa0b4654f90861a3cbc16bbdcf2415bbb083855b73e1a55f53f9989486b455873366875c253e0539f98e5d98ce21ba2a787ab6466055e5a4c3530661a1972e972f089d0a90e5ead2135fc5b1569e18794bf591961ea559c5e7013ba29526d8e4c93f6420d52109db237fae75f7040a92ec28434f1f1d32cd9d6c7d8e39e6417569341d1d735ef9ba9abe6a19bf07eb4f9490f1aca216e2c21bda5312449be939b8bc5c29da017d2f2a378c9e0d6204ca5a96a4781163aedf637f04455a7d04977cf825bf70c7069b029cbc1510134acb312eaaffbaadf29393cfa4a2812bd7d3b2f0f7bf47683969a21b03edaca3485870eec6cc4d3abde02ded94e837920bbefe65da5403d06a6b12cc2e9b55be72856ce7885590a7dce1a3482f5b29754330f5dc32a78d4ac31e7b590954b8573d0dadce9a8df1aa3a6f9fdc23687c596a57481237c91f576f5f71ffc19e827909a06befa241b943ef6f6ec3e5743f0966bc66587bcf6e433a739aa7a440f516f71f3d42b123cd9390861bc336bebb881f7a379868ac5fda0582e14101749df455985bdf059c5cd3c721fa1dd6cbbd5921e88fd6c13946fc3fa612c8023649b392b7c3faa878670d48245bdcdddcae88a11ef7092e49b631bc2dfc58f49a1cb62ee3d03c794c29c2ed48828551768c6ef5d9a2255b6f86303cfb1ca47a24e76e7fa5465be6f2f2a965c28cf41f16fd53b56a0598e1bcdea8f86ebee2aae5efce50b9c10d67c332955413f93138b23809989212315d60c670b5090d65213d4e1ba4942c95701f418092a8dffb98d1d49287aa43ab4a5182e7592dbfebf02fdcabdf4d0c136ef85b5eff3a0c2b54ff420abd13d869976ff5031377d5e0819ff98cdb46954baee1cb2a6c62d3f86e43fa918e1e676dbf1ae76337ce52499a71081de4e8eb72c2eb1cdd3d7cead08b790975ce96660ed329ae9b561e1b8f6ebad21ae44cb6736b0dabcd664a548fd0d916a168b64a9ceaa1256ae27724b3ea7073f8845af8893db8fc7d4899e64ce98488c2da570606f4b997d95a4d3927c1d60d4cb74986ce9b1b4527cdb7e11494cbe1d0b8356762d4ca88352f0b7f67dae06e7fdcff8634a003af14ce7c87092cd3ac3ddb3d407d808ec42c674ae6fe7e10ce4ea25917b455a9f85fd64b5b50a36818df9717441182fb143c60f2f68300e080346290966cd435efb67fe95fe7d8c8d2e688b5f73da403ad62515830f5ad5a01691117a6321cf25f65b3d84a396c45e0b806e905b00ff12203d1ef7d788e20e4c2c12327cde28383c6ac8619133d1f4c0f90fc8629ac39416ca3bd5f2447577e5d2bd9905189d927123076ae918379867a69587602b677823433f94b8eee7670a022c4afd11e8e197df9c31887a011e6123e22e3a80c98bd862051c5619ff82d82d1a2c2bb3783e8a99fb4749bee357627a428fffa19492fad5c7edf4d3867a9c22b08605ac58283ff3b14ff358f73c5755f2e3f9937c4b5524c69f3b3377fb80919780c05ec6c8af33dbbfd252d1ba91c692cbcf7c0854ff27c5be5acd7e328e9e028d59ff501664b3a399b00c77514f7ab5c87482fc322a3faf238c5959a8f0cc703a0285d5866bca4d6dd92f7c3294ce559ae58e66a364d1a641cc23be2822394294dfa1f6fb4247a7ccb3048f484b507a3d06f63ff3e5ae142fea45b2db40d7485ff2325ebbcb40e70918c9551dd84d94ffb35f8190e8909475902bc5e1c7d3ddb4486c64dea6cacdd9920f6621b0896d7d6fa6057f4c2c9e55a51b56a64df0047171f4979b1d0629ff8055e6d93c798f559573391a378219f4bd905d675fb9c6b2e4491a455eafceb37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h998f2b1229fe53744e2a59039445a6c8581f7f9290173e594afbf8c1e7b0ffcb7614d78625977b02f6a8ddebaa8d88a5122166266454e8449fa253e21c8fb47c16fd9f9e8df05004a9d5065d2c23c30886696c5d2331115c7b893164141acf6393641ad1a2f812fc3adc2ee34e98514fd0db84497a3acce20b7fe33fbc62082640d366d53b490176e898e1fedee4653fa882ff13f286f2cb745d5ce8ef189a337864863c25dee5b167bb8fefb45bc82aff1df0bbdc5d3caf786d8fab160e6343d3e015d21c8b70130721b28e272d663167613a295932ae4f03b6080cf2d0ee508dabd6ba77b867aa81cc5690de8ee12dc6c4218d6f79e982eca2f793005d08235f02d66e8cee05dea742af7d8efed16d4c07c9f5d354b555c743c8729c15e7556279f82227fd9e78e86413b42b65c44ee4b4c0e4e3fe6c7ce4b13760f4c40c6341a438b7743fc09a88090e0d903c37710573f0584c733c86f00cde36eab8d1b9cbc9d519d1d7e68be6dfaac617fe22cee89c96e4e6051636858fd6cf908bad787e0053425dc5ef67d84d4fadd557f69c87cad76fb2dff747fb39e462a838694973cd17e90b62c4ef927ff8f356fbd9d48148dae80e6c52ef8b32147d7fa0b527fc1c190b5fd1c68ad40b4d9e78e693b3e991d2d16fba7ee862d486c28e99bef23d9515d7cbb7ede6b0a7b4fd5e5191a1a74a98e4b400e12e3cd39261769ce0caed52872624480cc17ab8140719232f8fe73036abf5f14882bcfb5e08f56a462e17a2fa4e49cc3edb78102e023b17b7ba0a73dc2bf0140343b6bee3e67a0e54fada32523b318a960a986764f2127fa710435afc105f81f430bc72b1aa7cef12ebd947a1a5b1dd25eb2822c5a1f610e629b6e1002bed1183f773c304b91060722060e5959b45abb79d1929ea29bf3abd0fa0365f56ea46f17a0b0ea26a9891f88aaf3df10b37c2e2caaeba287acf9d778ab2a152227dafe0911c35fd6d3d3a997316adfa90da3f7691be1492e5b8b362676b29680d8d1baeed353481ce3925266d01f7481a20e2b357204f4ab4290ec74d1fd5c19b4a1bc14d7a7a7da7623544ab57c6b95b6ef3c351bb913872f6016cb4a53834cce4371934d0577138db70efb29395d33f006533349572a4c1f24fde8626391c10cd4e00205a8cbb7b3f11a7a9be5ffb4a928b8b7ee745132a9e0dcfdbb447d92bb27481bbe5131694aea29a901a039e44fa9f993ed049cb87e457c630893bed2d080895a28ecb3dff129e8becc61d0e42f9d19ce59832db18bc167155ab758783550dfcb68094b2847ce4c49c05218e554dcab2385f778be6d5a7a5664f1755166eeb0ccf968a0ff571d0f7f15848e3b7b0113fac5435034ca1bc24281aa9d47ea41bdf04cb4d43e751fa6791f2f8c1a2268eac5731ecda783f770d1ee178504ea35502d61fd339071665e36dbcf8fa0572e144836e28e03653107dccc6d89e64670257bb5348c403217cc66cafdc25b64062a0df0ce56ddd3fbc8676059dd981e8b2f3cd391201407dc35576ae32fcf02eb9f8a91dba718c44b627f710da71300dcb52991f7e51076d7855f999d404118a26daf5b835a263126395b9a75a2141141a60f2714e2e66c82c4d923d4dad7babfb039f3ac6e607d588f13688e82548d7d1209c877bebc261a4e868b83a98222f39ff3a104b27b85531625361a07eda514cdc8a4ca5226992c722f69629879d2118d01edb11002c0f1bc5db4493f467f2d2c264b9673cd44c313ecbc51e3b8efed986bf66be41491570ca2dc20dbb4a70cf1af37941a3cc464f2cb04ad231f7bee649760afd94116766112557ceed3fae7f0eb2729149fac6d308f4161dff400f3fa7c50b71873c322e8e781c93b8a690932648c386c521db2ffd473e3b8db2fb38805176dc189b4d4ecb620c16cf2b612bb2a5d8954023f9bb0e4bcf66b0ce37f07fe0265f2b7584e6867fd016b6fd4e6cf1f9f5895df42097c9c62f9b1491358df7f37a8323542538f747ee453f948b9613247685cbec1e2fce1df9df52a9c966e2c974068114cae91372eadb4c17a15a02ce124c7c8257eb0c994586a9bafa88e5babbc904f8e5c195a1d0236013986711471a87b4c3cc79bb9a2c662c066ba40b51d89c20e965faeb819c849cdbc49d4c78f60b803e676c9e4a396c2c84d4eb315e82a52f8dc86568741ba19a03911002c8ff97814c2e1b7fc07c7648c82482fa467c875749518054c59bc1b35c8bb800cadd1376d8e02b6fd734a4db8da5981b0f1380993d503dc8b535d6295eb91224359f06ea75bc64fc0d3e94696d7d574bd6cd7ec7b0ed03036b17e3c52111c262e7b3f69c2d97bf6f2992790c473c0b6f1fbb1299e808b790d1164656676982dafb60f46cd61783deffcd92c268b09fb9dc93a5903abf23fd6c74ea12c2e0c4c3284c2d815710776587ec98029ea9c65f3614f93bf1dcc83525e07a97210dc091c096164fe446c1d317ec5decbbadaaf58a31d974ee3e5cc15f0ee5639dcbddeb27893f00acb8a07fb31d06a042fbc61e8432de1cbddf1324e941c67a3762d8aa48ba112e5c8a3dfc56f29c98a4fefb020229f9a8dffae223347c453a5043d65082c2e1c5a4a4872cd01ebff38031ef11321b047e44b04ee9245b524e0dd4f4f61659654c7a37c25819673f8ae301cfa768412d78d648bb7262e709fa37d52eb8218e5629ebd0adc708b4de339c6e0662c81c96c18e1462fd4658cf3c4a3492fcd8c3b5b5ffc66b4c66859c794786cb56688b2dbf54fbc5fbd2c7940153695479b29cebe30c53d724cf49877c9cc858deaadcfd377a2c11dd55d3bb543a985b9cd1ee643f42166d5c0049887d906c50fc62e3e08a38870a2f8a007829eaefa326903ad86d8cdb0e858a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h53955495daf8ad0d5dc4de97b45e8b1f07a315bbb20b4928d0ddebab0a09949bc2d811d5e3d3cc93f5d25b835fadb61e7c286e4e80b163c61fd466068c4b09d0614ee03ae7eb5716aa77eeedd1be57fd2516878fc91db646938c37634bd26a2c974f94f073af7da2c711a4513872738fb547fd6bb974b972f97b116a4e42ef13eb658d676c5b7af43db545e60edda0463b16a2f03913df470139cdb4fd4e736f8d1f577c46aeb59a1f5ac4662b6dbb97e05f5ab9fa48530b5273853c6643573f093e07e02031164f22242a97394901b51dff6b7ad14534b1cdecaf5824356e199b5e2a2dcfca8e147131f0250366e60b5de02d69cd9fec5772127d716de6527c8c492c1fb185f6e1b30fdebefc338ebadcdd2dac7495e5bfec9a232a030c8d2aa55f87b5d9d3ffd8a6bb4c0d769620148d1c8c069b10b7cdeade64fc00d2a9dfc11f475c95034db616d8405ba1aebfaf9c7303c66eb77f821ecbbd0adaf11057439d4e598dfafe4cf2990b28e01c14400ae693c33756df8762476290f45e3b8d865bd4188e84c9070229ec72f94cc40e160d4858c649bb6d7caba1afcaebee0cb97ce68f10fdb0c8a970a74da16a03536318e865827190ef0fb0070b6d095509f089811f72415d5dd2b459a3a7432a33069011870e6537e08690444af2fb6445c0d0ada78e60ed2d5266b62ebd4f4f4635ccab46cee00ce7332ee3e18e65bfce2d4cc1d54a10c9a73ab3f233545e7ac174ee7e3d8917a98f3ac6ed35300f7f56710564540e1797b719d2dd07fcbb6451b5676d2ba15c139f24f346c5cd38a6336c25e7cae656e0b8746f516667383052cc4326d7ae3424be359ff2b23630a0f37547be73d5486244ca7a57d16a7518b8a3b2ff503b221eda4cd9d0424b2808491f331249ffeb6d6f8dd738685ed5205833a2e07669095c3fcba9e63fa3babb7330e83be6692822aa7d0555a5fc473c489313112daf1898ed50f7bba6fb26374b5edf3ec32c47c5cdd83b19f128931dd6a526a7d4395d4ca844b56efa919e95d0f50bcaf503a8188806766da7c2ff3b81fc6f6678626f509485022703a59635cb00f8fed3d68cf42392e853c7291c656b1053662c6fb2d6032e66ffaad469f5ef5714f8f4df27dbc85c6e0423452d19d525db40bb05837fd4c24108839572e6e7e7d1bbf990032efe2ee4548e3499f49908e1e80d6c7cfe2696d1be142d34f535c0df4dae8d580cfd8a99fc221fc9befce5ccc36b9e9f5a5676ea6189c00202436890e9ed704e6ce93df1d87f655140ad01e02d142b6077fcf58c0866c23a5546e48279233dd4a0be21a86e4e91fd985262996d06e49f015830847ec217b6655fe634d385b261467bc5a97b93469287924887405354fc5fbfcca5ce8cc9d2d712c6605ee801216573cd0c886add570b8aff289e106ba4d03f9996494a36e388a853a9bce46cfc158299a563fb5156b356a2aeffb73730d14db496de0b5f198739cf632e2996784198e821e4768301bf0fd64998eeec211e6b762c988e35078cf6935f87e6ce627193725aa5d89eafe9d5cc280b6d10298d155417b7b8e1c059d24b0a02f32666339e515fa7977632218eca9955aaf9c8040d4424ef3e47220f689c00bddb0c7ebf99e452f5bade45d0b1e659aaff417f5bc8cfccc240753109362f902ed70369fed0c20535cb1ecd235b01ed911fd72ece481539824a58ff34193198a10bc223691f94920b17a90db7dce11169ff0d42b70149ee86976a6cb30b0d5479a0a0d87002e0658b9b736976cca95b6eb3dc4e73143c4fd9be42082e098b074cf63e30ff69343702d98cda20966a8f3884c7a2122be95205bce59f4d20f6df7ea7b9f346d8e275b472f3849b38f586f411bdb9957aa880b104fd649f8ca0b9fc18d3c71c32640ccc58f7ef3a9d418c87320e2ab0d75cb4fe057a231e7d04bf06be7717cf285e65f062f58f86a89ac8986b19cc9634700082c364b19ad01646d2c6755228f113090629ac9c86f26b9141c020aea4bc26c90c336f321c68689bef67fa1f485d3fedb453794994df64c7305a3c087b624a12aabde74f1f167cbe2ea8b0339873cd85d841e2d5a8e5c2e6a266979f60bb012f52be683420534e2fa9c1d1a7eba1d2a46a81d7640d260e734d7ef4a63266bdd7d6cc0bc0b8096f0eda0d472f86ab00fe2f1659f052ae8bd03133bc8dbe9692b43d38f1973040d1cbc5b848b608fd4d05c927e027e70f8b878ac215eacbe56c7d1628309cae9b5d7eb4282fdad777339bbada25a63339877862cf8894bca7c35ab50a3a25d11d7889c625c14a95b8ad96322e30d3dca8baf9e2fa2ef56a26a205b4826bca9cb82d4d11725920b5351a014d5f9585f06d68912ab099e3841ca6ecddad63159df806a8ca9ceb73fe52ddb7cb948095b1a3a377c40ac9d2aa86a2e4cd5a4e859625da4df00a94e6a5eb89d974c501437fd51cba551097a975597e6bf89a2e9c841828787448c54fb20476cbd831d8ff618599fe04ffb81527641668a23b491390ebf0db6b18b6c75594f9460209350aaed4c385627f68c389b4caa288d8fe5287c0aa3a86b8d5f5db4f0e82453657cf6afe648e7c061aa7e2a667155f5ec98081676f6b733754f267ff3baf94300611070fcfe2ec8edee69f2a2ff064d6b4c2a5f22cd78aad9d26e421ee2476f5c66ee4ca14473ded4f976ddd52d9ebe4f96098d9998713d43a1e3eb32672746f2d059e92dc5d967b37dca5e42687c4f3e32e202023b1b5ca6356588ae001f3d2660b62d935dbceffecb612562ef20149a29c27db1ac6239018a0be68e8257ccb1d88ecf20296296089fb33d2be78200edb2429acdd667e6d5459e819ce2f7bf5e7c01d9a5027db0e59ddf1b62431c5371907fe02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he9bee3438ae1c9f7902c4b8c82be0c0d364807e94095122d747aa9fa7d798c89d5ecb268b2bbbf0924dc43161fd2de57140e5c89a3ce0f1b428915bb452cd4a14da2271408147e0a27f457b8f73fdb95fd962c140260b91a4f674482aee7594957d8d03268059f8176ae881374b110735227163602611b34c2a470fdc395f936f1d458c1c3eae42f39f6d8b38394313d0734fe72be2e063e9b9ad57c2b4d70ca4dab85b2952bd256cd6dd18819fd5a20219c9bcd164597d5ca6cc5caa55b68c32ec83a5ab0bce6b5d70558e0fd6d45af6a0049bbf503a6918b6e885a2d951a544bad0a93c17ec42e7d2f183f0a9713b07b4950278d0bfb74b3d0871882da1473c9845589dc4fb4fb2bbd081253671811ae80bb6dc8685bdd3b8b36ad43fe217d7649a0d7cf3d7e17f7546ac700ff733e977a902bb7e843af4ecf95d35e9a8a0ae199a6895c3366614ead3bb37c20763b19340a728788296c70744d9c66e00f01db02476017283710629e491f38859b59df42f016e911864e47334d75dd115dbe5de7fd6ecc5ccd648d4bdb8669c9c186acb6117cc4de1e463372852b265c10b5ff84145e6a470725097a3c20b763d7966609688c0052c073d9a28a6dba77c4b41eaa6cf8875486eba2955aecad6aaa25a2970da1c7a0d5db1bd688412ed31a8653abb6b503089a8903b54242b0961f526df2872ba37d0729e6515c0c4b15402bb12f2facbcf65705d3af55631329ac2a13ffd4fab56280a02501a9ff28e44e9be5ec9fe2cb3674ca67ee22315f046fda7d0de8f38e59889fd6c75c1480a68b0d352c2fed4eb013e81f820b525c1cc8a5d442c7b4e84e951714c6f0aad742dcae82dc0a0fc03d27798a032dee435c1989f187519da398c42091f630ca293ab91114e15850086134db32466a90fa7dc0ba77769bc3d2249281a45861815f18214827346a076f319b2cb86b881f06d5359e1fb9431e866bbaa3771559d89e3ab6c2e5f95b576d3d58b4e63e7ddd37d26d1ec4ad5ac5d2af382bedc28a3f2a255e3e3ad5347fb8f17a9818c6062b6b1651dde2d3f6bef415bb3a32b6cda8eaebe3d5d6ca832965fec4fa2ba41733834e1234b86c8d9bbe013aa6ac9e8555cde0adb14d9ef5f50556c9d7454bdebe097a9f3c4051b67744f11ce4e6b3fcdc3f7936fa8764f63eb12b17437a5dec58642b73996d0e72e0ea8d173c0599fc6076600180853cede824e847e6f4d6d128c8db9e61aa1f163fa83e7c69fed77b68aced6fb599c63c4d17caa1eaaeb2eddd58923cef4c5d1da7e38b893204b54227a8e0ee6e9eb89d10f38050af5bcab9976b75234d390260c80ae601c4388c4d4d7d81149e895e8f5e99e63992fd999cbbb74ec575da22a830556b41689d0e907eec822e3055fe8eb576e9c03ff77d6ae9b5e02ae37d287965f30ee3979356b06ecae4407090a0c0593ad6fe72c00e94183e245774fd251c65e6df879b9c4ea932287902791d5d200ccc982a0b6f3bf88c8ac5d709fa2e766d112f7e3a776a8366d5ce41ef3de54f19098c6293f841b6f1e8ad7810d176b6c8efd194f32a10f362890eb6ce21092c869d3882cf3bfb68ff8278d235915bde513c5e2618acba8a40dae90ae33acf3acc9a3c391ee13f90707c17b5c4bd38ad26c343c865687df175cb86d4b9e27f61a6b00293d50789c6c5cc58ece2cd252585a7c6e5f701328bf07273b4bd0f05f2c12cd535db35c81efe27423f0e64357f3321df9685adf84bd76049eae5850636175202d03bfb2396d90462a92aa112e903ce807ae8016e1579f3da2ee1008db36211cdfebcbbb15eb8b48bc76b3ea5e54654a32bd6976501c90e32eb3048a96b75f37366f73c75caa11af1b46551ffbc3ed886448e7917711621e73bbb8fc2240a01c5f038dc556cbc326ff7e4c9af3dbcf2a92a00665565dd322268ed59434eede09480bd8d9ba06f133f6dc921803fd51577cfb918afd05aa8caa4c6f9644e8c1d7fbb3fd3b859328308d2541c01ef156c0b37a951b68dfc6ea63e9f193d701bb29af579e315f52b33a2719e4cd72fcc498411761c1eab93c12a5318c2e8f4ab813b6d6b15e985ba3d5fbabe04f700713fa48d270d0b82f4f5458fa1b3788270fef18448c2c110cc38f4b37901f528b19de39091b1a52f59099499d8f7c2fff9924bcea0fe1f3473ac0f7d7b46e6fced21f636b20374bb77b948cf69ed21eb20eb55c1693c83763ea1f5d509e76a68b736bc7a6c712062132033ec54cab2e17d22d04a8eb2da8bba90b59de54636825c3788ade94c75f904b9315b3b5ffe42a7f150796b6ad0455a172d6fce6c4bb21d1b4c5666adfaa5d0a80281b5aabd183f7af36455303cddbd6b522ea64490d6c6dc84dc49fa6cce372757b346e0682bf5586e6507d89a401f23c618d2b2baa543d84ec36f7a6fd96322ff2f43a74caf926dc02575d1508e88ae4f23fd40d1275e3ec066476d4d833dc9d5b1463fcd723a0cf5e4734f25ee2a09a4f3f1bdb08b0690de09d50dacf4dfd3ef3f74662b23511c34b203c8faf5ba6d141a4e3f5a08aa8f457eb4510cdf99b98b841f42aadb036953b8799f0ec4c5617bbfb14735079ca001cf6479b9d1acc84068f998b209cb52c4bb9ce2cc90835cd3122f4393f8f03b9f469320c23ba5368f26e8838b97d6d110d84ceb086dbb8ecbb14ac969b485850c5facc9abd1e90e4a789b54f54cacbd6147a2def5755f2fdb73d7a3a2337576567a394d1ebdd292645e733fd35088b5c3850172827a3037fb500306463ed305150ecbd34be58f25fd9c01cc35f6183328aaf5559cc60e486d8edeeffca7f4219c6e3ddf0dc597abfdf57a7bebd8663cb8dc8dc2b0fe4dc3b5177ccda94416164546436f6e8175ff6a3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h521b5ad8661dd17713e872940ea572869f3396a3f19e6c5d214bb80826998e9242d367ea5a145a9ed608dce21a36a61dfac8b9410be288dfbe3898e8f7b2a4529acb837d4da3a308b1ef26fa7135feac970d9240190f89611d85c1f1f9011d7f7d0ed8bc210da3e3e35e0ee0c83ad1b15c9a97e9561b98ca99ed10804b45bca9910edfd486da43271ca375f34dc22069b94e9341c461e9ee75fcf92e4e0bf44bd0c51b649cb596b52291d0d1b4dcc2f011d28300b4cd91ff463d049413718598b6eacf7653a4d5a224c2ab9370d2e53b171b30a0a573fa5f0fcb9e1009f5960eb44a24092be30cd6e6a9e77780d9626515f12b6fb745a1ef77d2cdac579406fc48b482f6c4f24d916da8ec748d07cf1760257392aefdcc016e9c0be8eb71063f4d8d9612dd553a732552519f81237428e53f1146f565d0e36a66be3901921736382bdee44be99b59cca12d9f7c7d6ce328cd0362153dbdad9417e996b830072b121ab12db7248b2187f44f2e6dd9eae5b3529cf1ba989ff9b640ef62c2158fe6858589cce8b0609666239c9e452533ca58ff714855aa6e64465e29da344c7535f368f03247d4cf4600eb40a002be32d57b9d122fd505e191b4c9d2f0e72936b4753140e3350a077f52d5e8f450417e3b8ea55f070e41e235c2448c7b0fafa85f863040c5c5cd6c8791d06328a2d0cf35ffdd045e2f8fd60ec9868357c2f6a6568591abbbdcfa56a76dbbdb5af3a84cd96eae93d7d09e06a503283a8f40e353d096bda664abf92c98e18e725561986aa63032181b3a1759d9da4d6db8a6ecac67bb4cd188ba0d7f021e46833b9b89cbf677876f89691651b4b0717ba879e75cf974aa4d9cd72f9a83a4ba5040ea4b9047b6be66221736d4df3c0d2c5f8982ce75e6abc9a6ccdac6a6ac7550bb73124e84781d7250b29817f74b50a11259daa81d6bc557de31fdd1a5bdc96e50b68830847c7560dfec6b50f8664ef414a858efd9b408815524bc5b21ba24886cc91295cccc4fefd218b7c7da71fcf8acdea3bc41507123916273a98b4061bcb91d490c34f1911585e3108e80abb7e1c5edbc5ea43913d8f9ba9bebaf2246f7d620d53f75d92a52b8fc67b9631bff4105c8158cb46f550b3302ee95667171825b35cc125673ff72f25f542b017422270c1a7f127c62d501d437e320c8a4ea0925484357cf890e9d3d0dcae3eafd702adf0b6670776fc8dca1c04e35b58ad02c071781fb031064cb18dd6b2234c8b4b41ab35cbe61dc0997d48fa1e17a3464d93c1c6f9ffcd099787d820d0ddc170ea5c408114e18143433e7f62b170cf8be4b90c522ecf70bb737eb03358360bec2859802c40846ab65dbc7128b6507bf3d791d97cb592fdd70e9e2f77775433a48bfbaf5bf70037cd52b2d8ecce932f84287fbe40fa46150410716fd1e915c17e16bf9bfd3062af84bd83acea062083babae6b37c9acdbb0e8d3cc376197a568f92043125955d152dcef0769b1fcc494eaf53625965e05d16e2395f471c00e5f2d6189236c7a7df0bd91cb6c6fade001e0bc14613990915da3e8d5d02b54b4fb001156fb034ee4295269c09b226982139848a2d3bbdd0f4cdd8ef2be5a545cb71f4fcc55f657e20e9e0871c74eff21dc24501384af0747f5da7d32695732a067fdd8c4e9ec898c9c8f7f8dc99ad69e57e0399abf301c0e445112a92953ef77b59429aa31c8adcdeab5e3cd22f7f7155983797231058322aa502a85f653561051f313012595776643733b9b0f90e91f7354e48f495ba915d91c5598b7ed0999432b129e04e2c2b8bd36574255b7b0c64032585cf4b77edb7aa94ce67e3cd4e9f8ac74b36f5a56ef5bfb6d8aca2c837142511e865574fb284c8489e4dd9c0b2c61bafa1898c65ab266cb759d65b21a3fea408807061704ceb43bb7ea5389ada4078dbfb914bad249f00f86524cb6693025206809f3e985efc9c7f343837b7667be94873267b3d2380e174bb7a49db7c08d6bdf78b5c7333a66e9a31c55807ebda13a0f0b3834d1552cda8d86a9feb1d9f982b3b235d8430118ca69b6039c0318c8ef7999369a30f8302eeaa2cd68bf4c38614fa7c32c34599b685cb90b354504049330db6e440d7c57fb41c3256ea884735a939e73eecd64652319d4378d8819434f9da0cb872be859a8f9a5f1a007769ef3aa46cf70f5d60ff836ec6da440a7f71e2086e8c4ea667ee7ba53a48231582712b1ce5de04b2b7d37cc1213329212786fdecaa30750215a68590d577574cedc8fe185488b379986f1d0e3b05306393f542202083a0f93792864f1df7d3dd67fdb36b804ee01c12f29dc75c214eee6c5da646c89a233ad851e13f81e463ed5cd527927d3f16afcac70b18b0af2cad759e09cc1ec8054a7e639e7a2322ae9b270d3a0a15f7c97ae03d7dc909f87ac84292cc4fbe3b2f28d3244816d68831a8de76590ae96ca4b83d6480ae8074a12ae94f69113f3d00b293f5b447571ca7512151417b941e4a8310d230c4f050c2a1ec6fb4363e17142660a7173ab971455622d9f54cdd58783ffbc28841268eb4de0714b859a9bf36fc433b209c37a77072ac43023517255af9f609985c0fe8f0a29c3460a755a80f0075355490158cd034f7282709d1a0de31201f65b290cef02361f4c275710934ec9f851ceacd8c9f161546b3df215743538e6d80aaa4507eb743cb48b8813b9ee7f820b91b81c6bd4a9bc46dff5b3ad9c0dc0c7c2abcdd8bef6513ebeb803476b2a84dcd870c2e464b871a09b0a0c90f31af0ebc606cbcf1eac4cab3dfa1ec251dea9ca66b95f9dabef583cdb66abb5692307d7952b9d439d8914c7b8b6f5d8677ac41b13461a35087f8c7cf49036f966d17eecd5a632d9f328bcd3efc6123f34c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8baf5bfd44b2820a006d4c2c654d13af956c144cf33d758f428cf809ac8fbe2365e6c1c4972dbb2a4527bb5a07a9e1264da9576374e745451b70524b4b881956f223b5da75ba2489cea97bcb93804f7600586fbd4e28689f41474322bc48c65691ebcbeec4b47827fafc6e41347a33f504c194926418786293d559d2a66fb7ad261bfe83c9bb1ed0c5da9fef0663ef586a3a424bca596514e6e2e1292907b1796f74adfbda5f0e07d7e3d79a7349875b5fc901760d8810033f907e686e7457fadf69593d7a5969ea190a6c8f92271212689551094c87c3492f582d3ff2bd26ab1aece8a0029cff5d23377fc2b7dd65ab08ed5c354a4cd7c6694bf5253e38c4d27c9cac57e3b8794022433252a6c1fb06682a753ccc437fd66eaed3dc153bdb525ae45f73dc5a0daa82bf8a23e1ce86e8dff10e7dfda6529fbe308d367acef78d3c51b54998d34e314cff791efa0be67b195eff61d65d5455fd78a41b9f6a9ebe07a16d456c98f086811443b6f7b40ea6b6fec8561c518d0caf5a06b0a6e6843f688c8288f0eee3a04390188569d0ac84d3a231482fdf773a89798108e4e407100ff54cc9f54fd9a83b21d4c190764bc1f43b9732de90de9818b39c375785f3a27c38460c261537e901ba8f3947e4cca77b6184c988fd40fc19bc3e4d35377e2f5678fc31cac07d884ab4bb44e34dabb829702ee240fef06c04044cc778a4f38741c2a82d0657133f4c33f121c01d344e43deb6b77c9fdd80bb2e8442d0d09ce72dfeb47103a5f78bc6c04cd51ba93ac3ab26770567880f3f22d64242775df356ad26a1f29c3c9ec8c32a030ad752c82b8f18a6a7e5e7728cce20fc1454d0580c861eefaf419d10c730d70258f4086bac974cb5803e935a6a7d4ca049c5aedab0f317e727ddb50107bf2dfd31743a3cfd992876e3b207f7fe8290590f0277c5e302961dc7d92187d64c8551abba2b444e04f6a66d26a050e957bb6843a5ac35fdc654f69e1100c0f8d49b5e1253eae332fe1860558c037e866389a6ee00852f4b417138697b7f395a9f3cfcb247f6115806c6c52f67d078c42ea880121e97cb3ef35df08415c29eb934167d3740476708a52d848aa5fa8de3c217a03bf85541a291587669b25589a3e69d6ee24dd2a70e9a4c151afddd14d1fecce9339d11b986e4b10f9c4a04db5466ab1a192e507787c9756247841af61dd63a179a24c82f27f9052d82753f2d5380232b462c9764c7c352c03c3708cb1917e0ecf018a4967088f6594481b446b8646e8b0cde1614bb27f695ada419576f3d572df704b32b122fc80a2e8cbd5c526f29e211ff0954c32e652da20da83cd4a7ffcf8090c3c3dea3009675cbb4b3eecd4b5a19bd05b3086696a6beecb976a9fad6f4e660309abd1527bfcc4328cfceb3682916d164f7af5b6586274be2d323435061c5d84e5e63aa6b97d7f58ebac687f9416616e0e2a136d016e4018d70debe5d29d7e7c10be0c035014ccdb14ac94ba50520016970a6370cb41353cc260305e3c81cc5d8978cfd2aec0179ebde391013646a256aa313e5371d7bf3e6af328ec60be2385b44206b96f3ad4319b5c40ce770d55d1dd13f861c6cc10b096fd3eefa3cc688c6416708dc55385b8ce3bc0370d3b87560992b3252ab543938576760c6e200e6391c8a6bcdb0b8501b225134b56e0a09d9f85c37167f847f39ba8d680a19d234c3eaa14a49a3570b4db9908d678045a4a7eba9487d183fd7e3b9c7aa71a5e8d009161e8fa05cc32d9e4b92032ab35ab0b29ffc280be7f3ffc7edf122d1f11867aac7898e331a0f27b16785b3ec7f5ea389790288aeba48307f25c7cfaf5f83980a166d4e9c4d0cd28e40837b8d74866dbacb126c15ef2960a9d54a11a800e5b03d8daa2e9dd0630e344b1f3866ee24a788cb727ee6450e057cbeaa38efc3e52472d05fcc018470adbe81a0956eb5562c994603264030ef6a4145c543a33740bdda7cd73a2f188e6a168c404b3777f50009e54b0f5a08c78b63a8b321e9f5a1adbbc78e21cd61fa394e334cc213ccd1356d77887a7ec302da3900ae8edd7a9e77c5440885fa74db0228573704249c45514bdce09bb5ab0c08281f97eab552cbcc4d66724733e2ed19841ecfabc842fd9ce29c2764f8c0fd1b20cc34b14f74e0221f249b51c8320cf902fb3d52e0456acdd94335936a0263b36851d2fc5e0c10c9fb25e1e44be68bb841306c9b18ab2ec0615f313c310f8062810ee0f1fff4d768be5f14947005a45ddef57834fc89857d8c9ce49391119a6f2b0095101c7d7f2e5e23494ed5c405ad62713f7081ba7094eb81521453f3e392907a0eda20ad187a7cd4b074a7c031573287a324d65ffff5fee28b5cfc44a047e100335629200e48ad99aa130a1f2e052bb5bc84405f2c0434adcc3ad53442cc60557774db15b826905280d61d66093637bf226d38da7409a9a0f0f8f5f62827f317883a43e896cc6d86606d33c565b677b7afd932f923c47523925e8bb82b0841e9e447428f06f5344e2ce30261285536752eb7309370aed63c77d3256c9da557f1dcf88cbd3de0042d93f55d641238d9d8e6f28b4ef6d1f72b45c29e88e0d19824d580dd5378f6628e0ab1f47f40dc77a832be55ba2e1c9a3d5117e2141160010c9b0f9f9c546bd1537e131f23ec386ee5d2565822c019b40b431c9b36c7e79953725ddf259b1c72a58be0de365e4a09e018e3ed0cb48469844f329b1565d77e2e53253baddc21022b468bf0a1c18a34f475ca6bf32eb199d81888259cd361d588e28d8483fbf40393742271c22a9a509ff71ad5cb7bd8e48a427bb2326be403aa000f6a24d5b80f65016bb93fe90de1a06be5ea2f2bfc83a888fe1ec76ed54cecca3f4d0cde25e0cdf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1ec88cd0382c9de3bf8685a4c11dfcdf981a3b0867904111a78131c9bf8debaac597aa8ff71adcc324065898ec7280d27a9ce6ca7fe435333ebddd6cab937315dd9ea636a60b43ff3d96c6c264825adebc3e27a8019995ece717925e721fab8debeeb9f8b77bf083c589b4381c63365f39e7eea7422be6f52109fe4bda215369697cff04adff50ff730f4dc9e74916b20d5c67da82ff37ee5fcb54b744b174e735cbc6eb912ee9dcbbd8481a017f32d52fcc45562d9a44388a33bc2d9fb482f024a55b35fa5e38dad0dab47debc71bb53112f0a4405097551597ce6b048717c1fa243abd55f19741d366cad3866b4d7f57bbd84ada90ad66ea351d6e2e9a8d096ff4164d97177eb27a7986058708a32787a89f461608e636aee58483c5762369af4e89a9303dcc305e335b43be2c6015f9b5b878992f88fbf91a505d3c3957088cf2a2e92f7831b18419953fed279f08bef3680ee19a04faabdb5e23527acd995327c4e2e1f63143701e7d4a671f1aa42f7f3d04961c456a44dfa0577cae078fb3dbf871fd379194e263c91617978ab47c6a592bd97480293e84b4176f73c423ee8135dbece371cdc24cd1e2fbe4bade44445e5ce123cf997c241b9d4dbe0a72cacef724bdb5771273ddf3933ebaea418ae88531acc5fe8fb848e56b2658b55ca397ed204ab229310470fa248a5e355b929a738f58c9e44abf371b30f6d830cb35db9ba61daa273865fd07e3840c28efb7cd7b7573fa94fcfdcd58568f4def89d134d3bf65aa40ba29a7cf80568019efb32d08dbfde0c0ac4a26b1833f0e63a8c2c2e54e521824c5c0574bc1f9e90864c58996a484e76b3f19519246a241bef31158b00961b840527ae17294766d51ff20b7254c82521e129372f69476781867735c20afdaf5167b013b0adf73909dbcefc7723b73c3e9aa35a7aa39b0678ec199aa7c1e8377dcc99cc896ef261a39b808ec4b6ff4b20c633a6d88b3d5851f13065be007cfeb9f1ec1285d1c5fc169df0e8cd34f06664514fa48d598cdcd7ea85f566ba62e93cb38ba30f08111ec268f32502a2c2803ffe93f8ac800556717f32d5cec96ba5eece7d438743de43409f954d80f5487e5e48d4ff19321e18dc99a1ae408ffed909d5fd82606aa7e60477b548fdf0bcbe5e3011a09f55ac2bb92708850b936964187cbfe360f2ae7d4aed54726b6337f65d08b0ec8b628b08d54d544b517778d3932f176c7c39e7ac040892fdf33d854fc214bc93c88e212a84a48a9dfd77ba35b5f892334228f87b04e2511874bbaf45e8bb183c4f620a4bc3ac948fc8c6366aa061085ac4224b5003f1005fd899b4828eb65bb4e47d1729246974c505be1ec5a9475b8731d1f7cf07bb5c4c33a5682ef2d064ee758a4e44de06e344569c4fa41a2c530f8c321a30dd52d10d21e42e54766f2162e3eac281daa45700ce36fe4ca97e6bea4fd176e2c19b2b2c2c28e94feda3b6513cba09ee1596517cc0580b042b4a48e872075b2b0c24564d717bf1f77d7130b370c30d80d276e8df900ae5b954e33854143895f61fdb1e043a53166a7b001987fc159be643de16a2e83ccfc9e7206fea048f024744cee71e32ae87be13411cfcd21e29872e2a8a7a09295d5e42958104843ab44028b416b594e48b09f521d89da440f037c18975f9e7f111af18ef106417e6b3e2880878bf829b9ab7055c88e84a23b8d5eabffdd1fc0411a287271b8d8fce8fbf53388b9d314894ad8a4bbdb24dffd1efcb491fd51440a4306ce8fc9d76aa1b9f236826c13a61c314375785f32cd7b5a5a860adc8d7781eb649389f74a55781e3e07f5911963dc05a65eba1c2c3d4c2e6e394d4e161fb9fbb35b2aac1eaacb63f3895c23d700e07200e030001fbd70fec1fcca6fcf5f8a668dfd02f030666dec3ad22994a88e489a32756e4ee554d53e5f93be103ca76a89d32234e6735033e5cf11c53412fbd019e8c5fa608bdbcaf584002cda1cb1306a40431b5e5ad1172be9eda79849ef7a1ee036366c3109888f930e9c7d43a868eaabd661e0f2fce15a2828f4d33c5c9656aefc5d255281ffc642ee14a083d3cfe8d0a7c42b99ac0a471a13d21bb5af1b64af57a06e2a2a146ecddeaa7cb318c5215e70308927bf71f84a8be5f8537e2ff1bdd5ee993a5305d5ec9863590ebc165962d854541e1f77602caf1f738b0eee4f1526b385e3a62e116848e4d75ef9b7490665961b597c77d715257d78ebb7583c11b8023da177349f1ea056bd4281abab323fcf8e37dda33d4d0c0e01d1a9135c3f984c5e71d9478379531e2687556642755025c3aa8239638e5e981541570b001ba878464cf49b19b440341b55ce5f9b45e52c1535c88ab2f96b66f3c73851d5df8cd0bdb6b3d405840ab45d5435b461eb4c25a9a28463feb3ae03ce102e0c4b9df57713f136c75456afdeb467208a4de97e37810b24ba80ad381fd3b8b5d164a3360d7f4d43be6fa01b7e438eac32ae5b1003a59e714f644cb2525c7ffb75560e143199f69bbe89a206af0ad6e3bde933ebdc3dd00102831a96161dccf48b8824933cd8c9006a52ee208ce2d6a9b21dcda370cab5bdf066380fa7a79e176b413e0a80272f373578b8e191a929f37b9b1d4e62909d1f3d5f01e1f5c90007315ec381e8fba2a5179600165b455b7707102d3f0e92d1ce3304bf2e2117f13ab8b36f28aae1a3578d43efc4032f0b318125e48ffb25721de70df60d6ea3b1cbdf519f163294c9b21f8f1371f6fcfb7050868443949430205f593df59e3715c0ef5cae0806cdc96976d621b259451739947ed76c1672bb51d6efd7a54fcede7c8dfa1d04a52457777d252894f21736629667bb875daf5cb821964a52e37338cedbee6d896420450728c28718e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfb372afcab2a524ce12f3f494746350094aafdce9fc5086c27684133fe87a6d70d50bc56b5129c9740591ad45c246b4f629f9802a84d1169d1579dfa5116e81a11dc01fd7e43971cfe2dc7c8891fb062536f96ea79a6773097c1364cfa66e7c301227d8b72d6286969c1a1b51c73b106456829e8a2a9c59e286bac6d54d0fe32b9bc7befaac74db61fed6df8190e911f1a7d23d891ef77e35de7561f13503dfdcc3fd1e8bd44455f7ec66cbaf5a01be036cc56be4cc0fa5f3239ecd75e1651052ec1002b3c1426273a744110ab39a64385c9facd88399e4d130254064483cb9b3b628bc5be01807ac5a68fc2de53cbcd5fb3c6e0511ed7fa93779e672562e3c5d9cfcfd397e542fedc186660506acdf15cabf72c085ce3bdaa36dc9c70ae78e35da484fa923449caa9fd6e8ab42131b3d54d0d9e05d403651cd7b9b2efd880698723138dd70a55e609669456fdb9be4c5598c4386dfbf9426f3fbadabaaa78fe6b71732b6df03e0c8588d3377d6d3e50ee51120447e9c19c4bc24868ea7708e568084759b07a35c84b35264459a1c00aea1e185109bff065f39504d977d67f18f92897d369d8f4718d29e153f89147929c258bca3b1a56b9495c502e23b2c3b22fd854695606dbc5905d3750b2aee30c6f0ea9850fec15796b6b678020d79e01a96fe93937e03dcf9b580c4ae62b69211ef4000a6a9d3deb5dee5af3306d3718de57c87b5dfdb5d8315324496e05f0729e8e14b83a65606d5deac9fab94ce4b0034147258cb7fd02d8ba1f056a897bf62fd758e45b291e7f43f2727aeefd36fd97f40ef35777727d4d62cf200d692c42ddb3cee702de3b3963dcc4925b1de0a9b2538051c143883ee196b990c49d2aef329ae50ae049dfe38f854994a3aae25d87d3fcaf7b58ae2a03110c474f9def6a4a3368c482f07ec4a26afdf80f4d626eecf6ad567d76efc73ff36c7a1125160d3e1529a07daf65ead5e13e37c02e42bd7f9561277fda26f1fb5efb2231a556f01c47bfacf84674a6a058da7101f50cd9b26be5f4c9f5eb0a7e8dfedb01be429aa0ebb3d133913e56e18041e10845efd72fb29ea115daaacb150459056fb353cc7059cbef800ae8d8c0404bf1b1912c66a6de9aa4707f6ca544bb712ee9877b0a5fc362f144eb2064186d2e33fecd88a9ef5d4c3840083eab15776bded74df4393243066a8200a9e374d914ac63a99e0637a2eef0cdab148abaa392e152a6ba120c69f8af0a449978c0d7e554d92973727bc6c865a8ff56ae74ae4f0e6887fc13ee622ad00f02f68086db9498497f6409a5412dfab3cba2579aa83883c1c543c61cfb0d417803a7607f45ee504a91a39dc1db71ea95051a7382d1ec9e5ce2958c05af2750ae542cbe0706974ddc31ca3a829b3409594e8f2c9471b8c712cda3a27c06d9701e886657c108deb07f2b9dcc41bacabd7cf92f41a5b81dcbb4476994648270d205417c2c0ac56845f46e05ff48c10a6eb3ed1ab755f888d4aa6cd3bcf41ca4f8651705a1affcf920c5a7d572bbe578a444f81f97aa53879ed25f93619293867356d45804c3321da2ee6db4651eddaf58e79c680d6601b85f421d123220a642bf6a734144935f23840c4d0af88bd6f4d77f16d4d5c67d672c6e4efc6e07fe3a081d3637ea8c93c0f4b7ff7b9b5168b66e59ee64559dbbb5e98ef2852a49ac8d01ba07bdc4de7a3b221a767016ca1f1ced0ccb82e9da492fb9ceb9cfd33b49c723164f657551b53d3eb35f649972430e9f5e19a322eef2071bb91b47d63d228e8454b1f1da3c46848e5faa2eeba1a3ccbf0aa0606d3589abe63c9f0ad9ba6506e93e773e05c1fd03f008ec317eb1e208abda4df49b261ad8429118b392b1f9438265374cf90b68be73583aa953fae3b0d23bf72c1ae65e20ba2ed2d5741230d5396901b681c0ce31fb444173bed69191cbf6c9668cd129d0ad0f0e6ac060508d19a40159b261882b9414f497a4381934622d946ed6e21206f0ed22b0a7377aaea0ca4c23b4974d3418786fd44127ba8057044003a3df9c369a7d2a4d38a929b0d22b3a518674015277e95bbe41e9ecb5b9145c772ae8acd078723843d30419a607bcc800b5040c99387a3376914943d1cb7642bb6abdd1e79836c4a44f5a0404c13524b04565bcb6b434f3c53345944ce90683195932d81fe661788a7243d084b721d9e11d2e386ee8a1302261d5fd733a1d66a1a2078cdc8af9afdf6a02d7305aa21776601be85a6e3059459f2c76daece1a48c6e3ffcf07dcf6fe051e36e4e86ceb1d6a735daa4f659c8141a15fd32a842996d0ebaf344ccf502fb521149c101d3a5dc6aaa624842d5b54dbb8eb637d921b8d0c5f0eaab7624336d456c780dbec272d6db23d36669f378b7c8bf70c9b59a06dd5e49cc68374dec4cbbfbf78b199e44afbe6968f0dfd9100f66a872fff4fc5558f80efe4031b984ec5ceeb0784b80c6132a14d9c474ab9be98087d3b42a27ae1275b3130448fde7f0825d691c5122b06ab2b10194d19e6038825b252df0fd3c9e2dab2f3dabdf364222c47c25facdcdff2a12d118968f7027e400fce82c137a6988d611c7ea96bd0efa85c19cc8c918d1d4e33b0e109531d224ba8cfb511f5e6d75306dbce2a2892583ccdc63e31c92c515dbb0d85d468581d35a8d9766231822feb838aa7f9c2d4eaf449e97ad6fe3c4f65bd582082d756f4b4944a4527998f0f8f2b3b7d1d5d1a332d6c4de456fb55e36d5a6965d5ac0407de24141e63340cf5f7f5455fd7eb6aff5a4af99ab5401531e469738382db6c5474368de4c16115b8629f48faf7c2fd67ad72029ed866becfa7e5dde67c88d5c8509e751427b76bbb52aa2426d185eed9a43d09f88c514eeaa836b4c44b230d30a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6319f357787ba41d4772e0f71c6e65c667dbd30939a9f8e3bcfb9e96683cf7c22aa085ae27e37abc3824f6c7e2302f0dfe8a44f73e2c7143338b520992926f140496c5362da1afdc758760eba1eb21903985900bb9096d91fd9c891219da13705819174d19014a6d0feefe41a29725ad2e3668444849ae72f47a0e1e9d4ebf60ca0bab62fb328b1573167dfde62c63132167132425985f30c3b53a535db53cee28914172cf5261f7875e8c6313ff41fe4d4d99c74aafa0f71b183e0470fba4a4c0b58c48005259fb2b0514fca45ecf16343b8b4bff9f2628ae0c7300e83f2850518ec083bd1b3592ad9d06c7f144d8b44718d1735da2bc60685e71581a39f2468875858d03853e4bd6ef635eafa18f9741517a16d208f16378a8d85e032e643513b4ba5be80353087e0238d681ed133effc2cb64cc9e992bb6003b492128f39ce2c2271e9f25f536d84e78acbb2a0e9433cb4a50e356b946d39e1ae6119db5c55a4993dc90111670d456d3d528ccf55d0b8689f67ab0444adcc63bf29f05c7fc0484ce7fa1004e03ac4639067f4ee91714ee66cfd955551670a0c882f11ee4b1e376831b4ff8fd4f74bcf8647f0859c49917ba98aea5255b2cd5da2d251c66d076ebda1b491b8e76cab897696278c5ffae394c421417a26400af86b0a35d4d564c1a9282be2f8b1e08b92b469c7ba1ee3380b0e4f4b1ddda3fcc1db45d4fe977158245ec6e0b45b469d40b330256a83dee1770d833904b9bc364c93eadd2efd3b3e82b433e71e1a2cfc01413172abd99af108b133e58f7b84a01444599f7d8b0852ebaede6c03158cf61725c7d4528a50ee528e101fa842eb64c00ba504d271154ef145a4302e62ee1325bbd42b9bb080a9ae187fdf15481d048a80ad243fde14b2123e3d4336bdd78c0230bf18e0c73873ca2bf69a4a0cb480ec167bc38479d4566f256c411b47f1b78c5bd7dfc7998bdeb474886e78b60b6a952ee15081bc8c5732f4bd7216fc1c1d8ef793f9ce74255fe56cb03ee29455e7254e9f180337c7864fa4eb4b7dab4f49375bf40e7331078c041dba4a4f9c2403f6f37692ff55023cd3eb42f8a236a11c414e38fbef38783949f755ae0c149ab683d04152b8ceb9b247eae960b47360bb1614be4618f77c6597ed9b7bd24ccdae50cc45f9c2caa42d7afda45f8ecc54571355f4c91a0ce5705ae35a8397cd6f34e9b33d93afb7f1512611608a345dde5e440c3f9ed07790fa2f85871e3a2dbe133b8f9cb2c7ee4ff30692220fc609ce6f1a71d37572eb4709e7abd1ed533db6c25b39d26aa249e8e68e11b08f9bb4cd908af0d4c0977c91029c0ff8aed9b991aeb446edf56019a1a9bb1c83b4597fd2a7e40202b448ac9d1322846fcb59a1d7dba2fb4fd7bf528d7a6e07b11e0c3c26f4de1aabcd63426607ef35baba0d41c5a15af6cb78e6cc85b805eaa7fe2ddd4815a6a9c7cce6b3004b4e7d097240775ac236cbca8538497800be95a93cfc8f96dde6b4d937a1e51c8df50ac95e2031dea9713d221394317106c477e2d82cf5d54901f38169a74ccc699f5a92446b028e4b07791bcf1a3eb9deeddb867418665235f82ef3530737a487b01b94d654f543716aa98903763f4bcfdb77a2cd8365ed31727c0f33c35329172d9da171c450b8954311e60ac08138f97f1948d02b841b484ce34d5d0d40eaae7c3012b7eaaab1ecb2cafb2ab41a2c21a232344133f60d668adbe7bdecdae30a4e12fd6466b1ebdafbcfb80a01e2eba7b0339912a108445b67ad358eadc0d6d9be517b5547d52c1c4a328074c02683722c0488d43c11c9ce7d1db728f11279be2d025ee7334c0f29ca2052de7acd5fa03562b08bbbe52ea9ae79f376e8cfb57d18931f2a162d7cf5d3db17b08ba84f55c20c0d2c107f9b6da16149b778717d0f6f1ac71470d17b6691e23d0bd79d86c2fb0ce7e5989bc5c4111cc82ad7656d3ceda61b23053e8110d57296f742112c4fa0372c8782ca9be658c6a60afbed3205aeea139b5bdd8459689f54c6ed33f0a387b04d8dbef86b0f79ce7bd3739087974dd83693f5c711248d2d1aae6323912a66b366bcda4f088c179aba7acd6f36edae46a6e9ce8e6d39133073f06c567c55799dea6b4d0178e8e3239241719b523e3ddfe80fb010fab217cdffd201015b5c38d72335c3e6b4eba753d36285fc250a21118e33e87291309a48d9de6dc5686593da2c8b0b82679b232320f85f2416f0bd1463275f8d69d3b8a32eb508c2a9684d3a17a694382a69e11667dd61fe32efa242b8f3f77441185ea5e76696a038e7f35f18e92aeb504a9b0d9fa1836d02718b61b6de6329ab9e7833673567efa2b8e924c5b79ee3573f1822ad609ae4e4a8c3af127640db9fb52f66e7f027346883a0799780f1018cf9c46a3c1afa5e4fcf2da6165c94f4906d0a6df785d76a3fa10853b2ef8a9791d4c7d034284dc2bda5214391c39ca560f64533764b143115057145588392f71cbb00359d228f965c0a01a63cb82a7a67f844c98b8514e6458bae8241058b88a7bfefbcbe4ff1cda1735f1d5af9c7c2adc6699ccec5d9a739a63360c4a81ace6f7a50f4a9bbda5b074638480972273dd8166bf562e58880d1b1601ccc537d57265ee6d319079c240299e703bb9696bafa7fbf71251e4349b6faa520ffbccf00ed88ffb964396bdd8a6b34cb4cf4fb87e8e46276b3953894bba9bed7a358c795e5222bd3bcdb2802eaab65fbc33a64ae9a3ed388ef31026f64e66f3b383448bcd4c3784e5a832c7a05f444e85783391d982200c33f61d8c472ecd68d31585290e6ad8c90c7f24e855388d4a42de3d34a1243ca0b257e39618547d2d0efb9161c719bd7dc3982d3717371177a1501bd8e732f3e2146b908917;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h73b23cfc3e0d88f5d465b98d6efcd858362e5f4301629a9750d0b807e43aa1a5d0ad3b92954f42f9d9fe7c59451fb91bf0eaf89516267926a29f1f5535838f62d485299a2dc063e68027e52427ee366cf4417d9ba458265b2958b07f9803cbf7846639a1523ed1cec3aad2c7035da61f8b7e767c02ad9019b0ae10d19daf2678f36cd0bdd6d5be36792a8eea4eda22cf6d710551631e68015dd1c5a5c50689dea6b32bc5d57ea46defcdb27d95f98dcfb99b25c950605eeeadef8805220d6f566026b8d63e6ea36900000bac0fec4677851a881bd744815c380ad740faed3bea0c3f8b165d14285f38005b4ce6f47d5a86fd482884c771177fb0a35773546c06765b3a789f7760d918dbb1b2e9e86ab21e94056a80cbaa7841f561e34d7483e0596f16a1e1c375652711c17d6945be29bf98b2a7fcfbc94e929342ac1f1c79c6e5f1b8cfbedd252d8a72219f0ef9e351e2b29731c1792044ad290a493b3dd8fc8f514216632d19b05c8911e528e8dd272733c3db2447a1abcd4226f5233b3ab40ec8b539c5d07e0493ba3a96aa249e9d390789467502d53fea3d5f2a23de8d2fb8d34ce71bd66175137e7092085b652cb871e9c450e856b32eaa85028b30d9d46727631bf20c81048d10e85e4a2404f47096bb47291a8c3c06e87b20eb2001c9ad1b6aee08a17625aab60b0ad95f6c7b62f1c0723a4c01dde15fb356a9c162ae47394ad38d6a30259a54f3bac2f2f6fbb6dd46d3b0f299103ea3cfd04c4dd1e43dd926e0f30dac621dd41c7df7b3db93111e4e1b07bbcdac02faa20deb4b7fad39951c1cac4e555edaa16fc70ad6b1253c8adefaef1a72bd2ed24e3475e2d2a40c1e52fc2131b5b323b392e2c12c703adcadf75fcef9f2fa0dc3e8d9c46f44644150359bdc1a371d392945c9a15446bd527fe77e5fa75e4030dbe54e00a214616ed72d41da1fe0e2512adbf2eccffa7a941a5b53088c4a2b11b7d96fba1c8fedfd525cf7321f153c1c57f9fa49d2ae271f74b22872358258c6ae0478dfe8949db7fdd79548a901002ef6ea322530a2a8f4c66f0ed29d374b6bd0dd37f1ad9b0d15d7a70eef3d346887f596aa5b5233b1631678557b712653d0a57263c7f9c9b28a641f7225851c14e21a344c2a8d941c011db92617cf6c647d8eb4ac7217d2f755f9057c2d3e5785e9b5d4ecc7e4116964905ff0c562d9e5a885e1450b868ee094f5e74804972c70795060d16a0334810702a924cdb83c4d9138e2a99babd345d6ee85ffd58daa070b776cf6bb7b770bba6b0eaea517db08f548e9e4a13b79a5e1eb610c1e7abc02371eebd5c03ef83b0546413233f5b250478d6eb56a23c7da568f96748aeb9f03750187f0923200d48ddcbdf371d80d54bbab66afc175fcbc147ea34fa5d443b282194647958718ea689961bd43ed6803901a78517069d6c14eceebe8f56b440bccf847ba185550514dbd76ca0d6eb7a80917da013ae0d1773a81989ca9ad391667c0220e7a10b7707a8783db382a7f744f262cc669b67c7a086ff4be2e956442a8caa5599a24cc5a8076c15e365f232792d40f58bdbb2127240fa18690b8e0d4966d551b5789ad49b0e9f6e0325a499dd71f1a146329682c55dfbaabae9b2f8433a9bd15628304a5058169a11522cd4e107ad992e08ce1e26d89397318a73b6d5deb2bd1dedb6bb6419bcab41c4688435f8a0c16f9b0d6e9621017205281059d411e1ef342efb7ddf3a4a53e4acdbb53478ec548ab24a99d9816462bd4fd2ff4d2c60073759802cb22ad50090d58106217df9bf94c922120430e5a8ebeb23927d8bfe804ce3af032cf0d10557db5722b308e8a2ac3e7053fd8858a62f3a8f9b50679ce6360e4511a04e56c610b2b502ee0bfa1af0f72411054548b9d02fd9fcfba030209433ba70646d1a3e4c17e3cfb02282a6602e460cb45297ec0c8dc8a29ce945e5a4116a0a7caecc865850db4ade84de006a606cc28db389b25a75e5dec52ddc878d6e1facfb410149cb4f87a26ea73794d74155efe89e30611ee67202d9f3b7ba16e6fcba9c64f59896d5cdb5f0e0feaa15d014929179175a61476830c3d9c08625f0254443ddeec2695ac9de84c011dcf1c5a1662dcbd64952895219bd8d210ff04354b6538da6448219ff78c0331b638dc0116a04ba7cf2a4bcf999e5c0f480ed4ccf987b088fdd5d8162574d8afc2d440af368d233221507e61e06e13a8f536e62ff0288b282704cf0791d838684dc9961b92cff7d4922fe9f4f2252532f2293af39eb812b8e2a92085dee5e9b4c08a6ff193828e1331a68b4bdd0b64d87e7e8d0fa04c38f3190a8c06c2bfc40bb726af36b8716796e37dbdbaa53889201d5d58b291d0f66d11f11059f3d340476e0f1b0923402c3a2e6d0a13a684bb21f803d9b07306d401ebbf92ccf76a4d76734c4a21f3b6c6c2c5b55ae57e0eabfced4e49273fa7766bd90453a6fca87e6b0a657b239bedce963cda0a7e729c42304e23ffe19a5cbcfdb8bcb43c3a56506e2c6d86e98b825930c4b675db04b338b4697d290b24b52e68d75d53be31cf2103b87174639d34c87460351030237b58c64bb0a96473faa2ccbd5d8d1594bc12edda53645bef1bfe9637364c3bead878b7708460596af4ba329f92fc6a78c5f3691a19c935f4b9a9840176cfc4d06622a250d3a623e79078c5c8ad6b67205df2fb54a4b436ba7b2c781ccd56e55d81d22350cc4b82b15a5835965550c3c7f2cb5e4e1b79ab92c29b117cf2b2622b7b461912e06d29564730ed5395c8a9dd51c20c892ab1a30816030200af86b960ebd757af1a3725a0ee321a018fd05cbeb48bbffc626bdfcc3df45b2a82de0152f5faff1685d065a8320d3706a9444ee289c92c1a2cf4603124;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8dc7ba29c8216cce747e2d8df32dd66184b5388191e32408759f8ace8777f69fb0fa64edb5ae9a7c26cd9fb4c9c1cca4c10da5b6beb9bfa6f2218cb410954d627c26b981a97627d746f14d7f5a0fcfeea39f19fc9d9a245374dfeab6e44fb4f589cea145dae3d850d5de16bddf0d791f272c99f985bdd810c867f2ff87097858fe95e87971a8ea3a97140df11fa070d075049d87d31e651874e27b9bf05af96d6c1097ae67fd7435d4e2d30a279f411f698f3f12ead7cf6c8916ef2aca349dc424635524243b61180912b5ddccdb4e14cf335a2a75dad6fd0edba52af0da56a6b3004189df0e914adddf3d87bff9aefba3b68442d275888da7549ef579ce4bd2fa10af2f8e848355afbb03566b7987b9ef63b5ee1860426438a0ad38eca9717731a69543d2f99dd273e60e40c7b2ff10aca46fe78708020f04d1cbeb25ec3d03feda537119684c8a694ff1eed378b98962130c45356e3e0b4e86536074f76b213b06ffd6c1a11a116e7f268ce6e4c0ba74c748b2ee83a89e340b2594b3a998aee18820519ac62041d64d3fb3d736ee8eaa58dd8def4c8463f6b428a4c9213a864c7928d273622a3834bb0d53c5532c2917603d8dc46b8c4d02a4f14bdfd7714d80c733adf54030ad8359e61e382aba4beda5147fbaa8a35d4cd403dea2fda85a38f4a2f2de0c158d4eb6f654d259cd88ad829c517c0f16e99f0fb5bc5d57164caa1716c6fafb4a1df9b2bb0b40689f73f10a33696cc7834c462705c9b13e541ddc8db57363ac902e8120fa6d0f0f689db87eeeae7067a4db5faacd7aae3a5b46bcd78cd8b4c35ebc43a1b36b8ec38bffcfd9b0ae2bbeb96c4f40d10b3e9723908dae2dc22124fbf8bdc91cd0991ea265fce24e03bf3ed9901b0a7a1d20080684fa888c311fdc7d77f706201148e22d55e5b2f941d87ecdfd44a7ad974bef55f85b3302405c5cb6467efcd7701d1dd89afcf107b666c4fe8498b637ea501780a22ae9fe61d0da329ed49e69d49e8b1dfc89022bcd49a0678991dfbfe66e96814e36c10b3b08635d1bf2df598f144e0f6565b7d46d6a976eee44516c46eef70a28c9b0643a85a56b499f5755b5cb8302dd6e0aa38587259092c9ddab592846a7be5b679d2226ce30fcb93f95b354d7892431763955dbd73a75a1c093f81472f087ef8108ec8e0770af8ef9849870974f178b3f7d52512d697915edccd78094d2737b114cef68a81b31f9f04b71910101693d1f80e13674132898c686946fe080a6fb0b3cd9d611b9adc5983d7c4a08e48e8f1891c50703b8bbc8ff12df4ad4ff5dc473d25b2e349715dc1ebff89777a18a2f2cc11c2b7781472c07bbda6fb7d70bd585017f678da171f2f823de44a4c72899666f75536280d56567b44b0ad430f9b4027cd64fa208dbbb0065f98f235cc29d07e05b9cda20fe358383ac1ac4db07151ee78e63e03d79a5b9531c4bbb4de26bc833dd3f5547d43293a0b3201f5db6bbe142ef7fb4b0ebb911b342cfd1fd9e5d14bd283e199d89ffdf2179402a2cb56fda271e38753e487de6d4dbdc18d6aee2c197d9f6441c66d99dbac10e425a3e4ccd0285eeebe9df422443c409dbc7832e504230e90196ca73c09aceeda59c1a0aba2e5a3ed6b2ffd40591ed3eaee54833eaa43bd17db0bff907b672349365a5d3e0cf242a887b41f72b78f4a11dff44c974b342af62dcd484a62ec0b9998ee62683069f3877c01d8e043a4649fd98d040dfd0d4f3503a94ae12bd89d0948e8f2a565237ce3eb24f4324fb52cf0c7171e66efec40e2778af61acc3db9b3045aad41db1ef52bf98c940b15563561bdcdb85a4096952664371c84bf7b4a80fff5147829a18304eda39f70f4c13589f4410f6136d24b7ecf1fc6587e7f670f31a6b78f0142bd6bea93f58513ffdc002592fd74c8b3987107b678650d62e9d4b42d858aa627771fb44c658408bda121def936569cb6153940027c96c26c26ff1db44b03899b7126c8e1589a6f56685192267c88b29e16f380a82e99327919894c856e652a7c5fa4591da0105ed4b5adb0184990c50b66424514dc9967d98ff425c41ffd98c78ff0fc917e07d1de22b15b2c390a9a60b9db7194aa96f9fb5b584b57bd212e86c00af3962c37b8f1b2d012d82c20ffd1527acfc57df4a924757ead1f7b321f36d3738366509c069c9f6c0f1644e5daa9596371f06074405c637ba27ffa9a5656ba17c948020e92128357255664813043188e7eabd609a4c4f2eefab7129d5ec9c64130467aafafc5c4f1ff17c19b0547ea179030a0d06b38ea59ba5d43f7ad57d68baf0d68f6b09fb34e0d13caea09d423290099d4401019d45a84aff8060fa53af5a8f6dda3214301fca215ecaf9d8d5196c1ae97b411e7ad832a4516924f46876df48fb13a5d0fffe70d6f25c713af9ebedb89033c30d44dfe5281069af853436f432e4184c625bf58dc0e8a6cf629f70f5af7df82666bef082a4686b2abe6ff581d5ce348acd1edb79d2f82eaae1d253c08f1caf27ccc6c43c04179adba11b39aa4c631a43d8f53fcea1280c019f4f963f939873587962b02cdd452991cdb2c52c09ca104f13e0d15cfb661085614910e85b802876d7c5538e604224bb370ce0a11555edf791a5dd131e59da16b48351b1d070dfcff72f695bacdd2fead0c54359c5084d2b9bc30518707119dce079ac61ca55e0307295c85162f9548623391f7a399fd4c55dcad47cbe8e956a97af7c29cdd9163c3dcbac88b5860aeadf3089d88b89881cfe7e3f1d203ef78312154dbc9e7d66e42f8c8a0a5e03d98ecc11e1650e68c9a87ca946c81e69d2d229780c70a3d6fed3b7a33d456efe34b2b2c82984b3fc7742e4cfa447df18a9da9789a90208c33b3b9c09be16be86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h79d0c0868c94c621b127564f61d18b3c1d3f4bdf36dd88a8284dc76e7f8a5da35c9697c3650b8a02f3f0b35091300d9bbb7c31eba718d91a9880a20fdb6fa46682ba9703d40139b35f5de29bd9a58d84b5c8c33097537454434342a8a62fe2b659bf5a0e9b1ca4c8ce3256fca22125429c2b4d8db6bbaeb5484f616749d5d6672984ac5d68fc2801ff643c8d61a7e2e0ffabcd2f0e04c7edb94348c0dde7475c2c489b34722911a6f9af25408a48f1f3cd8ca059d96759432c0164d71047c0db07e5735b2d68adbf58fc6b9d0094b5149bf7fdbbdca1d40b1a22abbf9d1585b81957017308471b6ee5b6ef7801f0f08087ddb18496d9735f79871b886edf5fd059a424a04ac9e75dfa17fdba0b31ec556c6d42d28e7f87809f087dcd72b24da91e16850039863887c3a31a04a4b8e71d4f3540b83b8be516442f6e8466175c4a820ae71d35d831658c89fdcaac407cfb4ccab9b1cb2d0622b9b257b132bd3913478409872e40f1975388e7a447a29b2c9e06121f0f478e4867b8724399243b02a344451e4d054db8c8976e84114f380113cc58306d7184e6414469fcc2213d5085c9ca3ab9018afc823618f338765f9b426b0d63535b8de0a0d2335e974eb7bd507875ba257a3aa929189f6fe70eea49a023ef8d66691a7bca50b76db8569b5dbe8a43b40229af2540b857cb4a0565c1bf37399cfcfc61ce72e6ee210a18f0ea1bf8665fcd77284bdfab39dc3e4e2c417ba1bd369ce56ef7b06f5d69eae5e836c039300594a4f71d604db4f883a5eed4dd935e61f7fbd1ba47adc7d7400f602a10d070a1dcf430b9ccd30f49b0183ea1820dfd1a59271e88ff1f5a75f6f0734bd576a0b7d49455cd772478124a8aaab70361cc681be26a723bf3e1069129c9678296e639b838619ef9cf96e178dacbcdb4a38cdf4b3bc7a6add7f6bf91a29dd602f364bf9e926a76765d3fd87d5f9167d0de009bb3be99418defc28cc56b2bd2e8351d210112ac2b8dd7625bbcdb1b2d67490008c44cfd38eea0df43cf683242032893f145de067ebb4bfb2bf6606ad2895249535fcaca501e86368d8a15cc5697245f00e58a0c4e9d438f800c40239ac4470ff38abefb44de230c93749297659bd5b21f2a22db651b663fda17ea87b680f9b0b18407b90697fca01e031d8df5356358b6bc50eca869a312caedf7546dd77bcd5bea4000b1a9b9b95bd91c8c524c1e564aeb7bd0967ae5ae3587f3ba257da3921fe2e6fe0554bc5a29716464e0ea3b75df99a685a1ec4e8a884906824437ea5a2ffb030d21ecfcc3fab28455e4b504ffea6901eb9a5234885a499c3854255394a5de1e3eff2ef48c5c15aeeb369be3aa4d47c8cd56a4f90e7837b5ba4ac41fd941516cb940b9f4553a1bd9ffba00aacc53859bde3e056fc6405bcfb088facf6473c31d9f6b2dd698815cc9f39165fb5b4d41689adb9ce641b84ac33ade0672a7f67ff966e5836f09ac84fff4a218792dad7a8eb4ea1d31c0bb1b4ba9da769dcb81b70a728cf1fd68eef7b9f40df18491bea099fe8c52cee05e06ba157b1d69a7cd240a41daee3dfbe50546eeb188327f6bfc4ff06afb6ced5e044a9332126c9e87fe1e967362b6c22c9b050321fc599dd7689983e6b406772a910d0ae3cd735ca7e37052b7dee14e18ac2cd90cd4a087b612e133b947ac29bd51afe370c1a36d80d7269956a4f8cbfc65064e2ba9c2c0ced2a3011609f0c2627f33c491388c8e8b041da845e435918a4fc67bbb70f143b8ceaf5d4e7f0940f95347732a182ae8d8d0ad8a01c244b723f41eaf7e674cdb93c517bba957fead354b88f14a26605e60014cca06c02a16a59721d30a0bad718f19911c81378706ca331d44c3a1e6fb817d7796b25d0673ddb957185f632dda1649ee5ca784330f9a3f0b622ef188f0d3c7cc2ddd1826837844e9591dfb263660adb77d18e2a300822eaad0b1d5337c77883de4f84b3632eec0c5203ae4285828940d0d55567039857d8da360ec637eac5cf07aeab45c3f46d82e5686873712ba5dcd86d4036b155762785634de89fbae00f47ab4956ff3720d77f621c4087648f11555f63903324003d8c622bf6d42c9b888cca16ba583722838e5835eec40e96be465fd78ad19250e72c1bfe57234981be86423cb4c04332f155b9a9019e99f9e98e27691adb3cb761ed0cafa55a5d7825da8929e968b3e322df2803030b7d32e22c58d5793ed72182e6fd59bc5a7295f7af4dec091f64244013ddd56cf3ca4ac6b5e0b803f66625d2ea0cb0d8e992ab3185fff074d012f279e82dc25eb4b580e099145118ad01cad540b0a63edf96c068e538a45906d6857c9ca8e544cf90b42e9e4c45b6bda6b5775ea0ea0b63687e7237df787189a9b662936733b0e8b18bfb5eb746794f1356bbff609e9e56e61ad1632097525b038a6d2534305619697131c3a99e91e512a5df4826dbe7b77f9e7ca2a276a5204c2c5dc09afcecca2afa24902c070548992f7ea90e0b6a462f9d00ee0b6d808dd184824188ff28bef99877b02a0028ca95a4b8f489fd38f1bbf21779104a21340d6a652491d8c707ebec7c1076f83f9752c2b6038a495dda7a12354235ef6229e632109767c53b15378f4d0b47d046066dd2d9e0ad42b67a0445f0f7302d5cda8afa27aca6629a91030b6e870270bdbb7fa5d12ffa991d431d52874fb2dc7442efb69d02911fe20b3bc252bc6be49f8b4689aa3b416132326527f38dffacf06273bad3bd982402ba4a4778288e0e031335b69b098edfc760abce864861ba1243ca948ad028af2280e844386c185c56b74e815005b7f21e55a0b578636f8dcfd3b6f2b7506367052bdf1b8e74de39732ea540743b98fae503be6dfdce3cd988a911a21454197;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdddaddb7cd4200c951a92018a980fca3969d4825b8b01ca9e56ff2fbe886372f9afee6c427f5fe96b94d099fb6bb7b977afa7f28ef323b87000da060b362577d1e90eeff6f69a7cf2c809de2ce6791e3189c0df34218d5121e501bfd0a4db0111c8990df711c6146cd27d8fb09cb539785a0bbf6736e1817eb2ccdc6bd351146bc09558f56a09cd19c991788c60f62181f0c8f10832398d21f3f1a993097f8d67280fcfc19291e272550cbac34fcaf10bf06d8959b8518c19e327ecb68ed237fca9557e121c6080a0c0b10d3a059068fd53038a057f18bf8306d1647d7ef7c9e20e5c6a9ed83f582ae8166903e8137d71e71a6b6e31f736a09bff416ed89b5eec5d912d352dceef8c809445c55918711a1b107e7bfdaa3e9c24c1d3dce15cbf58c5d61ddcb30a59001e7473f26f9b59521f7b32633e6bd96c98bba3b7060534e2e07396100a38ea8cffcab86815a1874347fe0a7e0d9456d81c241f7a97ab788ecbaa7740a7044e0397bf74a9f7dcb10629d0b7e0b032e03de93f1586c354b65e23becfd61386d781bfe7e6cad04f703f6dd15a9cd2cc143a321fb8e70f5b7d9537b8bfe2f4cc204b1457c39ef310aabb791155ddd66371367d3337d0c37c60174d4542a35714d82534100b2a95cce3b79a9a3f480533fea2a21b4dac731f31764a669242d5e9d35c82fc68e71448357fdc311789c5ed4c4c05a2be1a719ee79b45fa65c8ce68cb3dbefe0fdca5af2064f139068de5ee1cf2862b9bd806fd88e96e63ce9af23b72eea699d56a53cf2e5d6126f0b21727e5cf7e342c894ffaf390b49983b3317d902e69fb0548cc01ed2eabd4bfbe7c2a4b5c06f390cf478231a9bd19ddfb28acda3deaeb2f934b5825f85989f254cad3f378e067d50fe50d0bea056fd5c3904d0cd2bfcd39e496b8f7e83a892ac29bebf131ac0c9413cf7de5312a2a0468373e2c3435de96c8c9dcdc6464f6c7b22e31e54ab49b17cd085e26d0f0e15bf0d9af8045f27a924cf54947128917678e72e77b8a2b0b093810b460556353f817058567e570b7a4e83343bc4a1a6de2891956bb939596ab24bafe29314888aef219ffcdaf930696759f5e86414a95734440ede33519968f180f43bf2bfb67834475a8f79e055e8436ffadea4c4a629cfd67dfb127ad6ec2f42855c6da425a5a6c776e93ae6e969e2045ab7e987a768085dd3ddae305d0170ed9e02dbee4105ecf55fef0227abf3df028e271017bdaa59e75a6090f8a1cd68e46b2b3cbeaf45c9ac1afd27a7399ebb3171b3a8e6938fc3c1b45dcd254f4ee2dfbeadf01168ead311e76d5b8d0d22b4684d119db3e9047c0140c15eb17b313976970681fd20d4a32c9dc165112a4cd73f6fbbcc3954d27647db6a6d981b4c778e1977807cc3bfcdea4257df43cba25e1bfda072e8a87ae514f49b03d4ac00d430cc5818e79bf774fc6e1dd4c17be9774bea8e6912b0c8c8325bd67bcd4c020a5565ebbd0946bad8c7b0537f3e39ba14187ced53ff261d1f633be843a6095690a2e0b9c1357f4a3534134b520361fa10dd350c3d55798af3f152bc821d636a099b960e89acd756451af991d909caf9a3b35ba96adb8dc95e6730c63dde265d97730e1d0ecf1eb372ab61eff7701074960a64594e4a4490d3d612994c93e3d97a7f1c0c12fe630d4aa10128cad7c6561db85d06684db0e0fc1f98b0b4308edbcc3f51d77a991939451e760ece16d099fac9c55107f9608638bdcb4f661c166cb107d7d96cef81767e198c155c7d6063f2ab754fcafd830c7c7cc914d327fdd486ab63900921c8a1dee531e37e2cc5b69a3a52151ef8471477b8a685cd4629c11655fe91b0d14935d2550f3b0762505369590df8f089fd93e29754f3129c3ef34c84f2e0c3b211b562b4f5bccf29c18122d646cfc416f5757f9fdae07ceb802a215fdd632d5dfeb48ab1fe39ce8a1021efc2c32d9f421fcb07d2f5a1ad9e17e1a7b6018d6af2c6f6bbb97da7101d0f4d0976ba581c5396f901979138f8802a7281d1b1a0aa38cd4a78e209bbcdeb38255f92c8a4c882f411fdb49ad0962fd0aebbb441f0d2da69af6728b93d374c6227c8763fb39c3bb4f4f212a60083eb7e423d43e187e5106014eaaa29bd619b5535d59626a290bcf7b4fbbdfc73340a48e884e75539adffaa84722239b4cc63915ca0f50b934a511da3b39ee628be64f8928642c11489744eb74562aed798a25ce995bdc4732a09cd1ad5fe8f916b238ba8b6b47fad3c48f19089f550eef45d1de8f186588fa3c9b7f6b69d948de1c20a2bc6a358515f779aecc5b0f75f3fcc668de23ef0242941b0d78e1e99c1acf05cdcde7ea835093d390a96752aaf5a856457e750b4da016fcc9c7b0b81d85df1cee07c29bbe8b687387610e350f95e5e075d26af787ccd256bb3501599cebbb28192818b6cf960f5b5c9943305bdb25f2659d9e45b9ae08b525a06a0e8dc0b794254d95315e4886f801da75c494d899f809b7f53bd30044210dc7955640fde2df26db42fa4490a56583c9b56d6f309f11bb357a416816010e69cd4deba74f536be757c3b7d0a73ba9a8cf02002f0e02b1b974eca5037ac4c4f22ab5da3cfc21b8c4e5e34ed646124f3c17f6f24cef33ddceae829f40c0e1aa7642e5f6627550fb9e31bf6e5069fb167a9031e87a20a6991d84039f193e9c8e46e701d1284da28c5f8e6322352888f3d676d974c22636b8c73ccaf842627e2ff68871c27ad05a18999a1fb2cb9e6ebb2b66bbeacecfb43799fbb3345e91c43289196848c3ed9c795a42ba539c99f62e2a1e4c394ed5c84b7403157e171e281432ea051e4997400e2f8e95428fc3eb5f6ba4d9a2bd6fa321414e2c6c5cb055a855e031b022077b1e1ef86398b2814;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4d2e7549fd5773c6df538b52f1b4f4d9af9ade8d66feb65615238f722ec8b838b1def2442f035dcac88414a07b6268f0597851324beeb03e9abe62568d8781d5f7bc01b3a44f512c70a57f56428dea9353205f0fff5b5dc5e86dfa7075e779f7b37f483e211a9a835818188b2e21b4c5eebd2aa8b793e2e926242878ad3798013bc12648d0ec15feebac4e74dfecadaae3df4563c32c5c3c4e8c2bd7ebb98053de4c6869251d696d5af956f3b26f9f188bf7c8fcb9fabd78f5f170faa7751cb36fe35aa41c4067d3f9e9aaf26392773488e70dd0fe6fb87e726223304692906122ba1b6ea15dbdfcf25f7be3278c5777b9674ab9fc02f4210c552ebad0bff2883b784c9591d587a8c1008463fb51f87a31a39c3e47ef850ea5ed7da12c19b471b12161944d2ba73e5bb37c8c1aa11cff767394ca1ea149c32f22ff436646e30efeac2c4577ecf3710563cb6a9125676efb13e08ed1f74b44ff04d28e7de0f0112ea261e31752d7243baa00041730e4530d24c735ac750f870c4744641fef8f12e2e5ac5eb0c450409ba964bc67385181878e06b3b43c5905623e8f76f0b028763935b3daf852984bb07c1dd0ec1f2c5e0365dc7bb1f963d289728f2fa4e6f9792e7f6265b73dc1813645517edf273a7648b32f59cc8ff4406e29bf114929a91be9180f4a04803152d19c563aa96b0132012ce3ea55adae6c86a93378dbfbec93a7c5a1c97f3fc1fca5ee168efa5cec36dc876d7c446c44ac0397fb45e424383b5de6b57bf827f5c188e4fe92d0955fc66d1494958d3485994a6b6156d50bc5fdd678602217693bdfb0c8054ea1871080cfdf2559bfc4144d94b99c057fae6aceb9db5bf138adb057b430578f032ef49f40d77d7a93f716e6ad7de297cb0fea75e3aa137771ab0e5e223eeed360275fb3a5370a38d6a9191bcc3a682c56258a0a536fe708465dd692fb301c6b28f17d81976e5236c8cc15f04d1a1e46e210dc6dd3394846927cf8e98fecc5f06328af7d540911e15a793d7ff60768d8998aaa271bf7129c1adcd84ab9a8bfa30a506831bc1d8ae1001f3290cfbf8560311e9195161cf37edcefcbd058b97f157ad2f33be3be9c0fa8407c6e1c04f8ee9a4d94813783bd4a50fe368d96d502443027d193d42342999c5609a964a1c9b7e4faa61a3f628b36c6fc30564c306474417eb7e9f6eea28d82d966de5c58839f8c2a20e9ecf99bfff727ff292bc9e04d5dc980a032b1af8334d60989d6efd73af92ff1021a44ad9473d9a40a3027eb0c7265ef9f4bfdfdeaf8e916ba3461504360e5aaaac8fe23a913a8359f3a899a1e1b37c61ec7cf92545ac1fc3e88b2d2fcf0fe8051012fac8dbcd5fcc8caeb686ebe7e43f8549ec3072be709aa97bb3dd2c1b144618efa05e586e29c4c6eebd5517158bd6c7bb275232fe55ddc606b50a47c98acc78647ebc93541d56f09815f65afaef0cbc870d75a2402a8abe9be1b1d10c134d4dea1e8670cc7d6ef1d7c5749343366f40a2a6ca255fc352e6f156dcf0d44ff79f559e020724f3ef472b36f851ac9a98f0d125c92876aafb63c132e92c9a4dc392d790b2937d77afeb6e0abc352cc3ccb2948fb871240fd5ae5d0a32f219fdc9ac4c9c06a264f3781c87746ccb2101fd1e3a661128e0a819ff4f10beab124af60cf5c9df01f2d2d76814884dca60e058025f8eaa087350ae26e9f3cc4775d4247b8210da796c64f1345ab391bf629a516028f0a15cbb33b31097fb666cc5c7b418ab45391220d4943d3ce254bf3863868b843a0c78cc552737656ba9d0ee4ef2788e3e5c636ef7f3de7c2571fc742f8fa1cadec3c24675191d8500be8c5717f69c943d5acf1c88272fa082e7ca3dfbf5af322eb495153a7a5d91dfd74c9173ebd0f5213617cf308147a90b3c72017c85f2956b3c1c75715c2611d83e1458d5fa509b7b2bde306abe0c7d9d47736940278aca07395073a14974b4ac5abbcc711ab786794102ab178f4c0b51e0eba34848f1a68c97247bbd6670cfff1762e3aa594442ebb7761c07048bd37d772c26d1be16f7a7b954d9fd7bb7be8e73787605e5eb4548c8ef54e7f38c8168025c8432093cd470f8146cbfb0763cef5fcf7577ae65dff664af84d2d43b810af17ad613233b88383677f113943ea8afb7fde0831c978fa0883fb8c068977033c7035670884dbe71031aac6e291e4f3c82d8c12185c60aa206a8085fd952051e27cc4cfd541768202dacbc5f2ee9bfce33160154640f6f4b5a0775c77000009021add6aae14155288843fe6a4e891f9189e676f0df123345b07b0dafd872219e2a753534bbd1a7f84c8826d1cbbf53722646157f54531f1425d3ffc71f158b684d6e08afcec6d9bf713f16fba21f1a874c532b5f7ea93604bd47196a7ba72a2cef95527fd39068bcb1c077ae560262365048c66971462a1e15f33ed00eab7bc6f7bfb25fd9296cbed730e589c719e0fb4e509ce0b50079dff8332b81494a6e206a93677b55be98e7e6d215d02284f5ad76f7ba6c5782c912148c68b9be497434573b7240964f2e26c325074466b434357af20737620e9fa8fdde87befa4dcc886e4671e10716e2aa41289646f16dcf3643e93002b5bb5ecf5ebcd374e5d5637f222d9d47122ca12dcc5f67202cda72425803b54b81908c99a719cf330f290e14ef20b170d1b4ef480e3bcc5733f91b2e078c39fc5e90772de0d2886df764b5bb3ef20d6e10a6ebc88b84cbadf95ea71cb39aefde09197e3779aad0b52ffdf520da5076b0faddc024c105f3073235a6fee564e1f616642ccc267e1222768646f2e9fbd0a82bf677e72cd33f04619f42889dfa4cbc5c60dda8f579f1775e04c9b4e7c8784dd0303a3d9bf9820e0d89175077c61891cff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb1d3a5462b98310d575210e81f11363a54a26a029219af41db729134b031802d4fdaec913c725017e2303b39e3386da260148022061dfdf5e019a3e57f68b17ea26ed845bf304d93a50646da1c42cecfc1a341c18a27fcc615a2b3e31058918bf43245a5d157295c6e4f1e2a334d8431752caf32ed2c0cd2c7179188bbf34bbcce1746ad0523c8e03c2f2cc8421a7d7c834708c6c01f0228a9627c3e5ac840513a1cd17a77bcb631ec3210eac3792c4bd4f060755f4d088fb1653b49c94b67a209ae9913c9e4895c28031e9ba33b20410034d0a7de74326d2c977dd996af19a7fa07923cbd756588033b61b7e2395a3ab921bf87fd3eb3795824f72044d1c630f6b7212622336d8e5d2027a1eb3f70e6f947df1f740c5ea096e69efc900b22f22098509795e6cbb262580aefb30f964a9aafd02031b7b4d4c95004d669af973e12e082ab78abb1957bee9be72fb842c0afc46b9d1b92c7b05bc89ae5aefcafc8d1c6d564d59394741503aee159c0cbce184562fa89c34be405c31fef3644eb60875ed7ae6b36f528c6b0b0c2bb7a08f95c7606b83175e278b75525551676b29a8bccfb6c5d74a56b4ae10a1547797f3c229dfd4d77ff8d4b4cfeed3078ed47f32e2eb9cdde99f23248a769718f470ce3e7880a3012e7f0f88e648890d014f6b4b11a6e1e07c509f5524dd62421a5c15d34751ef9f571419e4e990e1648701ec5d93714584bb3bb96bdf221831f626c937d5658a3e450bfaaf8ed2d1abfdd7a608eecc3e008e1e810ca931db9c1551c6e85729fe426586dfaeba673a7d3cf53431e8bee2fad517b77b26efec8e246bf4efa859c4757e68f159feb9c18195bbec7bbcb628642b6029b8286ac94754bba1b6b59b5d2ddba51e220970b07c60f6ed1726a41cc362016a7b5fe54e9caa256c500d79ec591a1351a3c045c00b1bb15e34f07297423053cb76f8f30a9276a220ec9ba23fcbb8783e2a6e85be8fbad8d4ca1f92699c3e9eb9a1a7e4292fa69ebbeeabca7fd906fe7e73573dbd91e1cd76f2c33421d7506707be42eaa1a7dad8811b152d4ebf8e5d2a1e204d3f75044c689d1425fb2e29cf38535da7afb7bb06c82ad1d381d9e79c0f8ae800ba5848b53d4e27efea9249615826411057c160a716c8cb5113b6ea503b70141259581b2b46fae70bfa2757d1a0ea9b8a5aa3ab60ee430e81911468b4af06ad070c9644ecbe84902f3c2f6d21e1951871f5584632d52857bfd765090e7fe4bf423a415f0bb5a5c1a514c3930d3efd51fa73f7a0b68804ccc85b1c9142a4d29630948d6fbfd2376fa882f1cbc433d5109f65b6182318a3bd8f815fbbd66dce734681862485192e22a094ccd979116f9cd2c9481d1b80ae6f15adc67cabe75b33326ca73f32fef9a864cb72266267cfd8418aedd7bda278601709023cb8983a2d435b3a40cfdef598319814b8b814750e3c25b5e83aa6e667325aba2364c906e221d792d2c6ae2fae15deec87cc6ae9482d6541a326d24c9751f18b6b12800609f13c57f0da2420d67732fce5236aad86cde26da85ec7468a460d71fee96a79f6bab4f4196a6e1701c03e3a506660e584a654f915738b01ab21631e3cf21ea263ee9f9ded8beea28eca5da9fb5713b3d484e3e49279d0b54231a3e389ea08a2a7e330db4d99fbdb9d57bcd648a38d61c15cc451980557456988c0fb63b8d872376c06abf7bc1f16fac9f4058985e9e324d1d4d6df647e91efa926834fcef1f1615aa1ef9dea6465a28e0d9411823684f1674444000026bbd4e8683a985a45cba4bcef58c9c5d3df016dfdc476ef0cc4b471b37745b06e0aae0c3cf96d0df2d8ab38976c97a4447be17fffbfccd35a8a095f15f9e7f614de389d3e5840a2cc6c9f550a62d2e063ef34f130ec040a301e6334f1ae45eaf189da47519c721ab1b082b190fbcad5b72ba33b787bd22c3c21dc5a4c9b9f36300c46431dd51cfbb8ff2fb453946bb305db736a5a63a285e60c7c43ca6e77d82ebe02fd6c66fbef2f345821bdc3d130591053b5d4ac512417595f28582bb299ac6c9af964c1c320ffc5b2ccc432ed54ab8db079bf98813da244534f4afc6ce84a8a11d79d4bef30cc38016b34c894e4f7788144830213545c5f4929da02cd00b798eef90fffd1ad81d8fe51bdf5c2d40cd2705a6b10387e99ebded54415fb8f13db9b04357e225f2246254d40bfa91a4c9986558fcd7623cb2eead5c1095643fee2b7e88c8a36ebe6ad649c503cfbe5d8005efa444fec6b500fa58541d71f8be3d1fb32bb2e1b905867380524d21acee5817ed7fa4d1c947836e336a63123ee375b13bbde9a16c10d0978bffcfbea7a4d12530d31501b5ef747c8531eebd427a8a518bc1c192ab8b30d0ae8edd0856b937f37232f43d388790e5624f49be751ff78aef0fb71b5e6f3152bb65e9c1e666b387c63bebd2afc3c51a1fafec976c772857d79422540404babc20b78255f22ee003d877b198e1dc0e5b489d24f98a69576bf26642c4a3b4e221a55b235b9d2a79d969925fd0f52ee42542e78706f2ceaf040566deea84788acb6d520456fead4c47e3fd5dabc0c563aa8555f7b0271dcb3011def57ed1c48ccf2eeeb898b3b706a547f68589c487f370defe926e233db22095c4d2eed3195e019d35350cf9df8f48253546789ade9df7b6ad7a5859b564070aa9e366aba312a185fd048775a112f1bb742296a1384bb4d1fbff546c375c49cf0adc9a1a31a1acec8f00cbd85fd1ba60164df6a8447a95debcc45e7ab6c6121b3f6e93f80250e3875ba8499ece2226cc2d239d258bc8dce4183b95bf60b75099f7b49b2b1da0da963d8cd506662e556786e27628327b164fdf07eac9b99ebd16fcef5702bff4f31aa3f908a8ff83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h921d23c77ec56dbc542ea7b873f086fac7fd5d8fe7b4a9dd9111f780bd05c49edca2698f5bfc708215c3ccfc53fe5060032fb97da630cdf2047e648f2bf7449e848f9d468aeeca8d1e4d2dc5c345187963b64ab22668b4dec41aa610ce9b6203b9143860c27796d4472e90cd97e7d2ff548dbb18ffb3d35483000076b8604e329f6a8ea0a7604725b3ba1c11533b03ee9899c40427a2b200fe4e89b8219ddc85ca2abb35c8c4c98ee8ac658968de051f2c063e1f2e3e5b05d94fdd53ad7d1ed07811221b31647cb2daf6d189fd313997e1031fe9db23fcdc8d82c3407d3c3f1ac76147b2aec0aff82bb4a3d5e6c24424b1b62d5e834a51305052424b0416df81f717250327f8b8bb2526a0327659af676750e507561108c5025ed12000c065bdbce0f28670b85996894f149f6afb327e34aa0947008fc787cd67eb9a1355812bba895d41a3f4a8a5134502aeef6490cc58daee58fe714c3426b9f43937c7f1cdb5517d64f85f45ab5c6b3e7afee98dcd97570b49124caa79f142572e5f6e2a105cdefd964421c3d8ba208a85ac7796d04bc45d3c532f4f0099138fcd682e5c0bd3ca08b27eeae39124564fdcf6dc9dddab392b5894b2bf727b2c661aefa838a1d3a4b5b63f9ce5858b243ae3b32eabf13508d05a863692be1d6cb8a632a8a72b5538a4d8e9def783a31301c42ab871c5c7b1d3c412e4522b4906885d27d1d4512791e84d42d7b6a76c926ffc9d94f0933d4526a0441f3a8b6a1f5f0e2a1712b7df8e6276db5ecc741d4fed6123d8ccf6c86d7263869c1f1fbfe6a270f1381e71c6cb52e93f943190b9e96e96a4d5c396cad679eac9f1469f12f984294df8cce4448dd8323fabd165eac7d558976bd33711b912df8ae8b6ccfb7bf5fb196d4415a407f7ab22ad5531d1c35ef4ba342c10b992eff20b24589edc3ebb6791210c717ab49703013c399500bce231de7643893c29d8e06d892ad5a3f2336e03f9760abfd257dfe46f466925a85ec8c8bd31c4224e9da90846da07d4b8cd9fbcf9ac187ec37cf75cb58d9d318063dca4a2ab06694c92d17a85c307677ab9c216f0f5c0fe5feae329296abeef1c261c22e17aae37ed76fcb5100fa2051a0fd9de3f16090b86a1a73b1c1ee7e6aa0c0d03a5734a205e80084febea15b34a4d17429a592ab7dacf5d9b82aad870358f9cae133bebe03fa9e3a14b9ada2de0be73a4b8e1e54ddcd7071a92986f49ea6df88fb26fd95cbecb07951781d33cf0f9479d9785e6f999b66bc11455b719631b2ce92ec6dc387b6dcf3121c58c3ff2cd43fde9d4d664336a8080979d9196313043b9ec47987c9d3c8b70e717514b6ec6f588243c099d5a6d83c3408a9c733bf1f8e83a3ff0ff99ec61eb663d3df96a893aa48b426163b9b3ed1e97d266ac6332736c2e24411067646f07a37838cb10eff53ff872132a5ad0838b8654b9a9ec808bdc690a75fdbf6aedcca79166f361d6cc7ad5abc18d66466e820c8f3a8aed0220e073cf6869c5f9bfcfd2ea14b29146c07cdcd548a218f3a6d9dc99a85efa98189cc1b974113f02df516d315c3de8bef391a8c101c040d0c86230be476616da291ea3d2d437da300dd8852aaa8bdbdbc33cf3865a9f4ceb7c71cdf54592ca3078bcc62bba22bda056e1aa9603cd7e65e2fe9483980533ddbbacdfddfe69a1ce391377ed5d43dd524bd466ba0d28f2f752bf96361badb3ef8277183b9b77ce0a4aad204b88bb6e6d6041856e2f8d83e6c59a6472b5e35d047ca9e07d7b17e5c0f798f27eb2a5059f2b687fd710399ff1f273f1fc25a595ecc0727bc079cd645fa326a992891f4e8be95c8c68e6dd5c5dd3de848b4e5b1172e856a5d13ac82b4e05e5e8c71420e3a703a808f6e0ac7d0b34f8025c9a96b4cfa1e4309ce04d735af507dc44a4dccd71781addb4f81a0d3649a4f470055496b665d5dd408c31d5f7f08addeed8de8f6c0486943da3dcab9c3c101e4b9392c398fcbfc390dc54b7447b4ed2a226dac7aa839d93780087d7e62e7a5cc6db5f9b361c763084f8b13d80226fb9375a7f3f27460bb3e14dde672998c6e936b8922a2b873df5fd9fbf22740ccafa133afe06198c76ac03112b5256ca3547d742b34f80930da32d43feac83327b8b46ea23226374494e6f9fa0564f893347583cb4245f8a6f9f1d3ec48116b9b5523349cf472c158efb8719f312ecb9a920842b39453d57a797c09ef077e5f1038db4d58c317b1b14c576373c004f4464c42de411b271fc35dccbcf25ddbd0383b3ec012eb42144b590c19f2349680951d239c1bbc70e1e029ecb09e208726703f12b1ee9d173af23405786b05bd8c3b80b1e1e11a51009a8291a918afccfcc53767c8bea7bc25cd00a3646c6b2522592bacbedba56e773bbdc11e2a62d7508e8a5c4457280fac7d723c1fd5bd6207ef320704dbc6cafc35f10061c099ebe48dded5a24f8855a6df16fdd7187f3995f353e9f2881d3426bb7e3d40c1eaac8dc7f739e7e5cdfc4d578028b97e8e049e0fc6dc3c359005f0b76150a51b293777af85852ff9a118d2c0af4b5b5ccca40752b752f23a0b8d94477dc03b2424162abcb84849cca157e43f4aa2694d116c6e2ffb95c8b4c486d86ea69f1a6e4f7df5730403101c87f5abd2170dd624d96284481cccfcd8271683598a990bf7a92a0a6a5293235cf44bb030f7618c5b49241ed061eef85c37a6aebc57472cecfb6ff867c15c68b0fe161618375a49620fc4f5c76873384d85500c8f9232560fe08994d83f76d21b0e05c0b676481db3a5382e48eefbe38e34092d4aee2a989cf2d6b1dea9138a354b1e836b948306eb47ea504b96f0573e75e698cbf6ba4c37af2fa44330834c14f51e7fdf965895188df0755e328a1af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd9b1ae39244b8ad64c54230e0c10c33acf89cc9b22194f0e0395a769dff5199de656772d12dc64dab39b33259a45fc9ec3c41ae8f1ba52cc3bf2ab5a844e82a0237a41cd6c9d5b5b22f1fdfc5fa643c1af99c4ba0e3bae0f8b50ca1191475a8889579bd5a7fef0f95a5a95865add42bd7ebaf2a2194728ddc7bc4b1ceefc799f38867acffc1f3be7e618465551b7684f843f26a8e369f056d4980fd56ff2a5d1da4974e692806b4a963a94d65cd5e1426b4aef00d527e2847d4d3bc4236c6b79040cb1242cbd649fc5e0c6949b3ac7527ab2712a1dc4d855ff27b5a3ef09b1b3eee5ca9e66e936fd43891166b3d879e3e6e032fc3101316fe88ba0347371f10cbfbce0bdd42e8ad6986f8006c1047658c7b2bf8b2cbd1771f2cc968dfb50e88ec2c48b52294c19b83c0453b1f80451a2a8e6553770867772b2a271beac70edc6de68435f04135aa738a70b60b4d569c41b8fc5d5127923fd8c2536c1850d4699bee3b8732f88140ac6f403846ccef71f048d2efda5534b7f6d8148b685e4cdf9e303caa6fe6a0bbdb2c5fe0a92bcaae8d5a8c7db333a740cd4c060b8800c5fd79423e4d3a77c7f75dd15895a4bd3945414584f362b5557f6c9e1ef5fa75080121815944bd08da9ed72c007ccbb5493561077eeec3567df68f3200964a900c7b56194610503243e6ae2fe08ca63516ef6fed190a95667d11f101d4a6cd86c51554de3be089fedb64fe5a0478a7ec696659a42d932bf3ef73c0078bb5b62367e2ac0088daca6bf35f508a86d24c755b2018c0c5f81f2f650f98b640a15b21b9ca49ea3eb0e865bb57a0589879d12750b44ce3b9b50eef1547267a939cbd1f143e0c6f87992ae7d3edc7acd79cdb14671fe822a4fa0250038bb18c2d0577a729d58f3a4ca8b6ea3d45b1f2a90f1a24f4d5950fced2179d67f05f81d1343591b7ded5142bd8e2d8b122c6a33735084d8ecc45cd3a8df51f80627f06cc10afdba095c49a2c9d4f3100da2a8414ee57d86bcc68ca5acb470bf0ebdc75438d3c805458a62b7a943bcec0f14efbf1479f511a241cf649524766ad457781fce7a988cbaca55187873df723895276b7ea0d76c20c22e060cbaf483b2e68f9b3955a0f84d8a09fadc9d8b7153627b5922812bd2e57dde0a1bcb86eadac35c9910d2b6c87ca53aa06ddab5074eecdc3b213d69a2c8f9535f4ccba3da041a2a9654232d26d64fe2e378247e12cf8164362d73ba8edf1660a3fe5b3c96bfa63b212193256539577bb35232fdf2828f44af75acc30df5077612e767f1f3cfc2de4072c92e97bdc65ce68c3f6b7f1c0c9aa0eb44693f85726bd64ca395941ba0b24243982d6649178d9f9b3373f41105cdad4b3d0a914ad457af6eecfe042b01401b4b66a253335ba106bc89a854430e2409cbceae44e0bb5cf3a7bf5d8453536844886717bd6dca9cada7168660971fa71281db8ffc8646c00a0368f26f6fd07599b62e8b571a0765c6ff587f7ab2d0a6f2cb0f728f6b4894fc7fbf2e0de5cce3e83b98fdea557300a793bb84642f04944931d33267f8e26a0c50c198518e0cde0428be41c13fd6236997ab0d42e26dc36c809499a80d72679e18f54271105a4433749169b580139dc23b88584829d5e81cb6a13260a6f08944450b87c212615acbeb809a9912a47c14dd255907f77c6097b86970c61cfd262ab72a2769bc55b74d389a6da6670038d1c92148e9f766ec7f596a7cbb9fd7f7073c39e0e36e0cf54a52c38b21f9e53a3acbada8e59d9c1275b23845cb4f59bd9129f14d9e033903dc9527216d0814982d8efdc32af2602b11a521e5d47a694ce58e7b05928837bb2b3b3475b9ee2f640c729dbac36058af95ff6ede61c70d9acb101ba29ba6ad8bcd44f22a23c8f2147b8871388f2bd1a65e729ce096f4328b25bb816f9b313a97b5da7c570193d31912f3646160a712ec24875cc0569a68c2f4bff787fe092636aa5d3e0a37e636a7d636c5fca526502713398b5cf85d355640853a0b51b96448c87fcd934dea9ca3c8a009e52c95b518fb4ce544173b855e541cfb40928c4f27b9fc312520888d24609bf46797563c5166be42035c2125bf357f07d286bbc38b238ce4f6a21e8444e587f041fefe1b95f7d77b337d89b63164bc0bde43f7b5c1d7cf34b54e2e817b1a6d46db749ce9aa01b0e97bf1a134e1fae364d712f4633007824828985f88e1c8e70418e7ee72bed4cc67c27db8ecdbc7911445b3f5b8dc853504b42defb79670611be9bb0e1a9ffb44dd4fc98fcb74702750d0dad54b80004f9ce7b619c84aa7368df8b44f799e6158c33dcd4970140889a9e3c0861b1f5ef610498d963aca1ea71eb2baa26624b99a2ab29d22ff7fd029bae2c36a90b65b8bdc775d431b9127eb2b8d99410f4041196abd6fb73e8afcb0f4a07ecc89dd1b993c927f1b9675cc2b57a537de86e015e0b17afe56ade91e035415c2409a895aaffb39eb8cc1579054276faa5892f36de4f63ff9de6e505c97a355878846e7cb318e41baf2b556690b4570cff89806380aef701c8aa74200ea833fec0a1029b1bed7dfdb05f34ceb5d9f450579ff29908377ec8ffd33a6555e0d23d3143cdefd7937ec5e3c429a1d902f7402a6005b2b2e9d4e88506d1a3ef2336a0aa369336d16c722fd1e500d4018ff9c4bae5eabd8d53ff8b2e97735704630d11f92054ce35e79e91de2b86983ee4cc92929f90ec2111580bcfbf3cf18c1e2a4fe3f292ecb2aec6e311651096c9daddcb59554544fbcf570410a0a208e15c1df50482ff40ce5ba3a78676ab389653fa2563e126fac601d8368d07491390472d595b3fef033a0919644b3f4445b73ceca22f84f11f287d646deb30d45def759c4525cf4bea812844afeb499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8d6296671a7b09182026f4360d0e1f6d57b4b33418ed0a825d0264ebf28e4b231645e82d6eb10ffed8e01e6ae398f9d0e9a6641e7e560e2323acea512bb2256b7d9dabb10e868bc61e86e2a425c9d459f102af7c28bcb6c24e90f3be5be6f5081e456a786eb2eb7a551931b30b990fbbc319d9919034d40006f4094c97fed668a74667a7f15344b87e0d1cdee00ab9ee8aaace70ad425fe470c2154e872219a7b72a62fbe85b6801254912db220b1d6d8832b8817f13a10ce5b7f643b7f15e0bf2b008764fd37312109a1fc262ade8359e2e66bc17c0024ce6b60ea85b48eac82e11e215ddb370179a37abdda9d5e5b5ad3e7b46582d943b603f461399bf12b0face318056b97cea14ee1c9057ac1646e79e2e079cb6723353527507f82af7816b1c5ccc6461599f62fd4cf3858cca7b121ff1053baba90210ebe840b9b4fa1b13c9de2050f6f7076a1b79e0b6d5e9762466963275aae65a0b87a7d071d62d6258a8304bb183d1744b40077adf5def83658934ebdd9f61c4f21a4c4d860b35cb79cc56691fbcb10dbf5fdc4a342acfa177d77afa8659f250d743727d073b7e028ec68703a3b0e62e2c406134d80836f4565bdaca98587d5ea011b6855a6abb32fc2a2c9f234db387cdb69cea4db8bdb142460329bc0dbeb184e87c955212258ddac8c4aeb719a121481214df967677e356b9dea8cb8c642dc81fe916cc454000f6329e9fb87bc8250d92b97a979ab3a79e0a99f75474acd20a90f6ba9c88e3322100d64c6c9eb5b2a3de8b24ab30a7bb48e68f1439932591edb556a24d690de3e8cc88f2a6a774685ca85009f4b0553f8ddb969349aefbe198ab8dd487043048d3db3e0526285fc6aa54c785c8e0a128168efa69e8f5bee6e2f3f241dea12719ec4410618999f798d5e96379b80885c06361c69614c36395c80b2638f1df2337b155b2c397c4fa9958f6a497239828a84a567d05a70534262f5e7d8759039ec3e28bbcfc3ee26e12f6091f7161161c67650f6434bf517dbe3d55964ea676e4a6bf7bfb61364eab0675f030a29ae0cfbdbdcc2e5be91e3a2237042ee4581514e9a650e4e859d80bb54f5273c63f6eb395946773963cbb626060518c22f85f522b39baea017e258a6ec240c79f5ea95a42bfa7c0f40b2774d37d93feb87a0eb9e7b51a27252fe29079495047164f8a52e3d3f94e6cc1beae4ca537c33e074d20dd195dba4954a1d8fef5408712e4122096809c7e2bf4bbe7fc299e10b66ba70032a48b58503f5b5157bde3c577766efabe961fda2ba64d0d0b5813b54d50d3e2536b05087985afbbf86b91a83c2c7b403de1b9d2cf26af900044ff12d10d44785cf93949205c6492245548f916ecd91015be7e109649d17dc90b227a3942b0846107d759bb40ec3239b2306a8d15dd91355458df530f4e1071299f48de47895bfb988b62c5c8982416ee1eef321d58b90fa2be80d2369fc129acb659b7d72b07afcf5e94cf8700c951bea604e8f2791eb6bd86a3b802263616086ded95a9968b9e964bfc4de6ef5cc9d21d034d32306aa59a7b769a7c30675906bd9f418ad89195b40fe8da61bf166578a05bc38a8bd9d8a75b46f16ad663c36d4cdcfd3a889f455b905be42e94d28cee5f32249249e42064a867f752b00dd90a6d40055d1c7ad49dbc6a629c981132ad169a4e38f50d35ea1b81045de0370a07a3d32719370184661810ac4dc3647d7c1afed6cdf4e998392d6e0c7f98275adf6951b42c98a6796c088efe02cf1f96f244bbe5f01c4eb6dbda943854677702e180356b35ed5e5074e47c1e1b8d504c1f47c72dd32a57636295e30c125b9a3240102a39a7813c7f3614b34b3d7be1fda8f2afcfd96e9c2afd4f0bdbce94dccf8b37be30a685e142688274f27a3b9abf9fe9d2d3c3e4c0011129f3d0fe8003c8148fa9c5afe08bc3881df51e44acfc7c512eb11d9eec834bdb3d8c90508a1efa94ba35b0b1e2f8881eacf3bb0ab6325e6e3bb3f44381c4771c8604f4f7659ba479c92786d01cf69032bdd811998c0e3e0e2d38924008eef7d7544767175a09282ac302c36b7c82dd89c32490b39b4ce1f2f70c9df9140d76b172eccf2a5c75a38756c60c14adc101dac314ef1b6eec1092fbec5271a24676d9e21d94d61f83c38db6a77aa7bc7ef533426b3e423002785accc0e59b6f81d38779342d9af908bd53b248295ff286db8f14839d9dc0d3a2e3d1f7b83d08f38b62c0ecc28ae3f6a348942fb53b990891794087723d553d0c744224702f2778197fc07bac0cc1c6f66c595117015a12f2704b034c6134333273ac59117fe0795e374231c458c252fe7051bd86c926f247d9cc0770ff836b951c7f4bbdc1ee07e33e8914153517eb9dc0b8fe87e1dde282dd62862a9df99afdf42422667ea9884d4f9602d491220c5f9d4d2d60810bc804d59f11e1717e7b891604bf4adfe00373a50503279711997d9548f8cfcfed1292ebde15137d2f6b19ea7a2bf9c7aaafc2e4caa84d6e29f1879d4e74fc950691c87909ecd315c459fdb818d318ae6dc9a937beaed3b1b2ac5da74af5c71a65613944e1766b0834e8a9b3a97ae3b25e50ee16c4ada25ba096a0aea16faed794b42eedac1ff718ef12f00b1d79e69e5e88fa95a35ec8f02593d5bd9df4b8d4b1768b9f7098ede15a20721691f5f855cc260278b63f81699a04da7014e3b8c0d34bdcf1f79a9f7dfe01f12b3236206c02f0c862091f10713fb88c7fba8752af642720d04d94e4c7db0ec0aa15d2987af3b2fb13d8b4f1a8430f3c563d59950213a19723a08483fb2c48a5041e69ae2e9588d311b414763da7b42a47ad2fd80349a5a2d94d34ab94b692ce43888ad2a5be1bd2a80db21765336e9cb985c4b70b7d6891;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd7d74ad30bf1c0924210fa79ddbdda8cadee8123ada417791e8238f8be1b6da798f6adb9abf141a9b43d6d0cacd2b29d670a196c87167d3ab733b7aa942d5cdeb01b1da13b63a0e8c60a21c9e3acfd52962be72f49e19799fda8a0e2c0ecb4c459fea79d0393d8ee7eb7900423db2086d78f88d1644d86b6e52373ee196216c091c5c307467744ca539b4f769a3d7767c6f3fc5a3f757215fccfdaf9f8387678d5b7fc092c533f6820fa1857e491d9298b217ce68946f1fec2476be45f0182a727d98767994aa015b89f71f0f133bad7317d3240f44d87aff02aaeb917c386cf621dba98f6b86066dae0b3f8f174fab502d9d7cb389a5fc7812fda0d813d81aaddb002c0f3f0e9936c2ae935571d8b3f2a58c9d5ef7b1e2f28cbe4c22f9e75dca1a65629e9549fe648599e2ba070f53e9fa1edd16cf3f80a129309cf177983c5b8daca51fb2f0f9b390cb19c795872083ecf6a1d871f852adc798718a7d17590fc2ef830c91930508fee59dfb289e866cbfbb1dcee5a13d5011d145b2d7944695bdce51ef6d5591cf492c89df540455c3347eded9eb55bcefd9b12aa4e15cb7ec8f55689c203a14ccbc3e716321d5930c0ca09b57fbe1db1d937c8acca49bd65a7e6916776fcee3881b880bf98ea9c908ea4e08a3cfa0b0e99466b40f5b4678482e303eaefd95e15bc8b71e0201dadd4cf8f6c7b7c558ba725db25addb5b1762053d9e32d4a703c99c7f1a78896544e1a460a086a727a057e090b2081e19486cbc25bc1b3f7d1158e760fd4ecca507a03a5621aae384831cdd781c228de9d279adcc71999c0faa38e1f868ef0f84593f50035020e0f690ab98e31c00ca4f60b245f598a486f44af15b89430dfcd8f80d85a4f1fe82e6c430547372c1df2a4283450125d124da00757acb74dd7e6790c70fd77454db76c5e8c2238f3720dbc3113818c0041a831378e8a64743d72b953838b2b09d47fbcb7097488d0ec1ff6b6d28fe730f2e89aa0bd59fcc667977edcb4881f68a78cf5733c421dc6a45ebc1667d53fd976a80454987abd85cea7adcb2c4e19d2a26d685009c4ac6c493ceed58461c98f9d732cc79bbd7ad1c786aeddb0a9654b7215789a574013300e81636c74d9ac6166ad7bafbdeda1f1a07d58d833c29edf0b680cda0aaeabf3871237477adf8286eccf105463dffb2c29211c84d59878c531ee7f86a1837b2aa17c24ecbd37579ed7b9019897121ef7a8d930d283f493c02d2c1b17cf25d1ea8ecb91acfc54d9485ad42f7bf974404fdfcc7e8f4f89dee6b6c5c8d8311133ffd710cb2a298cac3ac7bf4f21ee3b0eb04098e7904fdf00dbf28e8dbd74ce8d362091b16d70c0fb80553382a03f6c2997dd30acccd5e4c32773c076f48e8f0550a28b18048277d263507212c258692340b4de617d8bbe043748ad546199162bd91e9b57c426a4a5d3571ac7172a4140871b4dbc0e3c81e2d5577fbad76165eb53aaa2d70cdc8fd6f42fb17fe986f3e77d82fd787d3c32ed0e95cbc79119504869329112ff9e376853e66797945c0b09500a3f650c2d18999967ad8259eec1a28f25433e7364376dd8bb869d3aee1dc48b8d106d4f8da89064f104f22ddbeeeb4d32bc1cbc99f5cc972ad5199bb90239928112a69d7f2a2df9329d148cc9cce5a74817f1d5a7a7d564c44aadcdbf621ac34841dcac5f1fd2763f93c3178bba9f5d2e8cd37dc96e81107659f2f1560ae5378d7bc6d61bf8a9c184b7cdf34efa0eebd7d2562f543e4c7b29ee987156ae284c89f802364e3d799c5232c59e74e3cae5a0260041dbb9e5c6fde9cd1cc63729271df2dee69908647b9101c2146a035630134eebbdaffd89e025ae773a5ea6ef5ac0e36ccae71ce1e91e6b12a7837dc74c30882be5a98e429ea4d2c295053d21649d241a1e5d53280bab958fca323f71093ac3752c19e038479ceeffbdce1fa4efccc0d59c3307c8e76c310fb2cc64fc1531167fc8ec3275dc4a5f6b477ac18225cedb5bd577ba01c1c566f7af32c5c11a4553d1666e49d1178d2cb6d9ec626b4fa83160d4f0b8e8774beab7f4636f5f914a8c4849ff674608c08666461abffc5b1d931b20c257053c4b3f0532e97ab92834421e051f39241f1ee6db6b1521e8111dc8443336a4bfecf611c7968c34e44f642bc1bda8e90ae0c6f1610b080f1ecd454b6bc72756a4185d582bd86fb5db6d67821d876cef771a67bcbb49200712a8cdd4f58c2cfd0049ba0656770054b5d021aff335b891b5724cae1407670edfa949b7018022b1abb0ab9e45c8a9ec95fa3032a85042df8129d7cb2d84a827aaf529235c82a3c63aa60d6d691a72f81c47e11fc2b08eb3a8f96f76d094a905e22160f562845d827e27c48ac3d2dea2c3e1cabeb7416d3b4aabbd621f380a1fbc7e2d2905149ce12fe7347b38b5d0f995daaa984a8014b4d119c8c532855a2f399519d7bd73485b4da448175f3465496b5a6683f845cf98ecd1f5efeda18b608d5a88d30a090687ab21b0705cb30c29851eeaa63111a65fdacc3695c074f2f62672569f4f639932c8a74ac2024b0ba4288984735b25ec85e53d3ff43cd413f1dae8ada9e487e222e03dd8fa258204d72337ae3d91985a51b5a53f2cad8a22f00436d6ae77826f91ec43ac09b41ffdd3a73cc8bfff16111ae55dba36f3d2cdea429d737196a48f0b358b50ea5c21397f71550cca8e6a62e5c578f59a0da0b56436af8330a944ab0d3789fb3dcc39bc1e22a12b5d4bcca220dc09de4eeac3c2670002a40c6ff3c185294d3210db667da9896fd4f4c158cd1ed6150ae07c89872fa32b20ae1a6becd83a2e568d71c3c0089b441705e94d74124fad024a324edafe4f5f8dbca18bf5fd11351b8236f798f460f2b506640ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h476769a6be8671213e3caec4886e5ac55cef16c97bdebf5a6c21ffcc1f5ea3f23778e8908da2660658f57ff2cfad68961f6e51d21162c683ee2c38d8807c36731250d5b940a9cef3b98fd5b998f5af3ec698b3e2def3bed09e1ea4388ce30529d00d33054ab9d5926e34097f71465f8de6722dd2162c7cb81f6f73511055bf57f16336c516a4153e2ea8bf8231e77103247d4c90aa01551f0e329a24b47562ac811dda1dd784db748aa18b00aa379ba53ce87df47198695b68b66f4809ad10401e8657379f89d510480b056d87fe86144b6bf7b6481937394b400c7fbe066c16a9d1f345aa6e96835698ac7566333bf5bf59ea69db562fb93059fe5a097caa8324a1027487628d8bab05d7516e726a843183c57ab68f743cc667392849f41ff14d58b5cf36a883e16a7196848b489b7b082b500d387e7dde4c7b637cb6aa6add49fed6ee9dafa54ffe9def8e7140ad7a05d2e73c0407ef1be4172a092c758eb2031a91971e07794df11d04639c52be4423a18f6b45ebc4ab4dd3109bd1c80a0137dd2dabf6f0080c2c02058261b9dcf8cefa4860caf72aee28c1875e8420289c078d0e019f5d454cd405cf2d9cafab1f539598f0bcb5d09ca587ffe7b117f2839cb89cf9bd8070e157e498594e80f20dd56a5cf3a1f97a0d131d7e1152051d1a09ff4bcae84f4b63804b76ee3f0210638c427141abdd4f35dc8ad07473bb013b27b12c5623e40b185b178fa3192327e9630f9667ca8af30725208f1c1d324c20695eea1c73dd2e2f21611e8e61b89de294e73cd3b9aed5285b4c784904dc9ce829b4c8aa747dd6063b7d66197cf0119b22fb69b7a35125385079a66eb19ee46ee27d1c9996a5279c94238bde000147fb93a8842c1a0f5ccbbbb45d28a747c93327c54043258545da042d8d9b4a6968014b97837bdd5fa9f283709c6ed6b596bc6ed023bf2f13ffcfd06523b33b7fb0af7d06fdda7660f476dc722a6ba73ddf895c152251063ef61f56c0ed38e92b4a46a01ae1ce9827663c0878be0eeeb4a48163c440b9d6b18af40cda3e8002e508b242125b32e7fa5e906867475f8b540901f2789f1fbcdaf10014f02e17237b55d194d648854c5c7ddeca4cbba765436003635e449e0c7b22653cfacd86293b20a97d8d283e14a8bad2ce64e6f82207648965713ede1b97a27f290cdcdd7c8ef8e4d0053416b176be461b431a0221e71bbe54fce15b679bcd3b091666fa27a2609a7804c58abd668410d8870f1d24dd193a2ca8086e18fbf32284b8f02aaddc8e75a9391554211b43f37fcf32f3785936967b0ada99cba14ec017782e08b3d90d1b6d8f37275f323df9cc08937e71ecffd518bdc342d219144eabe07116dbb388b53f646bdffd405769d0d9f8a6fa044f17f41b67cb64c1a93758de7ad633c4937873be5dd139c3a4eddcf5ec922a7ffe4c318af41bf5b6288e4bf72f93d6dae7cd9fe8b55e51f42a40c78f418f1b420d2b441d374df81c86eb8f84a68d9727fb237b856aed19a219af8226dd1a66e8dafae995ac03967213ec0964b435ae37a9ebf76524b44fb18629c6bc2427f6a8b4c69f6dad442d5411bc145be5e5b33c834ca555b1af9a1c531e905366de0551bfd2cfb16f2be79afcc633d249d47d5abbe9f4484b7d4f1e8383a64ed5358f3d8df6352810a985b4419fba66161698c8a9527a9fae49707c43556d231c8fe5329be73586949616eb2a06010efd44bc91e7f0baaaa315b5a045bf0f6a634ffbca90cc8bc414acaf244c4b5f707121b7ebe03b7caf34e777e593ea780b232e48833dccd8a2a3c6a68627cf5a82fa2ce1672e3a4498ed24e89f1545d654d27dad48c45f4e091cdc7b28492365abbad3153c5487d290a2845ac6371890db20ec75dcdac1e356e78c9227b5ef05b372e8eb72b343d36b93e8c73098e3e4f79bb84455994e43e0ee28425d6969a15ad03c9f038b04d9da8a9f8c2fe8bebd690a61b0a1af7d893e9f1b0d19db4a516f6387b757101d5cab0d2cc9c07dafd13cc3f301acc3c88b84fbe90c12b0109dd0989be6bd200c4a8fcae5fd9aa9981d38b20131092423b1630b8c323c217e0331ea94fa41e9874c93b9babef9499f8e1d2604e88d0b8b69a43ea89b5a6d3e804ddbdb06bec593440a408c8e7e8d84cfaa8609e9c122ca6e8f65f8df912568629fc5555cb3919b63e282e6003eaeac187f13c60aeeddcf5c07317a3e448465724a116aef76644537a3a806b301d067a9c676e51276a95d28cec4305dff84d637729d1ddcabaddf3dcb884bffec7a59d99b306bd345616d04b886a0a407699b41de10580abe89b29aca9d785afc6d08c3091383c92556705c17a744a343cc7bb864cd8a0d39d42f1942e7d7281be92fa4db9cf5e679126ae53fcd9f4add75e744aab08f502210a0767a140c83f2aed5d4f55bbdb67062e005a00880bb8a401a0bc64fa70b27b5800a11471d0d13852c4b449033dc32bcd23bc79f53b6b5d1ec206b90d109cae1074de7777cbd8ad3a99b3aee079c94b0af720731dfb559b43794ef6a1fc121d588b7b800699e98c092fda149e37ae3e04b4d4a79b6c3c5d53e88ea88bdda81345f4e6f71b9519e5f776bb84ab37f7a285c06887f478e1a8987f27cc5b89313084e730525c51ca5daf59ed120ed411e7468c2d1629c4b5889984473677da100b55b66dc68ff0ca35a1af7e0f387be2d7e28df61bce7c271de74dcd4b365d44289d58ee5c631880257e7041b9e55e2e2b0040e0a10f87c862814cf3afd6c33c86b0bf0576fe0ca5844728198850ce8813997c2dbbbb81ba72efdbe6d8687638a11452aedf3b256ecf1d09e03cf1efa89ce3b7f082df4f26b113ef1cf764737d7e93897100669b60d7c963e71aa99de74c44f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf72c49aefb99a513198dff459b0d17d7dd72853eff7c64711a64b0e047da3d53858a95a647bb7e1212d143f63d84c28277abe9899da3efb6a283be2278f4f13e718788c22efb812410e1649ae4300486c1cf15f0c600fd2d0b46cfe5c15fe01cefbfd0d41644d56d966637e19eb9575db15bba25ac6e90096b388b75688a31ada0cb1b4bd2cfbae47761d3dd8ba81162260724df9e9a5710b6afed673ac508f2a5d874248400ba7a4d9b16cf13a7bf6e277d259d9e6ab16d75be6d23b4623446bd967bc0ab21b50b40a978036a7c06f788472f8c486dab1f68ab8fa464684c3599168f2c98cca6347c656ce70d50a86c933ce67641eecb86d1e65b8f5049840ce5b117e6160b1d87ecc7344c573f2d87704c545e6528d8e65f45e731d2bb3e2303bda12dad78697a43e54ab566b94076bfd67b8201d0db1ca637d7dbb0624c630372b59ca619d3d41afcf6626adbe54a9cfb686e082ce2210ab1bc46988156fc2f855dc99698aa55322621854fad96651a532c8ce94c58b86a3ab979ac85e09d80f492e50a01e3e4633f691a5e12204b39ebffe6a3240f6a9ca51c12a7295a3c06e98396ce7d7f9cd663d1d5f957d0f4743aaf8044ee95c143cd330a7504e891df74e9e950d8e7d5b83fad73cd19bec526f1b457145cb2091dfe1ffe133acc1c61607a14dbd8ae6915952eb8a4c63d13fc5381532358418d28ce7809bf4e0b90a15785a124de9c4acba49dfc2f7fde51a38671cc3e67eb038fbd3667ce307964f2b9953a5a443795447a1f7e73f5fe754813c369fa832bc0039d68e0d990b44f6a646100da6208f6cc31866f34fccb042c585e92657be5a04bd73e3d5c83b6f5234c6d502b2a647c186b8b915b890d503a6f8cb9dbeb361c916390373a9aa516cf163ab98da4f1635201e86f9dc946a8e0bc4e4e04b45612851aca7c5ef705e5f3ed3a4bab56aa3ff26a3430ff62e37433f8d81621252d5b1faaa975dedbb1917b2069d1ea754e5fdd056b1dac64f781b6aee2ebce386b7a365593bfc1f94d5d528560315e3e6a4c83275b203d2d4e9ed1b99ba5a22c048afa71de275127a05ff4a6dd146dbf2a8701c95a76a6e60b75497eda2370d9cd6e6bf7753357727c28e4e5d14e133784da9d28d769616f1dfa24555e7b2bdcc80e664d86ebb2cfbd663e6d33259cd49c5ffddfa9610078b2175f5df71917b32f8043f983dcb7775fa0cbd9efb34e3bfdb0bb864daf07d5fe21ba671687f39c17ccea5cf3c13ce03d8332ea9573c5fb8d35f52bba561a9bcad9c45082a92aaf00dfc3fba2f2db0a5d95617931f134c7149347857ec4c9c1115001f800a6dd2337efeec077763e779a6765be21f9bb0a050bce90de79d93412871913ba9f9ae07859942eaad239c26163375907f5ddebdf5f8e41cd62e453f72fbe450f63ed6abcefd57323cf27685cecae68f0e5f565b8d64329025eecca11602747c907ae0de0764fb3d512127033acfbaf4c81cae9a434ad075c4a9b4de8e5ed884b6c7226671ebb45d773d72765a8090d4697cd2bf9445e14a15e3ca4c803c1f649aa705862c8e5f4a516a670622991403aa20c029564bffc42825d9c21a96c1dca62fe8b89cbb37c31e9e98c7dbd91a824510a65bb5b1a216739bb8a469fb259493f2fdfb0a7c95cc76b7c999f44c3d0659afc87a2e491ba3d7a46c3d16da7c11270fb990754f46841a611c9a13b85f5fab6b0e76e9bc77602bcbdb8d8e0d55d1df21ea12b9f742eb28b98c0f444c025f03c8757e8ddd45bb5fa35fcf43cb8eafbaca3fa3e805d094f3d7c36088396e074e3463f355f75a8ccdb610c20807996cbcb80cff4532d399941110de3a0319240d235d61bd6abc9f38a9ab8c5a0ea30ac933dd3705f1cc5cbf5737251de355e1c7798fe7c1b2147d2e7cc2795bbada4f998a9ce7a93384550a3f25a3a7409b2b8cf8d4fd217a83cf14901c847048bd12d586db927b4883718d55b9036267f2bb7969ea17ec503eb2f0aa113e62c881f9bae51531021ba3795baa9ce2578f9c08010f782a90136d34d46fd01c73014032dcdf111da8f37c78f39823687e36b22bc7c415d7a581bc194c3aeeb3a4bdb7c0e4e04be62ee90135b42ffdbcc6d47330e8e8e2aca6066462af6f02f17bf9c28af5b1a69e121d4d7945c08be133eb0ba9ca9650b0a7da973eb7cd618fc55537028f26413443d7e9769567c142bec93f8981aa25f527de26dd692afc1c4e63f8122f909b59c3d86b48cfa7e80ad18ecb3c12fff4d7a968b1a0a420dc91bb2bdf7ba504a17e98311d67b5098305b4875a974dc54ac465c8059157f694ca7a0f1e4e7cbc556fbf32013ffc10f3f9d8a6842eba2a4261c0c7f371c5ead3c915a81eecdd6c84aa68555ef05f638b10ae95544fdfd024954e8686ad0756a36fff21d830319d6968f4070983ba793f0ab8b799482bb1d41a342e0b40b2304ddc80e47e4c3516642057d43b693525b5dbce1fde2849d5a8535d0296933c74322d3d663fc8489065cc84bb0abb468336af768947a227389a42f76793715c01a4227015ecb329c72334c7675a7b505fbfbfede65afa8459b1fc54d983b5a81844b78699ed20a24b3bf2c01089d200051b8d040cd2c4aace45972fd6b6440f9fb194f0e84afce48a7af705ceec454dec0b263a654123a52b9a9f94ea6eb7acbbc1d8258120d96bac22a747c98a4015530d2642542917e09b5f5e136a57e551be7266232618d86d289c6fe59a6078e1440ab86d7f7a21a8f73261b9f305a33e7251e33a209f68f8c03715be346315905881e9937c76b5353fb905fbecc837c93430fd8972157ddf7a95ae45a90fe6e1215ebe8b8f613197bcd59085335861a29c0b17b5f6a3613549cce8b438f5b3e130e0619b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfc43c68aab7c95a70f467ca10a77ccc333330c6ed210c5bad999da657fe6a66a34115273278360ea0a60c2dad3d17e99cf350024073dfc75074361f517d7861fc98e7643c04e3bc817d80a7db6ef088225262d48e41234a8113d9bc1fa77b5a9aaa01d6f12961c0d86fd43bdd79676db8d6483ae6d103243e80a6368860621a20e60c43c44311037a3192ca9f2c2265aa45ac58c1cebc94e78a47c20c2bbd7b2a79a3090798e2871357c726308afa3af9b7508170dc2ace39e8b41384f0cfb1ac3670130fbb83d252cddb0ac889a5c239622a1b9d0bc970c75bb5967e442cca3d339a319fa713f2a8612fa34d989c83e0eaa6fa26d0d5311c33af3bbcb1f8b6d865e2e1dfbc657194898dd2f0d9a9e95abd64224718547bde362ad398c231f4afe67b1e0609e6f4976e5bb82f0d6c7ee3ab22d5155d22ade8b15b341142602939be66d0be24fef25c59711732c23ea188bccc4cfd5655b08b1c8b69d53a26361a40ee2cb89f0a6cadf61dad32df863b07df385c81a8d84ff4554ea9176f7e379bec9cf7860c9c81a89cc1f33292a1379ec17ac8b818150921989a4994bca637dc1a8ca74521b393a145e72ed977a0d16868d1ae022fb36dc346c4ceceb7f30e176b9f6ce348f49b6c88dfa69bdb5b3f68f9e64daec208b76fd3068faae4d354e96f5a70373d559a69cea6f07fbff86ecb07b86773f3861f067527e67324e7d377feae1c91f0a644fd8a818c1e0b086729f0fa7526b262c17fd4fe563dccdc316e23b87911476a8b3bb729550a916a70b9f8f09b3fafb9e49d9fda07be3b8c732b1e9953c95eb06e0ffb72e73d1b6225a1ef79759fd03856f3e1389df3e4af7432f913492de1a55183931b53e08a4408e05bdfb11b553c757a7b9e37794021d9336c70f27ed097b1053ba0158ed7b0aed232d6d63cd2a250d6af3ce1e8a02c01730d902fb558105a7515bde4fe1f6319e0a7f25f31611a6f440bb0d432adc2050a7ddf90578e66c921bdff6115be4673d673b38dd7e9b2ac0a91c00cbf21c27aa973cd308df143c6cf94c8cf4b7eb98888d276bf25dd5e438c7d611c395530bb025b265170ea23603a3a58d661db14e5fd7a743a95c0551df12aae79226ab67701d757edbe503932bf234bdfd24ef2f27103546df9b2bff2c7d18091a9080436b2e48058b19cd00432e2567c648312ef7c4e4b2c1a24fd7e0177d8ab7521d9543f35fe2bbbdbdce62b6b61f268d72f9372fde868d8a1c8f4b188c18af7267d111dba3bf01c24c3cd94adcc81e851ec028ca6d5642e2c325daaad4109301899c7eb9498c24aaa3409eb1325e99ba4c7de463d02117055e347af8723dfec847141fba0104e254064e8e54a213e6ebaa9e1e0c312a3619737764183514caaacb3c79836ca630b57df7077b80431927d101beffa43a3586bef2673922c9bdf6d38273cce2cb7b0f351e1817c7d76215e5571ed11e89e02b1d7724cb382e93dca5ac8bc0f1b1955aa13f639e56d63ffd5c550c6542aae8e53de13b12d5bfeab18a84ad95706b9668cb6070ee086aa81a27d497d96b0c491c4e307f9830318cc1e686b6ab3c4d812c7a992e2eca6d17d5d54ef677115417bcd85bdec6fab717cdfaa6eafca0e565c1cea17230c163932bdb82ba8452a22fb29369286bc80de066dc1f014826d6d0b818590ea61804bef42774e511bf7019a81cc73dc1a470dae00c2b03a679e39eeb1cf92f0b22331285154363473919f35dfebf7e16dbd11b4a3b58b002a74e9edac0d561be6d31f75e89cf44a9713259d3e3c54119015e0cd7902ac8f10da1c6c1b0ecd6039a5657f0c94f446cbc83e4a5127292122a188cbb82a2acd8853f97246e6a07380f26f3ecab956c8f2d8a09260634d05407121f2f9f50832f896a23b498f55e7be369932fe8d1b19b04a280fd72ebb23125ab7e10a6c59aff8a54638a8ab4c38b0a716cdc36a8fcaf9f2edf44358427fbf9b7f56db26fd7df4f55342e9a58794e36ebba2f7e3746aaedff4bf4802a00310822f1e4cf4f456d5bda245b97d3318887e1346f3d62359dce0cddcb1bf1d274df9862377e3d3f72a3a2cb47ab2b17cd1f1748212bebcc9895b7ed3e7bdb3675d25d0dd7c9dc155ea0ac2ef6756e2dfdc4aa53fb1a0a0657b9f5a156360f4aa8898242d761c1aa3e820f384824e117bb79bb0f2db048e221850d0ae4866eb42382089d5c6b3d1f610025127af7a3345ed62a8425cea402338e74be681a36af2b5651040c19baddd23968507703441668be06f50e2c90629ad2d739aec022c2021b086a821ffd0cf5d1016c339f09b6d355a65021381c5eed38e8568f6a37038dbcdcf61ce2d3405fbec4c5859329db51e9cac7fd3e9523f57eaa10da0d2e29d222f46ac18427d19507ac91f42f4321e4a4ec2859f0583ad9c13d68fd9ca60446f693253381b7441f28070493a83dfd222fac369c8bb8c42bb0b3d288191224000d4fd99a2481e93c34299631e0550ee7559f689e2dc46910634e246b9823b62cee0788960c1845fc39a2c5567eb095fed3f020735597175a277cc219644929cbfaf78376966cee23933f1ef31273da8ec6afddc992c6825f7e461896b6d7a063c5376d712accc39578bb01e13600302ce587da2bac89e51329aaed110716e89cf1563e50e503b2e9df6132192f55511affaf0e74802b9028d76261924a3e5b84987b5cfc21a62d5197f2dc9917b1df0f035fa29f912ec328c71dd3c05c4997449f02ce4a8a4adcaa5356866ca81f7f394af45085b49baee40f788ca89ad1e49a8b408ca3b8fb25e395184b11ffcf48797ddcc409a3e4567197dfa6ae9c230eb7e8cef291fd63b5648bcb2e2dc30b67c161444b5783d517c250a0905ab2c232298f215cb39a6738;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6ba581d5e3ebfc010eecfca2e941e2a16a74b13b765899f2350bab4ec13ab9b8ca7ae05a8abfef7e26afc0239a787373e61a0659e5ce4513fa359edef9d90cbbaf0a7df63407379d207ee4a028087153e5a6dc543d448eb1f4eb377eabe35c78bb510c85b1f5825d8e24ccf0fae251a2e650b765bec3fa1f414dc271074480f4156233ffce704971e857ea9be22aeef2697e075a2908083a6d9d32fd8264c7530ffcc409281f1dc7e2ae4cea10e5ff1581139321915f7f969ac561e21b379acbc9db226875a015546768f16c9f7324c482e02a2b390a6df3ea6868fa1ba9607f6d4dda2d903ce06022511b0becd598bc10660469f796330a1fea2610eeb3334cbef4cb16fac63ce2b50f898a74865348cc7c942bd118af1916a1e863c83fa3822cdce3bf91fef2dff44c93cc1ab4299c860258199876887be451ed8b153896add158fc187082d41df167fb0836255e65c50da342496dc605dcec177851f0fb4d7d1fa7927d43865d3c3f885ee2f34293c8e9837ddbfc324a7d5e80c5c11466db3fd1862d958b11ecbfbb0f09cb5864dbdca0f7881620494e549ff20a8934f0c8baa130ab72cffdd344748452510a70b401e67af6dcafee57fb429306f682594ceb0509455797bb03a3f3141f1c4034c8bc5b0598e5b15b55aa040a65c94bbf2451ff200bd8d51b82f7825a1c97e94815cbd27dc40b5f0155236105faaa1ea57ffbbc1d3ebfcd5b98d5c6a62182fb54ede5fb37f20b93f272340855178d2c3f602eaccee9cd438d00cae1b96bf77fb4476fae75f8eb445ebf1e04657c4128624e989445806de3e67b65b869a22b28f0b57895b493e450d0e554f46c271b9d1859cbceef0192933e166ec715c8864822da1f7282063a906a6be17d008244e027885c821a1b8c1dfdf32124428b81e8849ee4a7298d64a63170e313cd4512248821db1a08af9164ed8e1eebe39382ce6f96fd66e8ee1011e369f222fade59543ad75ddc5230d03734f6c20f6c5e5c940b10fcfc290c7f9ce83903fe9fb27d266717cd5168064288a138a91348975bf67988fff77f65ef98d3820aabb52b205bcb8f29624cdef772c9eddccbda93d7fe530135636a2ba293d83877852fd36687c5b987df800accd04732ed75114565863bcf1b2344c19c312010f057a5cbc7fa97905fc7ba7b35f3b02f24962c8f4169a5a2c0ff48fc2494f6b1463ffe686709666e24ca2dea562a9901f49cf2b2d12b0d54256c944545275de12acb9c4720c23ed870c4e74fd038359303b51012e51b065e104eb875abaa58a774fac40cd27f688a0ffb80111982be28b47ae19982700a5ba1d401e0d20e49080a1a1769b70531ef05ecc3cb6b729ae05e19333890ca0e2cb7d14578dcad5bf4e568e1c4afa4a483bdafe6300808a0e5b62193a88c55b0ac30ea671bf3c6f78a6635296f6ecddd3972a868b6b352318590c269bf757761883e1f0ba5317b852e7d68bfb83420cd3423938531b10617ad19caf3d74caa3e2445b9fe4c43dff837d96119feffad987f43364b1ce6370819127f98a90cf93c0cfd44a01cfb5c1acb937a67a7fb16ff88fd52df63f8bcce7c3c696f1aa2e71e5894fcef8df1f6a03b5b78f476cc77c475c772900ebc1a1301f39142c7eb931acc2832a48eea9ce66252fcd0987c52b1103f3a8722e4d36f22b6cc4e35fe3aa29ff946c40b75ba76927feb41c984013069c07538dc07c5509e58d07d67098c7592a33a675509611ce2d3292cf5fd68c1e860ae93468c85af4ad3db822eb9a971fa7ef0152693d3ac567ba392910307b7bf7201fe73b08ff292139be5ca1eed467b3e4bebaa6b794ce7cba6a13e81b6dc05a8789282ceb050383f0adc8e8d2103f9218e1cf9f402b53f0c068136b4cc0f1292e4f941b11eb614c6257e32cbf5374a067dbd8eb8483fdc0857575c90f9794128a257d7db1f133d871cfba3ff9652f3015d470614e3350f0a09caf65cfe1e2e0a00c369fdbf2a1028640ef5fdee141f7f1cc64c4a0fb1c456cf18c04421b67d938dfcf7038df5d1bc01517843628daea24c77b8c719c64648584901e1c99271b379beaa18155c98363ec6289a6bfb18bf2e455ae8b3c8ce779d2505cdfd0526b5f528af1cfb90c242051cc16ae65520d2b84a0c2bffc308b387a5afeafc570f9dfc4c97cfc06756127eb42b37315e09eaffb42dbca379d938af68da78646d81286d67608eb5507439810ccb207061b91c038736f8c65f4a87a18c43aefb00075994ed3fb7055dfd10a4095078cb4b46859032cd7a96f5149b213fe09670da00f7a33e156f38033d9fb2f72839fe60f1f199acec8e6332d14d3459a1ea9df78db591db8440c74087d4b19d8d04d21a649d5b9eb8a87d6699990192986b62ba2179161ae4a55794e68735c430098918069481e7110c62b25d3cbf49dfb4cec2f5ffe649c8ecffac197187d406350cabddfbf5498b4e2d6e70badc951a3a77aa0de4d5f8fe175fd17bbe4d54011cb2d02d7b9014a71aacab5656d521f88d3a533393847a549d328356b6bb0c3f3867645caeaceda3da68eb2dbbb6158ff10fc78214157cbf10e3b44fe5adeb7330dc5f083fb30b23e33552a46226dff6a45cf7d5965362950086be66ce54a97abba490e0a7fa42718e2c87bb6f5896f3d56696e7568becacb35785e33479ad16951c2980822a65d0c76163c8aa36db76a989c1e8a657027d854c503fe96c9b9db2a719d9e96bb38b501cd630b804957cf4cb28c94f2ff0988d859ac893ee1d2a8aecea3b68ff1fc5bb711daf4ef6f4af03b907dbcd375672a54221dd0657495eea84b0d63fadf5d2ca056dd50fe32941e4f0cab0e7617334e4fd1e9944cfd3f6a1c8001a614b5f78c88d23316d0e19340e6151c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf21f5db418b0bbf8659ace253206771f278d979064e3a04246ede9f36587eda11202c7a3e934edaf9cf6bae531e61ed400a7fb05fa2ef8498946bb6bf93841432205180f41c4bc48e0f92955052db5d71c19aff7f991e2fec25c3a3f39d92f87e76091bca5fef65c2f5e13f333347f82c762663bcb420e1f79cb41dd35605a5f84de3329c7fc4f9ced14f9f6d70241e98cb74c2f7c71a3a44c544b32b7d63fc67c6adccdaf7e9f431a210face885bfd42be24f1f0acd54254797bea35a5bd915bc853efc4688169919c3ef888df1457c9f8f071643dfa8d29b659181acea436802cacb1572ed25b9620ff28c93a44365fd916db616922a7aa763dbe70ce90b47542b52db8a081dfaeefac3d8096d0db6f1da73115dffec703cf2b28f037a389937785fe15429c5948bac2a815886949ddadb51677a2c71f1bff4abbc1d994c19f317a37e64086ada945c08fc98a5221e5ac0548a903dfeac4a352b9baf20a72e3220dea7fea07d7169e182d1633fd8b3d344f6d2919e5346169754faf014f0d6f96a075ec7365a5a468636e1be5ca43302cc8f1b5563d37332cfad760ffbcf3d312aefa71cb59aa88a8046433e09b9b191a8056226de4621172dddebd6b34638db08008d9848838e269b1e27b51acab217e0773303438df2509b88f50fc90ef03691c6a9ae2fb96e423b114fcc38dd6f91b0ccc802356bd1beb0bae71db7c8d5294cacd85c9efc85cf2d905a9f59230e932ac6e4dce673f2a5867a003a9569942356a32ed9fd2dd1187bc77abddcd9a7851c93625811a5bd03c34ec0a5994fee4fb806f72a2dc86e496e04dcbe84a87dc42d56932d0607c4d12ac7808316591a644f348a9d2a9d6e7c2e9e7f0862114a368c3a8ffbaa7e03f73f3a09319bd7f9f97e5c8532123c8f03b306730c68e4c6089d0f3fb011f34e27759e42c9d6c382a59157b7079e4df58420140bd142a028be26282f4e7a90b6cf5cf4fe8036ad49259e457556700714ac33753d42c284298c24cf36ef946d24466f26258f68baf61d51552e0ec9511173b553919ca9f1b11edd90fda2d5d7fa9c8172a04b212a61386ac1b6303255a3ddd86f2f4d2993c158a20d5df8ec9870f915311251bc89e27c86980600bcb4422a43446f9113f7bc2245ed2220d41ce16767c6cf85389e76c7ff647d461069f9cf607c70929203c32dc4848f43be41f8229b5bcd6b3f4ac1fc6e708a40629e9e5f8e5c69fd256c4c3efcdafa02f78f94bdf6003a504c2e10d6b34a27bae2a798e9edbdc056fe82ae9acf455895b6dfa54b1e87aab79635270bffd669e8a4a3eff4c481e4aaa615b1367e4146db1bf96d31e3c5cee454598e05a1289d0939f0ec9f67b99500ffdea0ab5dbd122c0b5fc1588b204b35c16d603e285df9cc854a864e423ae36a6bbbb4243af0f847703bd9043bb9690d5cc59d2bf443b796d269d27c04b6f8cbe90cda3f7149bd0e67b9b87086230085dd925a3d8af325ec419becb4e817b17f4ea40933cf1ab0799fd073f23218a03b8825304c7ec164a7f2b0d7c262dcbc0b1c9a34aac41ad2175c8672c7f88584c37705c9433ac3994618d2c5192f4e75d9db47516ced4c6d8d10ee3f25495ff53f4c875589e9963f909225498957759733c73d8bd447e9e1af5d80d2f99aad3621f5297d71aac43fd3d0ae9e6466fa78b5ab94fa81fa0c06c452c057780175b808a6c0518dcfd3ba96a325a581f9d37a4eca17897f2e1cd654043a296db04903493feee5a927fe153448fb7dcd7bb7bfc2a6771fa6ca542e761cddd9b19902d0bef07cb343338a73b41128569d092d1f120951a04fb5e7843e284bc66bccee77d4e0158cd4c355e7c6423cf435bedb668879ba8985126a17d95974d939492bad3566db929e1b645672f4cf92b78ad0227c7f2a238d91a58cb98619df682bb870085fe563a1dfab908a5ff9f73502dd6dad12c0507f08d32452985819f8cc493f585e993042667f66007dc4de63dd7c0313a0f1547cc8a64e9ed7c97cc5daadf99dccafcbcc4c67575cda0458eb2b2b1d3d3238311bd2d726ff4a6edb6999a4056db1ab10c2a0d3c448abd4830b03a87c534574700b0303e0ab270340a02c007678b71eb2c702966f4fed6aa0240de8641ea342c01607d2bbacffeca8655a6ef27e6fce6ccdabf1cd960e481dfc69f5ac042248c84a4e411bf001967e7c51d04b514ddad04b231e9b987b5a2e96ea160a83a803c57c2397b5f26c544340e71de1109566ca6436cc5c2df350c5222eda6c952a300cae6c4feeed56410dd11c9f1de8a641c795d5eba04bac529488aa116df14e25fae94b3ef3b0bb1e24d08299793adac9bf3e7eda1821dc345a575365833cce960fa1b5547ff1c8f00b628a495ead1ba4135916d7b6f2e185ab69e5f160554d33ab1dd1358933af7ee21c2b2a07cc3c39d09b2ef9d720f623af719c9ac77698b2582576f71f323cae9e30d41d039db81106b3e0ad0f489d6a195b87c1b320785ba4af9c161c7b32f9410acfd035dcc0dad35c430421055ad5952eba58722fdacdeff9948e152506494f808fcedb26345432efb6db77e881804c02c36115215c062576008270b0f5369e8f4227fcd554d8f7649070cd9849384cb4f0f87ce50d3cc56d4f5c70717fbaa76c62e7b1f15e90e4667701ec3cc8c0170da816505106690270371e19eb242ff952d9038152b39b2f5d2e2e75ccc81949b84fa6505208c0ca47d37d1a870a8948b8436d773e2ab0b1080fe32a9938fd2e8bdb8563d03e6cb95cab18ba416edcb9d8ae3b0fa0507d3eff5a924ed40406fc94a8b7c302c992a71235123747216551bc95b4052e664ea066f562baccc6b1cbd79ab7ca58d16a5b02069e0e54c0423a7ebd8324674dc710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1d1b585e02a44a515876a3ff96874c538083f91add58ca065eaed9233f1e58ae67e2ab77fc49b6f58e46d75b16967688eede458e0df71adf8548854d5f39131ed796b0ae64d384e2c97d011701fab9660e206fe8f590bacda0f5fb6f6df468fce3c98d41f4bb1efe30f6a05dd0f4a307a84804696467626c532e32e747c6a6be1498c7b267f82fc90c4db1d69333e777d463c03d7a82dccecbf9126d28fb1ffbc93fe75b950614037064a1da3222f3a9ff3b054e78360504860a2e83b6622482c0da018405cc72389e152ae16c95a3f7edbb1d50c1145165ba9d8c5dbea5f6488e8f6fc46f8a2befffa90f580f9889425ce8d0c3595a65c56a4076a37eaf96a4832a73f88e0469917f5547f62e39ee931f9e7a7135f3df853b2303cd6ca0290e34e8f51166c23836d9566d3883141bcaee0321cb230ed4c93279f5aac0f63da81a04278d6a1ddc990438fafe1706723b37d690c67cf5472bcbc083afac3b2331e3069b653bc2cf15fad739d44f74e68b31e284a9100071c00405db9e1157abfa2b27b87a4b303227e8dac83b592cbb436ac694b19e9601e9a47340ebc84527869959102a76eea453358ae4347fc72ad21ead7753fa69022aa2947b760b6cbd6bf38a980553e9c28d019f053557f796f2589254f5f90530fa1e56ea33f740a3e2e9cfe26da715cbc09033f8039e3c6ec5ac7ddadc0207a87da193debd28ff86f9983d1bbde0e48ba7f5722fe2d454a8e33a12ef4076a789586cdf8cf9531cac866ab6d871f20f9f9e3a17cb2bfc2704e29efeafcf3b2689278d73745827332eab5b76d539ae9960fd63bc9a08fd0f88615264ff7021ffdfb5c16c580a3062a39f087ee2177dbfbd2553c2961b55b422df17caf85896236437318c8b7a7987410fffdca674cf29a252b67158e8094f62365c9b4bbd6920ab820d84db7fa23edd564066b1861fe09d0d25e8e17214ac6c824e30748af434e0137d5a2c61c98f9ae11563aa77e7473e7c8dc30b95c060a792309aacb88a19bc48d32e0f9d19f0b6286de835ec7a8be9c10e101192d45460d4727861aa5a1b2befc9db0d3250b9a30e8bd099f97edd89a4d99517a6700b8a1ebb4e9221dd70e015b9b7fd1875d2becc82abf3c5ee467c641b8394bac15214b780a9b68e2768f211b49010a793c51f14167274189a18b93dac358ec33caa83a6650aa9831cf279658ebfd78dc3f33793affe2e2fc65225a1e9d84e22449d98d95855cda870dd2e839301451cbc304d10f8f8a3c49dc9c256c68c4c677a2070c93bcf4d880a3c48c3f7b663d1236e1a619bc700127cb92d4acd55ea2deafe87d0cce77cdfa52d5947da08959db56383c1fac96860429be9eb93ab15dd19216c2f0f8e15e9a9049fc5837f849694b2dcc4f3080d073091a7e1a5e0bd15b21d1d8d2e6222d94493b479a5ee8f5f76535f14ed8d0f7e200e8b3414c227e3d0ef5db70483711ab61224c4cf3c0846cbaa180561423999bf540dc35444d29fbef52685cbe5bfdd6fe574b6c9834c1aee891c983a549dfc774d4044820f11ad3a2b181285492f5f764e151ac0d3656abb8f8e52b2254b47e1428d6fa6409a1d83e737d8822be0f5d2887af0261e74e34a377a7c94c0d5d6bc35fc24d6ad6079c0a468cfdc23bff3c7d39e178239ecd71a09f84c6f89525e64564fcf54521c123f2a01be175521c562352314ac9764f2905111a8ea060906bbe099a0cc6065a308f33cb929388d0d561135ebd57bf2faedab6b7c4d298bd9cc0ef2a6463d7a55b1d37dbb98803d0addf2cf07b38c6f8a3c3c3d61499a2713d6ec8474480882c7386316a01f1de1f97ecd27ff2c2ba77c81cb34ef0b999b9021518e95e4c8b4a70d4b3112d7a825857b0b941c60b29e855288211f896d036054cb5d034332d5e1e33d2f02990a18bd3eab20b47d2490d674b705a861ce3900995ef78d3a19ddd05c6629b8a224f66dc6092246103d7026d2188e6f004d262a631adc331b3ff0554f94724576254fd3bc1a214b641f80696e022462e107463f6aefc29e49e11098fbf48a1c186cc44707d004ea88893993329639e50965c9e9fea969d5a307eead1a9820b1767f05219f14d107fdbdb7fea7ff1fe31f094718d0d4c7149174abc358af81f3c16822c69cecea33a281f26c41dcf05870c5a1aab5b311942b6862f7cd44b1c46393e81558a236a190d3b54d32112f0d4e7f27a5cdbecb80760e3581cc690171bd49bf64040f2029775fb056afef302bf61031c9dae62eec7361ae27af21f33d0425b62e9d06e4c6592f2d7e0fd1780b5ba19952191c3a208efaf261fb810ddea9e6d8d36d62502465d61901e7e34d3cff58ba77dba00390d0788b5fdbfe542ee63ad2a1f17d20f10054e206ed1cea7e69c9e3e69c2a45f84e4d3af697a53338c513a064d3ad599fdc1f511314039cdd9941468923cdbbf7f0be726511c1cf2fe621ee74a1f4986588ee789ee399384967ae85a347d2f2eb43fe24b603115e56601f31682bdb0e40183fd043ecbd7e9fb3aed7d46e462b24fd7a288c3da688e5673552055fb26a89233366dac1807dfb3211441f94f1553d3fc7be5d6c36f05361bc51f84eec87b9c56b39857d50c4ad7284896e2cc7f7dda4cf797c5021ed1564d01b63c7676ad17c985228ed45a221b5465a420d3ca6b84a430c5c51266a0bc7f6272d304876141d26b33de51acd2c0300162ad4cb8f7f287600595e3bc46291fb627742ab1acff12abed2d995be01fa175a9ca835d91459043d63b243242791ea83e34c04ce9884da352ad21de599db2ca3307474c47af3bc6897f258fd2d4f302e29a403f0bd1ccb42e5d6a52636d9f56a14d55429cffd7f821858fd36d75bb6445308070365824485a8a1ea9ddd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdb5bd138bc1200c58098792054c92773799d88a76cc29d3c8cf4a168f7237320371bf31124c3b98fe1fc8c6a35191d6a2d3e258aaeeaa4add4d37582a3d0ab316a307aba08cd5644318628b99e8ae198b55bba711d7398a61ff193e4dba6e9fb9e6c8ffd9eef5659ee6eb27263783c4284aa89ff5731907cfd12660ccd686d78370ad8423808742f46ec4849d9cdbb29d2a81be650a6fc2c2d316510b37f09ef223540c6565a2ae9f9a9d2d52e0562c0583bab576db646c05e73dc373ef03c61645eb5a5c41e34ce041d23c45da657c172311367ff2a184663c38da74333e699a7ae9ab9c6c46b75da9ebdd269ba059eb4a5cbc010a88e958e1814d6826a30809053413c64d1328bd3d32cf05983dc2ad659114049263d1cdc0e04972a07210232edaf88a13dfc5588a015656e9f990179b8f78d77094910f4817cc0208c5d6e2a2a053d0110ba2f6e6471f6442d572668438b7f801017a34f2fe2d458a46f35cfe0d18e29f12937111b691f26b0e05b0283d5c96701c2f7f7f085bb96868cc4b76729347b2a1807857b287f68685aedff9bf1cfee66c50ef48203b60fb16c242c9df6f06945c54348c7e60ae4bac2b19aba005dd3aa7ad79c4d24cebcd0ad0f573fa41b6bd1f369c0cdf969887dd547f2bd04b2676249c84492f1b9d99b65348bf13e788871da24f5481fc3554172120b1167a0ad1c10f54880cdbb521acb31b66a0c5a71ba5b809b9f12e6493b53687974f24df40d58d3089fa2150868a993c1da01230daf9584498dacbce79f7668b4a3a4c378487addae478f77eeda329e8975cc3facf10f01107c2398611ec1b5a11e8530000ab7e9ca9f7b17e0e67204a68a9c2ab3fba7c7a20f9b5a0eb9b21a6cd8c65f2dd9eba0d58ebaf6533a9fdd3ed89f34ddb9b7b85db8ca5938a441a5132118e049b3a35d8ed8a99539473990dc01de52900cd1e260ce18d9297f4871fed5fdbfc8e2ea667333512fc7e3b56fda5283c4fc23843599db379f8986f6ad42080a5ef89d77e67030b496e782583b9a4b801a4f99ede0a46e83a65037e30d3c79985c13b75f88cd28ede04c2ea0cccd60fc454881dd2592da34815ae924845a495a2a0d439231e6d71c6bcc67de268181606e63f93069295235e18da4543149373e0399798770e584f808781d2a19d493b79586109bda39737ef1f548c62901acd94b3963deb3dcb12e9b759848330531bf635179b64e7f371c0ad4ac357b49dd2e1f4cc0b4e66eeacc0b233e03baac960c55636a2d4ede2c63ba6365821e6b2dd39bad9439d0f550d9ee509654ccb3c00abb2a09bdffe0502828bc641bd44805e127d6ec68218525346eb3cccdf1e0391675092a3f94374c67687b6591c32cfe7de285eef7fa46a5ebdc8c1f90ffe799402e5ce6578a3f7106f604da1337775b0054ef2733070c55460e05fff7b4625f8d5beccb3a4210bdb53369bdf024b7d768e290de653776c74186be37587241c96b66b7116e2cdb408885b812b36ea7a000948db16a9e963a8d6a848510840687fe1c15cb0dc5d014eac7663347bbff911953dfb9192c37b134c1758b207abe04817fb5e7c7eabe6424e0ce8c3c37754769396aff518c294d4599a863b8f5c9531136115941057790f3b8922335fbdec4e8cfdd06445bb61ef812931b8d22ca46368123099bd0b350f9b0432a2e9b87776da409bcd2a05fadc3753afdebd75884ed1a64aa2b50eb1b897fff4cfec6c7641822af20a8286c3fb2eb31e95d343fb8f64768c15c9fd93454b51601a645fe84213615302d2bd2b176a802ae086fbbdf2a385f22989471609818a8d2a59112ebc6c534eb5dd9ebbdac4c6347a0d662a08179568f6315bbd99f1bf032334a736539bcb68caf709106f88456d4c9254abbe5ec0770a29f4d8b2503870d80b0aed4f626aa7804f014379c8e35d87a894f7044ac37b1300c7d09ad7f192aed99dd32eaa981d45c1ced14dc35028dd57b110fcdcf6a8fce02dc9d51960c84c3e761858c83bc9f84cfd8ddfaf766e3d5ba6bdef3d4cf989851dd6c725912ddd786e774abc60020f775b04b3276bf6ad547cd068f8b367b18d191b95fe1b8bc4f16c37095a1d638780eac730bfcd7044856ad419c341702f8ed68f2d1e886a91ceff85a6cd1cd911550f4c94d4476bbc280c7a519a3065f01903f1c97faf250dae2c5b16ea7bca2c3ebf57d99d8b8e7e3063985c55560f8e11205ca32b7eb2af9fed2471d6867220e0ce22b4dfb786b11df388935ac535451800966602e015107ff6311de8843fa40e419238619fcad2ed710a4581b3c70aa7227a9e7008779553ac2d60054f1855f027af8f6532793dba5fd32ab5a6319852d3e85b0a38f4bcbad2b9c323c58385e3a8caacbf1159abb0ac2913fc7a6acea5d5ea186291bb5cc3103f185e0e61f1bf28a3a7c44cf4fdef000fe8d7f77194cf36e9dba0d8bca2cfe5a4fac7a43bcd2f144e8362fb9a1ae6a1d73a2a20d42e4785ffdcf8c6a5cba4a2caef37ca90b6df7f69b3b9f5abe294d2072f3a3f4f80e31c264cb03cf475fb5b7034fcaa0ce805f3419cad0c382272f242bc11997a516a59d9360cb0082f12db86ec12d2363749d4a0f3a232b7445d0b07d66951c3c445a5266d830ccb05a4a48bbbf8dad7efeb84075e03d51326815f79366fca5e36ea05c8992bc40ea298cde1d104562b266704999107c1993a296294295e776c1f9cc0fcd677eadaaaa7716084e529a96cb28753bb4b3f8e58118af508956369825070c62ea4fd58e5b3600f40892e337c73cbd50a3ee36d2d3ce21ed2b2c71b398c62dc91c535dc434aafd446e31053045832a54f6de18b9e886c0818fa100e4dd2c80720d004dd1097655c72e66bb00666d5517aa2ffa1d8b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc61dc84339ad145c19e0d61fc6950bd0d22fe001b3e8d7880d23609eda6a5f263ed971f82d25acb709fd8ac943c6a56229daa946f1710f30e0a15f9375c5016edef80f329e121621c840369a7d14d78c9fc7deda968d5fb8024077f57f67e12e596bd4a562170c20bb4045841a615fdcff3466a45e7a7305f99638cbae44d2ed020ec7b4c56d7597c2852557b469b6e6498e46b5194ebd76fdc3eef13a476d7e20b18d9ded49e78b538ac237e07dcccd8ab8fe08f355299c30305b23f38fceed7fdd8fd0ec7aebeedb088a6d21137b1afd89f120cc61d32f6383e8874bc6ae6c76544f3ac09134a5924ac9544532cdfe9d83be214ccf2e7a2896ed14e2f46095793d4ff4ab9e8d56a9c8086a7a225f6a883aec09ce1c4f914e459a9b14e51a3d766598b4b2eeb812c358bb46bab6a0e4cd45dd82f49706fa9b7d65824d1bf32ef0c15a7b8f7c20a0a8247accbbb846aa4fbf3d8184f60f10f1ad1f87071d8a78f2ee3b5d62edf4760024dca58b9a4b5c9fcc2c103c4e5132225cff4b58bfcf070634e723298ff559cfbfc1a3902d5b781c8c1c3bed3e94f5ea461609f898acb684ffb43bc3b126945b6390b321c164a52b4e449c12d3e3ec5e8fbb8cc9681420529a665b4f27b269f3b9d92d095f6622a6362a5b44c05d81f752481beda3ef7b50581446d1f7cd4aa48ab89685f9de9847090f864da3769c491021e291af2807a2f56e33ac7a2f37760c7810cba6b812f82becf1f8e181149cd2be491f8fdab94fb58ccbfd774f7ab457911abf0b83a73aa8065cc67fd6afcdd5c9bed99a77c68cc6ac32f7ef8b7803ade9e3ef88ee4f3dbce64c8f20fbde76b636692eb10fcfaa7d7893a862c093618d4e077e88cbb322c9bdaf4d6c3b21541f18c1ea1a4dccc407ff605e419fe85472e30a1d3cbeec9ecd326a88ef5cd8a6d193aec9d4cde92b456a1b4d8cacdb60215a4bf7feb68bf02ca3b05e625e872386f24913366cd8c7c130a78e60632cad3d53342d424d0dc3b9433ebec22b8168e5d8a358cd8bbbdcd74d40e4ef397e545a575bfed16b491342467880046b202e00fd6093ea9268afb869f6bcd982c609e21d6613d9b0febb710c962f1ab832e600bf925c999882415b8875620ec2133176942008754105471d6411cfb54eb2f51bb88005a635ef2d3a1f23204fc93e445e0c14a99a04c4b83f7daa36c49a266d22df4f32a4afe1fe84a457bb8bcc12c59650f7d2d4339bc31b9f24997b6b60d9d78635c62d215bfb7b987fe83703926954396c615b40b24dcdfd76acfc45fbbce7302cb140d78a3c5199fcd2fb469156e2759164b8c7bfa5eb8b472e952b4585249480d93743bb0a17c7fb81243a58cfb631edea127017f6302c165412161430137f5101fe70c44f361784a44edc9deaea145d00fe60045c24850a43af8b023a924fcdcbaeac8e36aae9d82ddf7182727f39cb8289ad4aa792d6a2d0d411bd18e937b967400c209df3d50888a64717699dcff954f1ae15259069737afbd88979ab17f33629f58d4d6bca9f417e4e09708f0dab117da6917187bb9aa66d62cabee7702df53d18b85c57e6ad6c5cbffa72a1943e3e7f70eb6bd729d4862706cfb0ce5b600ac74704cf84868d75d2eacc57fc5c1dd9295a65e2cdb8dc8463d01c9c7c1e01940a651dca234bf9266e31d9940f42e80ec5b1c0333cdcd00f32b0413100fd13bb8aa7db31e4c7708c2d2922a38b6117ca9c7f57d1a7983d10411b2e4ceb550261f9b663213e1b47a0585918802be5dadf08e8b5d91eff4b2af82abae870c89805093ffc7b7e878f4f41a02e8624233ef5a2d2bcd3179fcc8ea51575da134f808ce25a40e968db58af1706113f24f3df8cf767b925b0863e07875e634f5328d5a0d9fa5fe9ec875f94ea0864a2648924043bdaa8ea3ce95862858633e05438a775fd29c51b0d21decf05162b628e442a67cd3c84fa38c2a3c6079366baca1ec79038b991f70864a33ac458676682ff6cde93edc5d4c86b94580bd017356ee01fb878717f3c81f1fdf59f1214c1784a85633f05a3170ab19f5cc14b75e82daab3449f42c1a69a121d0bdd63d2ba01b1ceb1a6b0d9e663189afa23cca78bf0b7a392018dede62c044e0b00cbbf7249cc8a9662639ae3780da74f6d36ea8dc4c6cd2140aa4cc4ce3697364c56ecae0386cdec5129a07a5f62d08030870c9f755767d4d64519852ed741de540007c23c735d5fe35fa6a701abdcd4f895e6462515c6a4332e7ed4c09ebbda539504c18815736e31e4785fa81199686de3e1f6417f3afcb54624025bdd1a95337b0365559a9aa7ed75a84dec6164b743e807c81d8cbc9f65e4412a21532c9454f20ce72236ab2b07119e7c7b8d5491c11c7c1112c4d46de1df6f6b3277e74e636b327ca68df6b71b8b8de10c74f859cff951e4ee08a93cf38fe9b0dbafbf4cc4d48a2bc83078d35402f343f6fe3154b86ce430db2f79a9a62b68b4cac7e68f688dc5fa2b85a19a2a652805eda75b500d2ba8d6902ef12bb7b379d9ffbe5c3c89cc9fdfc17e7d3160712c9b2815be6ea2dc48e1ad4031fe3f25d32ccf2716952493f286d03b97a77f90d53b7b0baeaaa20822a7795f4c43e2f65486bda5f92a83c12b7bb575e9558a34e11ec033f6e275e6d32e36f6f236326e7b7b50b15e67be50eb1f47718f76cd2edaf3877c21e7055f7508c6cbd667e60169832f05419363b73577bfaa16efcec39f8c3e019d41f3b82f802d58fb2540c9995fd5adf08ef815a77c1513eb0d4b9580fa4a8f9b04aeebb34a3db14865b2999b31c313bed841703629e920605fe8baa399b3dacb72487ad04e06109742475abc521efa39494c032fbaf0e77a1b8832efeebc0a9ea9193b17d2a4135c9a3b8eab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf655480604ac3b8745ce678b1644645de2320c4544d4e0c0045f51e70d2022d5f618c38cac424e3be0dca2e91b3375f29cf983888f6832f91b10ee7961d5c24a5e67d6f84b28f0bada25bca88e406b47a3ea850a4a8f7d1b50e4de3cff223d2741b6e963fec9f8953acfba06786b6313eac482f63c8d2eb5df83196783f5761434a528aab06f49b07e2231071f748d603a7209b713a1d8884b70c0cffcbe0f9a71f5b8ec9756fbd8d19317d3a70140bd2998692894c9439d01b2ef2b313c6f55e7b3415dbe6a82176d83aa3d19e462be60d0ab9d899aef265bb6147451cc23d9e3334157e754dabf2d8b4cf84d601d4ec40a0bf18d648d2acb8f01fbe76c6c52a81431eba878fb0357c00bddf2dba512951257737c9108297ff96e08291edda003156883f3366595009906aa1fad92ca205d4bb69555457c9aab62fb9dfc5656d514d6ab1d2a709741f333e843cca15104cac29e2581fc78589bdc4529e0fcf7ea52581a845fd5c4816ede133ce07e9378e341d2c3b76997207689a09a61edec0f2c2490b977f9da57a857e0dad0a9fc0f1d287331090521d00795c87f7d8d188aee06fedeadd47525f85713bf42a99fb6397e22fce36423580073e55179089b30ec5dfb7eed637b7fc3ce8eecae2178eb698d3edecce7aad96fa485532a34bb8c6a764d924aef1f5b9921bf8227ea143951553dabcd29630912e5ae38ec6aaeb5822b9e80f29acff93ece75155f77d82af461b32fcc77dc71a9471ceaa573fe5d5f85e04c08ca6d95f1c3cd94db1d13ffda79295c276622a19701a8ae8d623c020fe6ec559ac7443ee08f88d1ca732ed958fdd8394aec72e4100eb9d4d8651afaa5528c5ab9287de6152e37fa279ffc4a4ae6e2713d0ebd8823c0422b91f4090b3cc76aa48349f606e3d92f51029935703ac113114a26d575f9a7894c210339e1ac4047c9d0914a63854448bef762aee52f5081106e4dd8818a4895d29d5201a9adf1a0a6ce73cdafbb1c97549b2ec7477678bba3089371719971b507daed7b1cab58007a0d4614e98b1b67c25c1d2b13afc309a823824495e8620cf4e2e8dcaa93efc8571fa41216395207374012dab5783bf1ea465cedc4c179995d9834b05f76c4559405f8d8de01e4d2db38db6922a4a644a419f8612afae8cee5eb2a5936c0741fc873d8dcdcf301e6c4d160c285460245d718bda6dfb1e4df370b2766885104b6a7064c9e8cd5790f0d4b86d3b4b62b69265ee329b40ffe7780a54cbb64d2359ce3c66e140e99653cd4e9bf7e09c3e228a93e7889f0d83063bdbeb98787f65f725226e55bba76251800df405334e073936a6b4125e3b00fc004be550a004042090f00a0161936c6c178017a7b74e3b5371b3e0e298ded41f8b190f79d8c0dc04fa12517f1fb71aaa5cfff2e46f067945a43e9f7150f11ef1e918bb6ab26b3c748d9a82116b1e11040051dc9618695d997f624e10e17d481807a017866c374cf2b29c4c43354ce9944ba15eef634c1bc853e2351702fe21700464fc0ef473eec61afe37b7140c47b96774f92013eb7c905552a7b67aae296437c83074b43d11cecc0633964474981c92c3dab1904262de4e841fd6fd6b8086416c57bea0c34b5c4b848cb5ed005f58ef45d73ad3f64cf8e0e75e8dba5c6bd8fd2cac678e1b5390e429e79f0a2ebd105212ba5c180d502e092e27707324328d341f143bbcb9f30b980a26d2deff407043c837af7da0b3e96c33336544429df19b0fca59c8bd2d8a16afc843074671a259f3e02c89f007dc18caeecfb4b692a398570da811f066e7e1a0a9d1d08fc022471e75d089eca1ebf7033b839ee562d0be77fa9637c3629bfafa16ab37fc556749209964d27d7eb8f64ed772d5a9c88d98189f2cedd5ff312cc57f981bf1bd81c313840e73c501af57469c23d5fcd01e6e3dff2cf4f5583f70f3d921ae9e8c920dc195dd2403b07a7cca9f7072493536e5da85457e01885d700521ba00201192c41101c1ef5139585c0c07f3511d35fb348a77827a7a4a106015ae22462281455cb4cb9c72e9c331c806521853a3d2ded8b4c6abf92944953766a88df4a471bf39e514c463efeabeff349d25bd39ad3806b75c3b000145cd17ab5d27a148a27ca202e6966432558e214ce23f202a9dec0e65e97e1d9e84415fe311d44140135363dd0df14e6fc84aa59c57344fb6a8904465af106dbadf48b7dfe2ab5098616f174e77a9684234d0df72af5bf764fceff8f28abcb6bceb18a8df1ba5bf0479894d206a023688f7a8e6c502fdb11fe28422a75eac397df01931886920591c5a437edd23d51df5abfc7fb14df38c5a910777d503383787d532b6084c7d10cface5c3ce81376686483109576a2593444bf4ff59d073ba12e14cf902a7ac063fff936c40898df4659eb486a168053d8d277ddb0aac16636facea28f5931695409c26a9cf906d396887dbddbea1888c024c580d3311b430e46891b9b8840151ef3563fa054267c07e904192886b5536c777d76cdcc9bf5f184559df32629dd6184bbb2827e24befc8ab8b3444460196a5bd3fdca6b1a1588e8f4afea9b0ad898a25b09b6a07ffea4a46e26e572115eefb244b43a828b46aad89e72048f6159b074b08b8db0440fcbcc4f639db0b310b80e5493bcb4100d2dddd6e14a75a384f7aff5113009c8eca88497201bb9adf0d3eec23bc6adb045a76acccafdb669900a7fda7db826d1f82e9919e020d5b05969f20b88cb698186b86190c7e2bab993246e6a633ff9cf6742f7730929641cc5c7fae8f2704694e14f5dbbe72b4270d45aed391f3dd1ed04def1e672c71230b1bfb9250a490d730de13ff2382d99ed3790bb2fc5d207ac441c0eea205d26fcd72a6bd5c572cbb07f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h718135d5823f4b3cb8f6f8e2b8dae431996510c98b0fcb29344fa36eef49b8fdb9647ebe0304e38c0d64dc9ee7ab99fa79b41f6c85af3978fd356b5fb71cf2b1f501c99928304b68dc04f17a0be7849a0f4ba17a60542b2e6c9954bc32f2cafee3741d0b91427d3e6e622bdc826e2dd159e5f078025994586fb83deac065d6fc8d87f8f055b80c00a3fe8f1aad2b066375865c17372e5e2dddc42054aec140e8d3841f9f4e822545c6bc29aeb0e7b62ed7fbafa880cccb566988eac2eb6dc5d276ef515ae878ab425da697959f3900b99e5e9691cf8560f88a8acbd28ebd99d81f19ce848fef02164f35e25a6b363745e479e881872302585467f74666fe675b69a0e129795098fbace7c8532ff975fbbc3d711f861290e61738a2ef6b602c1359f533045f7d066fb1085c9cdfe8a6bc620f0e974ea07d014584000e2fa74070c853f0120f5a4b1fc498465ab0f298ca3a5208f2037b0808ecd7f9258e090dd388882139c95f155a9d689724c95518f32d48161ab62c6d927ed1303e101c9f256f10baedb4bd483cca294a9dfff0d3a586ed5d83494c4a5eec37b5060627b00ce9a3b25e381af362cca5974bbb3b79b20a6808ac06d427abcb087c264b4d775453b29476cf90f1afb4c86d9d0fcd49e09b3108a64ecef7c5af25245c6dc6831451228ff309b07bc1e2ae4353a77ae54dd9c4d1bca4e871068cf164e433375d083e173a363b3adfa3107837f596c349ea6535e0e5d171686459ca4cf2e45d48a027b4a861ee22e280f58d3db77700dedc7d478168b3cf3fbd9494f2ff344f83f728b82adb3726ac57afd78a16d8a6a21c2d89385707eaef41529754744530e67c2c2253d01fa9de454e13988bb353348c8fa6a36360c5bfd4615f233741347cc273f3839e3b50b650b6bd0e237ac52f282a25f96fa0825cc9b798934d37fb796244f70bdd59ba8e258ebaafd1b4f2a16840c1b5d19eaf5d3e1f7a563fa79032a1baa1ef0d892c2dcb3be0adddd5cfdabce6708973a0bb430635893e0ed3a18a3abfe1fa400b61c16d8122de80c44ef9c6d6ef6a603c8ff3f0fe69c6c3653c828f96028e797e47d3b884dec5adadde8f06c7a5d8fd070fab0e3d9992ccd37e362bf216fe223a9859b720c2b71945da9287167b8d0979f016c261dc021bdaf3e6f68e5622e7f6dd149ed66e11aa1ee5ecd0a6dd332fe2ba48c6047e6cac63f55c3924e26f6a6f2075b7db946a775983415aec7aa8fd724fefa67e9b4424524ffbb39469afd050741a501ba10b53bb7180d7afb9feb44661c07f017f29ed9f2bf3e947a1b9ff8ead764ef484f24c0a5aef428d47b7d84ea426104af88e148b2e141198ef64c86591c8790ef63652212efc57c50f094beb92418c32862afc63b0cd846cf93a370f9fec40a20085b3099934c2e145e5171beb96a16b024aaf2bc76f281fd86d88932c797c4aa53978b4aa58e81856817bd08a43e2051438d3a1b2d255af38ffe8c5abfebadad68910d786281831c06c92c27f175c7cc25f97328835fc56d7b0c0f4b31af1a4f3682b2a1482f841da500b8ff58a62ed4e6036366dba2d987f79b852d43bfa7eb44a05a1e9f58b2d7c80726dd8fbabfb4f73a4397a69595612018a3720ea7f287e85d29fcccafe4e075a97056d1e7ecf65f3ccc096dae651a78123a352a1bf11b2fe9468cc382904cafc2c42fbe84debb32d76982de740a0e9c0f0d57dfda7d35cf9036383fd97b6e9829c06d128a165978a9dbc196ef7082634d33892659a8ed6f00f295b6e4e41e2b14c930d497e7e17028dbe47381b6574a3618ef6a2f7faee3ae6a8be314716796861ec9fdd3161df8f54528d42f6a9eb2d1dbfbe31f3d8fd0692efa4704f363a316d067f75eff4c70d98ed6e60cfc2f88b94b66056b687cc041e94e2646403adb821139dce991146578a272c136ee59c88d82dfc9593aaeaf3416d7f7bcc258360eb0457c606f9472bf794b5474a3fe0f998035a74f35d8af831118111a10a41830b9dd88af5698676d5e21205b186b4db5cf47baf963d055227746ad4fea06e71efac9dcd26fd4a7dfc696d146f6fa331da60d4f46b9289363429942188c0073c3ca671b62b5ad77e709ebb7d9cf621ff73dbf3dea65d7c4f19a233f8e120fd0b46a2a0dfbda92bc8a68291b7280062b53c0b3eed49b14761e010f3a3f813fad62af5dc19b301326e7217e0aa64359399bf11d4ac9e78785844794be3714584fc2523eb4d08ec506a093603aa8a66f7481bce46c5d5d5fe8ea3834dd11746198f24b95e65319d0bab4be235f15c938183b6195bc7ee432ec45b00986659d03f2e51c40b65ee869f3c9eb663cb2c91d108b6d2088e30095c8da88570fddc3cdf5579802fed0bf315b5432a078d6948f816d3d60e8a7a00fadc6eda6a74bc2f076da6811b7d063a0104c6b53a871be88cc42d7c33f05564bddcab547a7477691d3887be2fc3ca73a28a61c1553df269091438eab6fb44c4057360e77e5ca2289fe3827706a10aeb6421737d4595d33ae8dc85d13bf24255f5570e8801c36e7f67712a83bccd49f437c060034c1d62ea604fd361c88b510dfff06886054716972adebc0889b6d5f3180dd3f82186596ffa9fe863f6c6b3f440f7db1db53beefb02bd5a32798c5cccad9978033c146446015b30592b5fe4c2d0c1baf59eeb040b3973da522fc75aed9c7a3f79960532a2554ffc0acc358ac0b4fab6c9117f2dcac7728bd44017bbe81491408ee58da1411f1add61be90d4561d274840a7c510f681b3c28699b75a8e7e3b40942cab424c01e83c396d02583f2167ce66b48158d0553f6cadb0e9f4b1fd817eea0a3f60a267b6bf66ce937fe52df6260bfacb489ac055090945567f65332f0960b0f623;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h69e9d8a4a6829d1dcd6306b4834d6de0ae0acfc54b09531d29737e3ee83c6bd10df4a2273acfccf9295bbf248e40f5788765bced7020f87db78d05431d9f3cefc2d187eaae670a5f920fbda3b3ae2b3918874189f69c6b22eef3c94a9e20b234b58f1b06744302baf4495be43de705d4e54abc2eb867dadd8e355502397f76a3ab3def37bd9f0f7b15f95f70ce246cf89902d30d85a79b5c6592b36f3ef0b9fa6a63148f9b43edb6afe5ba4655dbeb6b657780eab92b1012c0456a5af825ef4a75125ed78da699651300ceec4da86c80994812c112e59c9d3be1e5a9c723868a9bae1c368c5b25c19cdf921439c0a9cb208cc616aa0de2b872cc1a48648083a0da90c5dcbb6301e0a4a78a767f96cf1310b1a380986fb9bf4ede42b8c0499fe5874375a99d3703b7767e9f83e374f8313918467944654494dcda94229e48c972b38b33a50dfc6b3a98cfa78df6d6bfd947d36d9e66e8e2c534180a32e4bc003e8ed1c7dac27950c829cc79dfe285260b007cd0057bd4300b38fb82f6e43c2f21907ce023aa1246c6a50c839f32467a5b7794d3383a22053098e10f39b56bd9cca3ce813b02c62f4a1065460e53733a19d70235b96cecccc67934cdca16cd64b06e0e67dd28a9c133c33503217fe29e2ca15309be3bd05a196616c8b813f7fb7dd1611b895e977e29c226092d8532dccd6c3844ec8fdcbebdac6ba23a78c4847f61a364315cb63f0d285b1fe5d44db8e9551c62681902e879d984ecff3fe52048a39f783efdeaf0efbd7312b922515c4271a7d3516e207f43fe3f4c311b7137a328deb1832c8c4e125d30cf5644deddaa7f63e0e8c97b39ea9d5c11832e4329bc115fa0d1cbc1c4813d99a442aef61384959375d2680bfc4f305c9fdb980d2984af38fc9191f756da8b3bb8c2cff451d0a7e581d38cc39da5a331cdf62705546ba6042f0b72d67afcfd2c60cd3dd79c149011070c13b589d13ae4ebf2f3ca4c7b861147503336923ad0b8276bca467c843dafddfdaaf03eddf61124d080b146f67c9d4bbaad31ff591b10f18e1ef41dcaf09e68d2292a5927942bffafbd54f03d715abebda21cbec2b0b2f8bdf82a1647984bd3028bb68cf0e593ab53e3c283c141a114d6519941bc797b0a05eed8bf7fc8984f67fb2f56f44b09efee3e25e9ab89b2bfa4a5b621d1dfb108a21419e48f18db5f80854b0bc01fbef272fad83dddff1972350df6e83713ad28001e48e86172d9c27ce0943562e3f6758abd426fe511bdb932caac63bc0fd7a1f38546fdfd82c2b2474df19714c77af8419b803e79763608d29c3609937239f7a256d6a32cae0849f34d9372429c3c5138d39ce82ff643bb6c55e1ca37cff4296b3b856e535c4dcf7736e04281af05e8ac8944f1853b2bfae2f56b5b78308e3b83b65fc3fb418f2f9b211d8a3ec6d3c2d4bc26ca56b4dafd7c19b746f726ce7c21f7a43235d1b43f4ad78862d695f59a0a53bebcdad4de3d1125d482eda7d3e42f089cb81843efec0571529587c6c3bff3a28d1553bc0c897769d1f5b355d19bccb337aaee5ad04e76d71b68dba58cfe8242b001b0793c8faeb125922296d2b0c264b7a12c8803bb998889f738d9e7ed276926af836bd381e50a335b8e5bf7e13e150a53c3c7b062369fe62d348932957a377092a2415329d78638e47fd219b3ac7a8e8a6ca1b1e77f1a8202606c46a22e7f0b18997add3a100c5b5b2f3c46de11900666e34378457b5ddf4a3cf0c0a54119782cf963b38debd76a562dce2f1bf522474aaa607b4432d31e2ff8375289ff96381709492af445f60970c1e62cd3337f91cfee36044c2f61743bf10aa55dfec33fc04a68e5493cb226798dd7a6e14bdf0fe412ee15871cba579e62f4a41913faae341b73f12c1c1b56112a864fd44a70a1ad37ad345fc479cc0d33b05c4eec26723722c48d47420eb66cbdf609a678c5bf33ae3d7d714bea89f2cd2d5505666d515a4045e95a9316df93da61bad4bcbc1ae0c3354adfd641476d52ed3fee32cc11d2559720b4ffcc1ea0d48429be4606d6a24bb102d161b017e124f7d2027849d1e715ca423140e0e6f4a40d70cece3e09708875446b851483f58513a07e275688fe73495986ca9101ddeadc318b89abaaf72701bea742fc74f7aae1ad93bad07b723a42f971063adc958aa44d30fc3d3724c8146bebdb95ed108d0208a401935149b5d4fef2d48851da500fb8cf4b00b7871cc4bde13d03e8b96f5b71369331f4b8e8be57101163f60429eea4fb472fee631d8542ede4bc7837dc3d8b7f6cc213f4b4b0aafac4d95a1b400a8357e15c0286d7b337483019236b278f38d0853ec91a3bff9fac4e3cb1ee868dff1cae4fe88b152afdd9d64813d739330529b9f37d0f6c300df82c038c0cc7652286fa736978d121a1a10ad70bdb3d9e7efb09b937565118890d58adca1e8d260bc177abacacee1c6de4e2762c72db911d00a27d397196c4099b6da6f5371f1162f1b8fc0ed1a1052aa123bf81f978bc871f956a118011b52d6c5f959ebbe8c17e039b59e1ee783423c19cd4c98221f22d94309b9a2aee968a012d17f6208777a6288678f6a3062714f600bcbad11db5a438cfc3a362a41c4707f7d890615ff25367152b196f6976659f6c6ea3b74774a16ec8476ecad68008b59bb3febed668eadfefc347dfa3eff52e054b5d910609fa0556d9c12bf29c346dcf54d462e6cfd7d0a39b96fe787b06d441e64e00d1c0b95c5d301a7ea38ef6ed7670610831e3c912dc2d06a645c5c0ce38559f2501679b4374e502f81d437d9d33eca14897f16fca281387bfaa651f890f17de4d949c63b77836c5bfeb3ffbf00172fc97347f6f2da55fe569ceae5d727b95df6eac2b17fe7183fc5b82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h945f2f7c100816051b84eb02ae9e2cfb78e2146153119dd4c9621f30971e3f3f74455e648f724470a30ab9bf55bd12233530143324226f8be6151ced6f9828783b0421807e3426ebdaff38018a05cb1da25203e5d337fd723d82caafc02b16f1d51c3e2bd47f77c287664a9f8adaabbd0a41afab1027a84fdc284424841f4176e7c6de6122a40d5cd4e98067182329ab2d4396e9d8ce3a66d898a029045371212bd232683c7c8f3f7896ecd31080c313d13b738faae7783e8c0c3301b8122a0906f2d89bbadf417823306608bde0c2d211c998f9efa21ac2b20de0cccb33aa57d04a20dc4392e93377bfde2d1a9282673b65fe6fa3fa02ee32162464583382892cd58094808ea032236b00c9610e4893822203cd54cf38db2f021c8b61e4b138a7d4bd7689c515938b89f418cc8ef68c7920a15bfd1d92e7bb37aebb82d6138e3f727b63855dd241d2b0baee5963e0647ec48464280a3e1ebe686c5e902d33a97034fc132d77c8b49305c5d215858eb50cfcc1ac550d2a5c589171e5a9572b0414d651e5b29061d8765819b57b79dc32358fbe28831884d19225630c08e10bdd3bcc33874c1543ba000084a64ecfed5cd2c5aa329af54df59952561d84fe2e97f85893b6923ae8d7ad914a513db8d71e063cbd7c44e8b5953e1e934fa01d2bb9ad9cc7d73a9fc667039185cc5a2d2d5970d18ef9d5b77943299a97239840f58009ddd14ddcab702a7c0279fb282fb937600fab3de2ad00f4b4e09e6fea11562536054cd70b72687d1d64e841dbe7fcab86e88690768972c816c1a47435b10da661ffff72c5e6a32d0d7b66f501e6620c86cf8749678d2c02a030c161b7d008d532ff05a2b776b94b5a1a73179af15b5958cd18b4a01b68c5272663902e6381c64071081ac03ca961ecc84d8bea2d82a871f4b394eaac710b926e784b1b6d2d0b85781bc8723f2ebe28d75006357e945276d8d921ede0b08c1c75da2cee58beca653790e8d237f88551c59ac40c9ed1cf52de797b645fc43dd2eb6539fd6feab8b9415a990c3cfa738c250c0f4543e9171f429e2de779da05d2e66d093f8b7f7885473132f7b31e8f8f731cec16d4a2753230f45b37f38cf69c0ef8fd118f6d45b98feaccfc5b184c5cce1cd38a9e562005f183c314a9a134374b1894e7f7c6a8dd24990749b267b56afee11218e07a430eee24cdd509388fce9d8643e16b5cc385e406c062197b6dc66fd98033ffc946c12ed7f0a281776cc2e98f44c84111eeccfd7917d35ab25452d6e9f46b1485ec6e1e9374246f835da719be238af0a4fa6f76e74723ae6ea9527ba312f461c5eff28776e3c262dd8ca48778ad1b9198c23098628bca7b85a00c47bf0f5ab32c9405a34fe1bf0e9bb5dd19376fbd0d74fdc0d2aed08ac83277cd501775d3dca8bad6f492f32121d374b5d0efb173dcbb6a1613c7fa6d478221ee79034cc83ddcd3e815a7e660909b4318ecb2e9251cf96a2236540df0ce1ea3c31b1ca7bff62ed4754c41e835fc330c11919695ba400d238c8d4e23f1bef683c26eb8bafe00774386cba498445af095c80bd9a8c542a33680c5ee75656bf9f7e19361847cebb470dfa59afa6284fbc7df145c70044942f44367324391273442c6ca0e287d7cd9ad8d745752e20ab1901357b02cc3ddcb48153edaa70bc3e8ed1f4df5bac43da445b4c7afda9f858e0ee8ecf4cc9f04bde491ef0fa62ad6f9d462b688d13908a66025c29cdc753a41cdb9f58d8c5dce79c030f96a7c64b7ff6d5faa1701d417c0f241c08aae14a96638841d761711f29fa96a18c261aed97dbd7e33948462a565b4247e9169630daf79ab5b176e9bb6c9833261c256532c6a8c88c6991062320e8b5632859c94a2a526ffb9c87f997fac1e74c7165f544a4bd8dc73b73227e4ec214fcbc688dd84800118290831850fee06a27262d4b49df5d55ffa37cb23aabe5988e109f51bb2f4ddee5107d788f5b1ed4f1dc588df692530ca67097b186aa41131bcb1c2dab2879fd2b96cf69a5df7e9e1b28ec35636828d93d9661f42fc73f6724607b156a34ca30749896e3441a4d4677f722829e13f258b3272d6fda8c8bf8ee1f72eb461449f663fa40279bfd56604a5842dddfae5ca6c5c9e2c0726ed2533163647e7f519c6ba799b771cedf4b83dd28b3ddf2e477b1da426650a85882ad23f609b211f1bc05f729a9cab97ee7b1f792b9e8a2e55629687c86fff1fe2133aaf4043286161e85ebaf1f97773223e273fc11b0def7a61b94d52e70016fe0235e7af63b06f1d22e5b8543e0b5bf9fc383a2c93ae846605638c85fba6ea67de574181ddd3ad80d706188cf09514443498aa16873213a6f0285d3455d63ab1ddcd203e7a9acbaf4dc2aaebecc77e725f6347851ec30b735aa43355a62a788cf076e6753d89c7ed34a777902d2b6f645c34c7eee90a1348a99e9801afdf3ef7c168f2cdd9cfa35e4a0df2ab1cb38b9b48d6431cbc65fe73a75dadd75dc4671551e90026a819e1e265b9defc7fd0b6b93666f55011cdadac0812f091c2c4e22dc79d9851a00006d0d6cbb894d350d3100b5320e7fb613dd7fa91d25713fba22e309fcb2db65da734170e9f29e209dd4a6c556ef56131b1418bdafff3533622b6e5672188c666848b145465fa000f5e22f8db553d22b474f2b3b4ecb1bc45f1619d78c5c5bf3219eab57e66a2ecd588bdb5d310e1d4e9ff058114625429ba6754faa30bd9a9c9b9fdcd5e7b7cf0bca9938540655631c9f52804cf598199ba24be57945b2c7dd048c4d07dd8a5030cf414d0e34bbd3d836e8fc54490c1a52f54771908bd373239ffa7ddaccf8186a1f0e7e7c595b3bcb8548ec3b519cf19191809f47fb1bca0eee04d26b50ab55865d4f4c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h34c6e7e48128678a8f48a47c4754abefdc039b85245ebfd5d01451f05892a484f6427d1ed2e525d682e780145d8715192e6bdfb3e55ad60f132fbda37b1a4adc90e2d9c9e5f9a3c8277cccf841663de3047a529d1f97bff1c12505d5da5d2e02bdb180fe0dc97efad3ec77b5d8224b10f82cd5cde100dcdeddfd38b785e778873aeeb82cb6f33af58e09166c87150f9a43ba1f30ad832b3124562160184e9188bc95716d72ac910088fdbb6986a0846dadd8acabae2365f3b7b75061a51186d19152d20b9298be1e4ec6bfd70a16f5d1deb4d5d1c396e6ede8b7efe2d81fbf7d25e4f562d6c226528c04e1c779a87831bb2ab17e9ddd39c94cd7e720713355ef7c1352a56489f054f788c0a36fc882a3ecb08cb2fbaa550f858122d4ab61fdd3b2ee1663b856662062fa9c515e56416e9a594066cb8d3d3e78e0da2602f6b8447ac97e156281c4ce3c01fcf98cfbee5d8bd00ac2c695ccf07b0d5ae85580add3f59b18a7908057b375be4af48d73841cc49b1ccae1af5f2711e3fd7ee35fed26a9a9453dc1e06a6b05051060b8473e6b622ca81730e9a4c9ddcedbcbaf67111ebbbbecda22c9f7127e237ad515c196fc19c97815c8fd1a833dea0266358c8f44a62b667bba63801472295a5a25c1870384f36c53b6c77dbbad7c2b65abacbf04ff501e705297cdc4ee7eb4a0b90f58c1c4d963d64d39b38d52e0902031ca02d12781c496ea8942ea4751dc9a9006e38994c32ea837049a7b93c041e508d27c6648ced484bb8c5e95389f49c98bd1a2cd763d73c96b1981b9b6a50919e3440a2312fd847b44964ee34ab9962eaa09cd3527a3695f41fb281acfba4bb66b7018b4866f86b6265208bbd7820f1ef38c2901bad5b850457989923f401e571e2691503dc19814d20efeee63987ad9ec0d59160735037f61f5fa4f8d108c4c7eb014629ba61828d4fbd809f388a58b62d8be6f0a8ed9c73b4b57b270cd9e32e0fe2d91d94a8d35af4d8e09227404580461ece84b6f27dd434b7b1a071e93086a998b8e2d93de1269881f2cec3bfcb567fa8846dd6f2c119325905d169da50de317b87de31b726e67f3237ba1d04e85f9c021b2efa9f30f48c0241a4182bb9fcb3ccd16dc5b75ffa9ccc2257aaad7007c47c45fd7d690cab75b90bfe7060240d0542df94b3ac923a546c1976a445a7d8f6651a3f4918a3a40ead0f72d6c698568ec238af3528699dff8d1e7e9fd12343bea377d3b0727683f0d5a6879cc07c539377581a556ae4bdd3b3ee2db0bc0e04af3cb054745ce25cc2e4e5ec728dc3c54e56ca492b72321f244391a847fa388dce1ef161a567b3de68eebb0c1a470b42cfc015c6f493f565fa24ffaae3e76b9ca2a0d75b79cfe27cc92a172747d78657cb434cde942fb185438407e526d1c2175bd66d4a21c5cbd4fd7bc8f5f40aeeaacec31d6c48814f446d0bfa9ba6d5b3cb97ff03705cb6bdee5eecb88f87cc46a4c5a317a923ce8b176ba0886e965fe615e8fd720a4b844e7c2795815039d136ff6714b625897118315b0818c7850d26532ed5350d7a2e824c45cb45f4fb707f2ac48b1ec9e99b8de26b3576400ba9bfcd3d99f1650ae670ccd6d16e454ff30457b494848ab1cab208a95cd085be4256d05ad016b37ea4621d9ad6d79846c4ff4e6e1bed5bbc8f1a983516518b7ac6544b4495ad0a470ea40120ebfa9c4078dba281136cf31573d62af39c2353404bd7114005c801f417751f294a6ee39a6bcb199a3de722486c398e1e01c81534a7e6459d0f2e379835710a0611ac47f1bcd9df6e215445c0030d6a86a788d1b36542ad1da71a8a66f269ad71416856efec9f5af34691c6da46caf1af69d48af50d2729f8e90b5e644f13ffcc46c5068faed8d0185f5128fd617eae4f81ca569d88e92a375afb3d6747c84e080c3b3c3e1a551a0926c2a39128351f6205c69fdd7bd1a1f3322e2bb4a39286ad06b2c742640d48916e2cf585c5d45db73b5813b32fc87362196946880f016cb01006a8140d4a5fed682f61e1b889a3fb779cbe71dcacf6778e5ab33837a1b8bc7a01c8faf3ff16a7e2c392d9f191f2a95da87d1e60c37c7a660b4b4726214e5f694fb899381ca73c059843762b6942f08bfff0864ce5a8ffc2e01d8713957c891e3f5d6e47064df6e69851dbe15f9ce320ac4f376edf3a78d43290260d7322832cb196095f06bdd56b5a5cfacfb104dfe5bb84a4d4c8863034a722027a66ab1e41d4de631e33605d9d2f1f94389ce8bfa9e1c304cc9622fb879658b8a3afe11ec555af1fc315d14209b0ce3b8f74cad2e2d4d0428efea9053555730db6876cf53211cd2b8bdcbd9581163eff0cbb71b65091892ca5e3fc07dacd63f03e2633eed63553cf4032708e5229d759892598115b21ae93254216364763c0583fbdd0c311e23f2754f91510208a316f3461b57b0b4bdba56147bbc9c1c7ff4025f2caece5823b721103d68a6987aa0af83a5393b42ce88dc2499c0f1c48689846769591c47b7919421a8be532b63470f5510e159c6053236a3436742f613b8082fa9ee79ecd35f3a153c6093b1108773782b077f20e190ebb22df2b9e9fcd33f5aa5af2ea3fd337afb9b23d8d4c8ab69c046c037e1cb207959533a514ce6aa1ded2e5902142725e45a92bceff4283b145cfc6d3beba395e3ba268e3d492c52ed9c060c755aabf7c6965393b14bbf02a2d6915ba0ed8211cf08c43a2375307c1144d15953757c80e93f073a08fd8b1735cd9261d36eebb3e2882a93f873cd2b5b17f640612fdec09f8247a45d6e631bfb1144e6a8c330ba0d5f24e25f7d9124cd700928915722ce266dd1fc9190ca059cb521d483e0c6c07f896e54c26f2181bfc467abffe2bd260cc1b2dedad8f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h36242f1ba8d94475e3071fee9e1eab9ae1e14a3eadb5833efec6dfa079da4721239d9ef9a50950846cad407b87f028abfeebd348b0598455832e3734ee061f0aa677e07aa01c22b9278c7c1e4b99b662e39fc81c2f817e198052864395b81fc5be22df97fc29e1981a7dac85ff3fd4eb8b310c52ba81e7b63f8329997b22b31b8e49fce2d922e98591f418a6e31dd6d65b73cfb5974fd507aa202d9d28b57c439cc971e7c307640c14a81ee90b9636164f027ba9cfdb9a949d6b5ce7a105a765ff63bde3991d15af91304d09d469d7ae9ff67fc7676f0a5d208a6ab4eb51f57fd9e50e407750473fb8eae868192a4d7c4bbee108f0e9e82c4e1d350c3b48e8a873b8f8d4b198343c63ff62e0fc6505bd20024e9d03fab1f34cc28449d76dfe0eef4a8eaf025576197dcf34336f0dc27cdc21bbc77172c05580aaae6f9ef216d9538656c98f7b135142465b740f675b900300dd8733dde71c9739c9ffe7203e8d39f91e30c3f0cfa72b6c116a58b6e446c927ce02766db99d5bf7c405172d44f229467368399f771351952fad65f2ef887564d44c652d661ad0bdaf45072f963e33cfc027eff03c3f4fa0d38f0758c241f49657808e3b814d7bf3aa874939a48ea8c5568bbf47109f04bd7c3212a65d71bba2547d50159eeffde3524397f400985ae30b2b051ae216b16eec5edd1c9756f60359e6649f0b13b04d5540c5a01b71a4003be1c80700eb391702fc43607c54bdc63cac198ab1871401c35285e4cb37d87ce380869e1266548320ecc6b8eeaf3c9cbacf3e983013ff37075a75bf2c717066012d6c58c0908a91f9e9dbf399d9f1fe456ba84fbd2b33192e14c9d27e87b0aab59303f5426daa1106fad75bde85722d46e7ca7d020f71129420356bee1ec69afc1547ec8aaf26233a1faedcb6a7b0d466ee5c3d6b021888243f78ffec1669730e5c3710d0dfb509259121bf2afe5ee574fdc568476bfa90e7641f0d5a21f0fcccf248a743e5eb44a48e8562d34a3b4df92d6df12dfbcf5e4523be16f5a24a79ca759a06dfdaaf1b2f34118d2fe226a14282e87e3b3d79d38e016077b398749c039f69c8d5ac839ffee89bd3a093135d452e1a15640845f1e7107d9fabe1bcb4b9391d1ec25ad534ef364146d6fbd9d6f9258cb6c3223ca95fc4186ed5b6366841de3a0086a1accfaca832365143c99a9998afee910b235b774b0ec21ece16be1fe6f5d389ce4dd9fb12c805561897e09bc52dcf50eb7c9503e0b3ce7e7938dff427026bb2cc4b654db0d8565709cdf1e0a5a53b2090312ba3582a4e3af498bca0cca8e3c017daf6122699f869b44e9e795679343ccfd219a92144bc02cb5ba1f023fb6ab8559ad2c29ec81b9dadfd1b3a6933a417661458d8ff68445dcdfd9d9c139612b75602f1c80319c7a1a4bd96da5e1758141ef3acf274c10011e02a5d2fdd2c595e8522d9151a72b8a8cf6bf4e0c99793e85d2bb5ba9fd6a0dbc86c1655ca750ca7cd1bcbf5ae5315bf75d320ac786f2ebadeeb66677df634751b37fa03a4f79f4121b1358b463c35117c0e8a6f660d662de724c5b7f34be8835632fb5e3b48f3083a2840ed6b8dd8d982707b3292d9042a7a222f0daf9840e1037e1e59f44b7ed5af4d7701975ce61243671662c8c636baa8cb9fae2ef91b6ff90e5bed2aee2ba2b97af5c5c5300ce1d9d431c31495f3b907708896ba8de800a82313f01153d74795f4e2265e7e0f703750fb1da47769db6bb775e917394329665ed056775761d192a497e8bc9768e8e23fef0e45626e6f578c2fb0cbd4b8c53023bd10ce4ce1fe9f04ad33afdef8c64e4211c94f240cd334dd05511f5a6fc6f89ad5a910839825838654120fb11ce47cb3a07bb35a256fc161888cb92da510607a25e149e345857730cf58e68acbea1a8077d3b51a64a8c20888b62c4cd79a3103fa2a889ad90c3e436c7e54da302064925f3e497613ea0e7ac929ef0b6e777fce9cc404be5bd5585b94a47c4ee734767cbcc57dc0828fdbc7f8a0b26491bcabb2ef0c285c501defef408d35ba89c049cefe6d8e330ddce214b8ac976c4bd36ed7af2e0af66d3391e3b282cfa1a82543f105f3f1663f70e0d83b3e2cad267407bb424edc97c84e3fd466c91ab62c2101cacead5c8ee7b1110b86ab2678347f34e2e2e8a93beb35738a257548cdfbc240abb9374547061d4cc08b020bff4dfa393a3985b65dd22a8f1a6e335fb4e243be13f47c5068f4541bfc4c82e6e56e6376b30122481791593ea9417de416d0ee0d6667c798c783b68cd5acaca63b8a85d6682fac8ce8553dcc5a09f0e5593ce013124f473e6206d257ad0cd324869392504232dacf3a417f02fc0554d8b7c6349d5535817fa0e1036c908edf300e73065d333722806efe809a8bafeb88ca641ca837a6e530bc7649330a0d1f5c910b2680009c42ea07617cc7c9634d9be89e7ec77f516bc24e252730ca61969449f089313ee6e2267861530c80487ccc93ae924e297d8bcde6f54ef32bf97e5d03947ec205ed54c8a663adc3a0ac2b51cee92bfa0b52e3b2105b64b0b9d9cc2eb3048c6af4777bbd43882a7589cffe5462dbc988697bd3f625c80e2300d8274c2e8499a71964ffcc6248f248c8f87d16729a548ac1b6236e9aa2b3ab5a1f0dc24dfd8afcb20c6acb43f060c72a2329c811bf1568e51450bfd7c4aa895fcd02b5762051375f5c902c2d916246f4f511e254d36fba129763e5bc9aa7b6b68a795250cce3a0b65a68881516d2b3b21720efe99119b51e6e17e6b2d1d34e373b0469e5ef22637930116fc5934eecba68daa41c22abb5d7f7739452884a2bc731b6506d5783cf99c28d2b14bdb8b893c365df2d5d693cebcc5d8d3a5f4418b5dce220e88c4a2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd0a68a647b21fba798911b7a6feeddbebe196cdccdbbc9b08130e03ccfb31eea769a50d6268b27c11c62c2e5e0d25d626bf9db169d8165d1a73cdb28cb2451058db212a8b29452b87ac7a5e6cd3cf9010fd34abaaf66d83e5830408af61c5b8e89ee3023f8778d67a29431f731c0a76002f62ace192cca093806d410b395baf5182b106129887e3a382b72d5736bd73eef7820cf3f4e1f3f1d22f84bf0f63607f45e33bc4ba7c40f74a18b05c94641e3d705426c3136f09c9a696d6d4810cae3d2243acbccfea1c999709987c303d03a25f335a692a5fdbeec96cea177759e63e6efc8576d02401abb108179490b0f8b238d0dd3305dbd8aa14940bb46ebd3e03851204abda7dfd39c54fbb19cfea787ff23731e713d27302aee584091335df7e6ca956e0b344e5b2bcbb4e2dd93cb31283e3bea6f122b035f47fabae0040043e89166ee3b4908e2dca07b69a5e0d8d80b72d223ffc47651e73cfcf7d20a0c7c588419d31b3f924de3e63531682ea299c2ab5144e76140b089a29b797129718ba98d900f7d5202bf3fea818f4f9943a1720d8c1620d64ade79d8eb55c258dfc1ffe68f9f0411e720b19ecc35bbb4fe425176f5e960b255b426b85adec93d45a0315ca3575397228b83f68a7ead65f6f8d1bbf5ebe7846f117b9365a20c4f8acbfb39615ab07039fe8451ec89e91d8e7e4268bcec62417ad73720839e4fda88697cdf68c4eb5c6781a8acfa04563d8b342f652d815a0b8b7c4c7a78be4b1134612bf8f49ebb3437c69088a5f7e92898bfca98f80a7b8f088fd42f50805ae9796da6c65cc44e03d187f4cc6494dbe5fe5745e3bcf483e94f434ad67a84188837fabb0a8d4ff1541f2850a673561d3137ccfce9699dd4e8af705a0549a1ce137543d6c107bec31608b2ec15310ae998e2257664861bf1b63cf50e54fae4c1c541666a1accafd7366937288c485df65b76d9c4dfa583e1df177b72e91e690bf3742168773b4f038cec382f55ce5796b38353a44471ef4ab1323c582b856779e5f2d4c88d2abdbc16423e17f02cad10ac2bafcade73b56ccbc34320eeca46fd0f25a70a3ff69e3bb598441dbada10914a7a20cd76e8e73cd8ec63569cd52584aa2799d8e46820e59d012fe10009580629949746d26add66416ac719aa66bd37eb3a3e457a610d26d9ad0f50f4caa069549e107f27423d53a35d4f1ebd79a32438c9fd8d6ddf09a54eaa9a601becfb2281680a2dc42e8fe21cd83000afc8d9075b35233af162f3f41a9383526726e37aa34618753ac608ad0a5188038608838340b844ad4e8961efc116c3b8ebfec99e3a65ea9e60620994fd2acb56eb554470ef9c9144a4f299cae46bedbceec8ed4d453fb59e5268c574e7b75e87589f24bc613903ac621af094e9fa5b4c5077af599af3977bfec9220660e28c4327f27921911cb80b52c1566ec7361dab693b1905c05bd9799ab731b69f12e20a93104a9013a3f3939b5f910f4285592aea525583395ec576b0f1f362ed5b435b98e01cb8d5076ec5e2998906f32b34e21a5c295b9990df4e6df486a7746956dedacfe68a07c250b3e5ff66ef8affcb00601ce0d92926a1dfd5bdfb63bee81b22e51f3d9af0666cbd260bdc51b5496fa853ff16aa13183adc4311db8eac436028938633ad61c82805e792c6c305e445573d23bed0c09e96c4d43970d4ad7f8ee17ecc675bd84ca3e76109d644d2c4039f6c82c18acd8b0327f19b4e33d863eb53dc22715b5e08efacdc9864aa39c6439331ac34c1d208f946b6aba5bc996ce468937031b7571dc6d50a07ffcbf7b8449504cc0ec227ce5bf963d66cabc593a6d5ab097dfa39fc5f562608056fc2c6ac6bae418d90fc6ed73db7ba76b353f1e28a8904d0b6a9212c602b16974de0e71fd2eb5fd0aba2cf831e98380d512f47c0c422f54b279ccadf1badf0dc9ee0341b622d603c74d504e1328e38b25147827d4918afe15f60786a2e40ebfbe8464836d0a74b3e580f33aaccaccbc68424128392d62dc053639d5cb853f9b629b15fd29b3f99249fc6ef25f13b73ab096b0f35006a0a4fdbbf15dc2a764f124a9fb438fc7d282ce0d0fa87ea2455172d3d4584c522c2a64c2b8c190612d904751b056d09404c5d69bc7d5b77a184ec51c990e3feec73fcac260449057422cfa08b175aaaa68ced2946aac4be6316242f2e126996b4720d7811e38a21babb8e0abafcbdb41eb38644b5fdacd5d348581fd738c0c5e9f6b6719b87af8cab99157ef87e62e42f6d0b18e9ecfaadc8c0e035010272e62775870c07e21aa2998342d02bfba1fc4dff6c8e5f3064e166b07df4cd1b7546479e4c1892f69a918bfe7ed7c20881139f39b7626d8dc61935f58d333bedd32ba67062cac4bd386d7022d32488fca4579d2905db1eba3bff6e0cc1888fb653de76856cb205f3644bc34b3ba4a0a4a0327d71bd446a0de097f8fcc887385b037477264b1adf364888d36f6b2f781cbee651b9bcf5ba6793c79962decf7a49b175c3d36186927917a9fc82159eac657d67c414e9d17106be85d262350d7fbec51dc53ddb087fb33a0672624bbb3db779239b26d6e063c1adbd0187f16ad1c2fce7fb1b9720a57b3f1e4aee5b2aa427f11eb9c908cadd3fe9f4f237baf0f0e8fb783c2b452b9418b889e29f711de7156b1479c5714c20ee0f9be06a9ea25c0dec7fdce3bb72c85c14e1e9e1921a41323111a005ad859f2f305655c107408b011869bcc74345b9cde802595107921fbdb116c74f31c4d3139b589d3bc04045acb1bae63414ecf65cea6e817e9d513cf482bf3ee7c08a755a06f8729d01d3cf1c146ace410e604f04ae52e3346503f3ebf042b82230e6a78e2ba864744505cd415ed12e669df35bdd3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h17fa39c6d053477140e872bbb6dfa791467396b90e6a68bb3e8db4db49b007f2cca802181352c94b59b20f4533d1a0fe32a15a73cb6c8d99ea2ca1a9d86b5f279791cb507a1487f40e17fbf6895af17a6322d1f2a17f6db73279764b0c51ec7e4e53095c4c124f2da0038d60cbd55d5bc42eb4d7022f63d3ff8cd7e9b32172b1572f2675481f305ee3f15bfb819928e688a2f9152082fa39d3bd43dafd32fecc6c7b96356e731b6aa7fb9fb570f879320c54cf03b3844f7096e68a7560101dff40ca8e36bc4688da8b8cd07b7367396381e253aaa0a804c6d0141dd0885f9fe476bf0eda43c8102e0f5f4558f6a1668e7ad9e0f5ee1d9511f2c455437fd77af6c865cdc94864030e573a39811da039fc0130b23edaa94f26d570d5b80a550e8e92e279ea709ecc29ac41e163cc6f159067558583000e5f38c807cd91ae625aa097543dfd29daf7631d3bd5a8153988abea6d2f104351d2f35a4a6e12646c6a85cb2fa50b550b663b966616f22e94cce739e7f095f4b5ab04819918c4e306139e912437ca5502f6b084dbc05178223aed8ffa667957c63895ab6fda65b3816531cac723d69cbe0d3c4425c630424c3fa02287acd73a17eac30bb478b85e3c1a7be490f96851edf10038117ee5139727a23b946a4f3ce840438f7466acfeb98619ec0ae23c7bb584567e99e4b63161004738c3235e6db5568ff26af3e8184241d10d66323c185e72eabcd34d312eb22f503c38eb192d9b856820eb9be93afded6df6d7e302177e9e8e4afe554a35fb2cbe5df094e52c2c06d431181fd22c897ba392d3225ca0a7d69429738108c0addb8fd9f56b8a084ed8101683539ab4f09bf1d2317c089c30502f5e3cf7eb37893bb9e0733359bae43b1f99b786a78985659f5c46a668200f8dc3f96321ba493ef6ead5e9657aa5219391c527f43678605a07e523a87ee49167fa6c197ba734830713e1e960772de7f8ed5bc0862077e288716b3e467dc57e0cd96cb4aae1d59632f734001a40e49675c74c8ca5be6af31a4d625c57940cdc38f327acefc3a2fbe564296d3a8c04c1492d2ba92245d474789b717f9fc7137f8a832e8c0676aa3ef5bf076a3f28b193269caa580b516fcd9604a3738cf59154890befa3a8dbb6ed037a006288ac4a26226a6d412186ff904120c63d7dc43034331ae63416e6b6df946eb1394be96d597aaa61a5627067e091ca9b2c6c29803731235b12b7ad5fb818f7878eb49a11d14a77172a4613800c43419cf345c002526a9b627b7b2cf8b277ac96bcb4fda6645c98dfd53f640b4ad076accae68334c117cacbc1e55ff8253651467cb9a5c709e221c799ef9d029ef5f28d49bf051c77d784e902d39efdf95628bb36bfb3fb13f4c712abacad1f825a4465b84a52c9501ae4598b4a772b539885b7b3ebd7b2c5eee1751d1eac746f8d6de4be164d9ec383ec8067ec5657c0d44bd414f577d317103888ee3f3104b7bf03a4a4c3aee7402c6ac6f00ba0bf016ffaeb9483b605ffa7b2b84727e36a554db519b308f40074d80b52064cdfa345840cd7b620850532be1ad433314d76bbcabbc90e424ef7e3ec25d8af7add292ccc8f8a67ff0e176dd54956d45c6eb4c2efccc56c9ee3153e8be7b4b39ea983ea9fcae6bf53df2a5237bbe7a7b09923d238c78035973ee2aa1cf80fae6ef16bd9221b53773bc55f787462aba2563e252c20bc32632561302f46d3ef3e4fc68d8e673549ee5b1c7917c7a21ce349c9a2d8db4b4622e01635a0a1fcda2d41ffd9be342745b26d8c818dcd0da7cfb7dc206baa7aea03d62e3ce5a726f06bdb2edd0c016b2a46038360a2f5a6dedd1807b697022c7a5d4091fa5b1dd2c73c4044e61d43afc4fe679584e51ca940f4fbe39717668d1ea0ae72392b1b60606f68742a011235e87a8d161bb524a2088ea22fbef41be3461fdea6728db0b868d6ae67599406a3819d06df4d4d6093c548125d02fd0c21ba315b5c35f171cfc69459d7fdfe93e5a0f1b4144912b8d023d755a3d78ad79ef395c8d07edb0ac4eceae1524eb27babdc120398bd7f085e2a3269f518336e41267d2af8c8e5ca4afb13af8644531fed57cd81695c1a9d1326e2c883debe67305a94e9b24bb165bdcb2c6ae4b016013f6cf4f225e63619924b37b2db6bf5240fa73aa3ad3488ee0746d78bb78a510159f5a48d8d1e1c505dbc6aabb2a91d41d0714e9c9f0e34503c053db09c8df8da60e20e8275bb29372d6c798e30d5708a641e1364a565494d057d271af3d97d802f562a3c64e98a9ca4b58111bafc4e571bd4fd184b99dac607afdd0ba3b1ea80b2c4cf7206b905993ffae7ed68f9787cb85965f7de6f47d355808e14fef3eb1c37cf0b70bdb8e26f232eb2d3c7ce27ce3fe0745f743ff4cbe360b9125e43e48e132d75a51f8eb99df4df7d2b71d1e444b1606435fcff2f8d50712366a4a9fbf67f364b8e4c911c1f3296a2556d0ed86176c88c983614a3862bb8e2da283a26ffa07137f84b07bacf4144e6258ef21d0884be12a9badf9a1f3bbe52efcd9ffbcabbce7dfe537c5e2be2da2b3cf99f1b5ba1baca848f146c8fd6c32d0b6a68ac5032913b1328e5eded46ada2b768c582fd88afcbd4b2ebd50f8f0403e30a6819440bf03e6286794abf79801b59836fa250ddabbc3a784d710b249d77d6f52adbf539ffe567c2756ac21ee679b9d9b779b999d936703e5ea43fb93696b7ed438bdaa3265f85db5b3a6ccf6e4a0ca61b7621f64db48f4056935ae167ccc5311d6b38e3e2a3865b867b57c2035ee43851a07e344e3ccbd81a2b57b37c225b691619c9b4cc7279e37bc033e72919b06e8744769be0830735db2a161c57dea6b319e3e0ece5a877f084759952f397a1e83e7d4841;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h557157a1efd6e08206edcd242e468f9915222484f47a2b50b795042bb1ba77559308dfa8902008a4d141d5a7a566fc3ecd7da1dac374f851b2382236915e736dbdfa8581fb2fcdfd00f1c01db3b835a3186bf39148ebed1cacc2eee82cfe8c6cf3093f20603427be1ccaf41c5a5d943d0acfbd9a6df6f735f49e13122f1efe4541260883b8b203a570a236cabbaee72cf93467e620dad323f4b6e6c7363152261b2a8f74df2c8e5ad6fff4764e3b240be976e7a7085addba49c069477b5127776450e76b498508f22d1f77c14d68dd80cd73d91bb7ffe640d906d781c3085a2a01bf2caa1dcbfb41c873af768c05e52d7607d68e60b5852b2821cbbda61b3ef09777ad7fe8936585ffcc3ac52795ffaa75059bdb34a40ced766cde351279870e796eb36fd512b77495606d40cab1a9694f15779fe34bef6440cb830f36aef4dc4fe00ec5045de6e690b13ae5789cdff7a659b711b08e2b67bad524f0926b53ceeced7ecfa3e817baaf172d54aa3addbe18004aada8ffbc864072acebea48aeac0c915112176cf8fa2ea647c5aece68bcd6a23ad156f202799159ba2961ac69c98a66ac4cde227b9c3ec8d225c5729dccb179cdf693477757ec429297ec3354c9c774bcfaf7c72169414a73746768898e4d041cb7f06787af4ad5d2497fae167f86ec5b0304c328497f7c5108c8b86b795091b533755def34cdb30b117abbb24d5832af0982fceb7d8d1e8fb871e88220e78dd0d7e4c33aa3fd47443f498d467ffa1e044350563c83041daaa6427eb03201964898796bc037a65e45054964ed031e74d9ce6579f941b609110461f84aff525378030b725b30ee81fb0e63200e4cd7c23b3e258db9b7e18b616b9df84450d042b489e1e6cb7dadc6d29ac86a39199f8236219bc42faf0f03d68d744c5d40eedd5b4036b119e6567ac675e6b8b870e1fe4bb29c02db3d4ed104052ed9a0d09883600ec76169d4c1286e69e56fbc15431441f7b8f6690c5b1e5f83cb59d6defd3dc85ba6d009d3f29330f21f238af2f61b92646bc04eaa0480ce06d4d4b09bd4347e4081e86a51ac48bcd1d38d1985b75a1498fec82a5d30615a54241ce732e9c49b0ac911b76017be739f68a63fc75f0f69419fbe95f81b513333b0d2481ed796d152e357014d6b7bbe424e39fb0f0b978dc4ef595fb9af473c2dd7021079ce1293f56fa4d9ef611f7154d15c21c87ee62b1b174ca06eb106f223b63adc452c5204474d72d3824fe20cb392f6fbc6534cb9c4dd9677452998653900a44abe7af7be30ad9496dca4d423400d1282b8a2ff0bdb1aa0e0fafb57eb5bfdbe9afd6ca473d76d240ee8b565eceab390d2a03704b3cb5c9ad6a90dee8a302f319a0a7521489737d3ac2791b5cf574a837769f0903935142442534647850cf327774bc80e88d931761de8d5c35b7bae923f7e91bb28c643fdee0fbef85c5a5508b40be2c6ad38f273ad0adaf5d82d9222ed89ec877ce6a63b015f086bc53887bf0fcc78ca38ccbacc6a3846f4a0209351901cee559e9dfaf56421c3526a2402cccb609fb53648b18874189c608e6b22a7c0d65ef9a713497d8ed63b09784f615e7ea462bee353980f3e72b222704b4c336013bb2a1a15624981288965a9e5368bf9688e75a3f14eb51442174e59960bd978c397049605c264a8972ed096d54525e2731650ced57c93c534927306f204f31e72b467bd8b6d8fd0bc4c56be65fcc06ad3e0934ddf0c92b821688409dfb7af358fafb0da798209dc77521cdaaf6137c9d37e41bbeb251ef582d1ffc060f7b20151f5ab2cf3ff4b3f36debba32105d92ee2ab8fd9a056facf379e8b1ee686ea41b66e1384eda5bc4d03e02d8457a3ba3f7738b40aa0bb34eeaba1a845ed45df0d62d885066bfda6755b9b0e1b8ee15dc0dc80915d9d5a9ef9ff501d45dd06ddd3182994f513aaeff66e079452b16f28e17a97e74cd25e8f73ec2631346f7abfc8e6fcde883171e37c98b76f30092798631e4e8902c32e5a89cb51d0b36bf1c3d42b3b60ec600a316cdd65e688a478b0d12b3a3461c987dceec8957f68e3fed4fc02707e3f1ad6f443bb25a5d652189a0140bc3ccfe25a03b07ec3a3700e211c667e2b51aa6c99ff9a681a0e9f39e277785650a2a722811dd884cd24363aab35b25a2f3a54577c7ace9cb68b31ce95c81983356932dd15647358f00915daa09ea436a014ff61d529b415ff51616879e80a9e2b6dad65c840e9ae1622c6093e3bd25b2269d7bdb4ccd81b3d9d46e0d30815ddfb1a25896821bdd99454ae4999e549ef1a8b355d69c56a56c8461d3557f9f7ed20fd68bc1179a968654d9a54d0a2d821f627f2943a754ad2c714407da3641a7ca4a6a0b409f69c8db5ad5232bc4c4165120bb60de515c70f8261650c4cc8d688415053b46f1ae627b11d3b270f9d01ea450839fe4c08b1eec513a3bbf51c81f8d15b4c40d48dfd08a8902b1ba60de2218f2af2d842f239a60dce01abc5292b794f32b4bc0c7b73ff8301c4e0e3bc4fb91ff1a77f7f750343862dd1717ae66688aa859b25d09e7b153bf1867e0801237a552cfca153ded04fbe06dbd3ac1159662f0837766cfa4160cd86643eb3bcdff12408f009d1089fe4e0160fa1aef9e5f36204af888e4db179aebf08f07ca2b707fa6d38cc55ef3855759508e6cda4cd53ac5400715e3781038a116a7674c1d2decbec368ddce0b334cfbdd4f50bb196f15f6f6c4ddc97acb2c9838699f1a731c198f42c97f74f3d8efd98962d9a126d1e0f9906b8d946eb386cfc2fbd4e1730ac719ed7b81fb886ffd008604c442b618973ee30d7dd3d104e1e3e01c7ea34e6a96f1656508d3c3e07fd527d0f0154daac0b1bbb0d493f15a4c57832355764620c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3bc16ab32d3ee61648142c5d1a4061c528ef959380cfd8cb1cac23c33ef76f5dc50f777f8fd8630f2a1224466a0457100bc643a18b851634403e1f3d76bab9c86be3a65e30ea2901d7b713b31a0d2fced998e037944078f077089af1dcfa5bf46c7403c0833f8962a52f167be7441b45b17bbb3f4717023d1128a99cdd4264f9b9ed3248500f112825df20d05f14061f1ff13b714a33f54eb3bb3010aae3dfafc3acbef7fd519752e16b9ff93441bd5e66422ca23c358264fbf502d819b9c98cbd923c801afee73f16c5cef97e32b4b427367690ee98fe0e471e25ff817c05a661a79f346abe2205a97e283e7e34b0717cfd038f4b6373f43bc34e8c7849c1c20965f41b837e7f35d92aa96e7ba1d63d3bbf0500f04fea0768cf76dc74ec6272f6c6220c7d701022b81103868e400743435083a38915697014521efbaafe8566dd6395f1ece9650d219c074846d040ef3978f8b3bd3b4dd646b295c0dca2db14acd2daa87fbe482e1d5b6348651bf1fec56cf9516e0a0d0c26f0caefe30d75b35578843adb6b18c64c1e65ab8eb5986f9d16a4ff4f58349560551bf0fab4afdddbac690377c7c9ecee18912db8511504d979fb4c4c6abda9588b10f3cd20892890193b13f8c10870652450b228286254d946365d96fc7c9fa22426d76e881b0def3405a4675d5e7cba2285b406e8ddeb9b53ca9d22c165a0f70bfe7d9cd9ff79340249c7712dc3159bc62c82d15f56e95bfe84164b2307dce9fe234228cc89e2bf444b244d98a8fe155ee9751b8f20415a31d4b405a6421875f1fe7f67fcdd59e9fce9f8d15562b9f076df1a4c454dd66eae395b2f793ede882fe42234731466c22e155d6477854f1a1521d55e3cc7f732a04c6c5aaddfd7e65a78fbcca42efab665031aeeb474117edc915938d8c2f261a3b6c4066ffe01a43ff656e0d78aaa479534be919341f1296510ffad10310b7b05636a8762c17b97a00ea1319afed74f685198e73630c5b105ce33268dca9c4a71eca0cb46eb332bcb0b2f6698d880c6fe5dee44b14f4d34fc38a32be128ff06159653802436ca00968e8e4ec0ca52026384afd2c9a103c78749cdc21a9afbf923e132108dd20e1bc0e84a8c36f8079acf31c5bf1605780008486200eee30587cf9916294b8b7e118f19d37d4e5ad3849586106f646d05f7e837b177280e3669e761f403b5f662690c26d68f2b1bde4de7838a2071a843d1d4636774b78115563f613d5f84f8a8ec488be865525e2d0647f993d8e94dbeb9efaf05642b684a440bcfb02742cd921e821ff0da04047313c1746b46594f0592842153f868a55804b0201f4addf860266479bda80759fa149e6899389461154b7c77480fad1e3326ea3779d0152f995fa6fe8cb64f653436d20bf9c466daf9f2e840307304e02bf1e43ada089b11743b07c8d731e8d3c2503e8ba8a2c36911d5cb65e4ccbbe89d91cb0a749c148002e4c5fd24d986b52fd0602f93816d8f2ead6e5ef30d3a91cce0676f147cee5b360f058baca605d07761073876eacf97d3bc640d305eab207b338e5d6b63a48b014c9fe930a581189299f2f73d999a6aacd56c8a078bdd41d6da28ee0617afba65ea92c606872e2faa6964f746e45bd3fd5de265aefeb3ce3ff5bf24eb0ff4f8c0025e879a1234af89204cf94a2964d83c71dd4acd3ed756ea6c984b0c32ce8e40486bdd2d88f44a10c126502bc74b7edb54d762709d904ba5dff373b18afa60b66c4acc3790c6bdb3b11a1484462cb99ada03512e3699db020383e91fbe3ed4505fae56d1d632ebfc872cd89900e6bcf1458f71966d507d7ecdf23c29af67f2a57c502f21a0085d46dd7d4e80f97f848b9c17d6f653ed9b5ac39b7ebd589b8e5ce36dc91c239f670d76af9b3dcfeb930bb05cc398b3ad99d2a4c3d9444e62bc61d1737412f9cd7c10ae468773ad4921437dd3d80edfdee4ade2d697a9e0438ed759c4ad89943942009b55a8c50436cb4d5f6b8d05a17b15c90549656775b99dd1dcc374895c6464dc987d5f21fa1bd894ab76f86c347705bccd696a66319553c6ebc96b7d8700f9bf1cd781058228aa64e6756de871488d59a17f9517e81177578722693e07fb63fcdc5af7bbe55b20b2a9979e544fc5302618cc9ea185a7f41aa218ad9fecf205a0d5a843c71dc268e27d25f5560385e6a5a00c8ddbcf49faf1aa12bb47e53353d1bb57e066dec4297a5eda40ddc24ce8f8592faa21b787331848acc660ebb0fd411ea61dfa43703b6bf5037f89231ca16d46751193fb75d3004d68a571514b97f9ab54ec9bcc473eb3ffa324f93f45a9abf2c527c3f2f0f48b19b069ec96d051db9cca84ec1c0b49001fa8e249260cd04a6e7b50085c6083fd239dc7fcaba6ff2b2c0a7a570c750b9aa5cccebbaa679cd9d4d55ff37fcd6a197a62cbd5416c12e3c38ae9c83bd3fdb951cdeb98628f6059b4859daa7a91d86380348a83177bb5d4d2f9e5b2f7bc5d52b4c4782119b68e75160a41924a6ff27d3270bb92df995d33b9f58eb8a0339bf027b93724c7776b95d6063006d7e53c2230b981be2c1fba534abe2a680e633c1dfc6afb0def3c4270adf140314aaee02bf3805c883a675300f047879ef8c247086b1e3f92cc7b4dd827f468e07665b744e5fcacd7293c1bac01ff129f2865c6c578d722fc214f3851c0fece7b72543d43611a67c4110dca0705a0147968916fd92ffe0b5113b185dc166bbd69966d05cfd20f00fa347fa0443890f3107ec2b2931bc5be09c5cf66420eedb79231d2858065ada56b98b6517defba1a0fc8b4a3451c4ec70d14568e12158db4c1b7d8b11ad45e0a8798df35c0ec6eaacb3f402bc4243b23bcd1c805dfcd6b1dd8fc5fb2f9f2a33fafc938bdd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h713946869075b405f8d80b008f91602fa9dc85ff04b211c64da83a5e6c818511d9931cbb59b1fa82b6b24558cd6d09408acd70c801d2cf88ed548cba00fb865d5da579de26ad77a4f34112f361763339adf3d93672d4d9da08168ba7b7ba79bc8c43a96456c3e39cff9af3699d27541a49bd183b33231ef6d925f0c9b2a46c78e617338ade8a9f005ddd37116f45b0f25415ddaa8fb22b9cbf4afe43670c95b7c1f90c7153ae2a50d3af7ed75092e3ddf330364901c81f0ab1f46c9dd5220079e76a49c2e1ac334bee32a52d20a95e4724b606c9b756b257a1a1c0e57b420ce0746b816d60f9881f5805589112bee33b014350442f9941ad7d31564c10e541560dae601ad11fcf0b81a9733d065d5e9c996e0f4b19193266d008ba98fd7a8b6fedd6db43df504e1f4f89aeba0b0a7f854bf753c638ea0f87d7b6111613c05dcdd71e27a729b92aa18a2a5ff4028c83fbade060bc94625119832106a445e416bfe88a0646b215f086316a4e5bcbe0d49f34734b61bb913530722a2e7256d23e7cade6b44767b86a9a477feee477e8a6398436c449ebd81b03903b9bee535d139b71654ed93013b5a9b5a6d6e20f82f104187ae6c822596a0611329bfb992d529a0f73d3811c2a113a1335136c91d15091f6348717ef524b18ca32883d2308f3f6acab4cffb9429b3cdc3c725d19f7094457e2d26b5714c464e7e9c0857d0c362f8051d66a7918bd7b82e2456cc4a72fc26e65d7abcbb1b7c5fa0f61c87c43cbc0381ef2a24d7800b7ac74bcab56721113661218d5aecb8c3feac7fbe4d8a92213b260ac2462e258b39c8274177965fb62d721cd18f5a172624997c892b469a7f50fbd4951bcc5c7727e2473ad6eff2b8131cd7c68d2532e9374e295ed7f4a6c25fe2e272ad55e88f0519c3cda2049bf0ead7d8d07cb6dab8e494243910ce78ce9e74237eeea86e99f150bbd664a33c55ad2e1a5215f7cdcc6211a0fca0824b13c7d3fc9e2a3db98013fb2341d0d351ba0013cf06eb7b7459ae114048a1abdbbbb5130bf2f19980b917e372e5f0e9d20e7d87664979eac7f0bffe91a96c2622b4d1db67ea28ed359ddce6bbc8d5611641fc940fa1e3d2fa6c449c9dc7dc6e7c38cb683f81fd1fdb6c942aefc429ef39775ffd5d350acd4a6cb0f2fca84dece370a753b4de54e3097b5e6a5054d90a6b0c791e2a8da52b8e93fffa2fd05639e48c586a2fc5d57ac8c58e0d48bf88577dcb2c87cbacd03c776204a9945d4359a099d5107cc33452d33026bc351324143de46ce7e25723d4bd5c0df2b7089c6037a8095612d601b939ab626c4d456f8a22f373f92199a8b583f90a7f93ac5a8b58f616710241bc842255f8cb9067c055640a748b86f8bad386fc96fc1878272dfcd941e9abf0af26cc38535ac578dd9dc4084699950a6f6eae4339e5fbbc0e123e1e98451be46080c2e4243a8c8e9807c74c52d0507e5665a721e1a29563056e884235688516b0a9ffcd756bf5d54b016e99fddfb8fc2af600301239656d0076a5b124be7e574b1db9e785cb65998497c34775aad08b27d1b415096057dbb65a5a3ed71d9d5aadfb3a4a6adeb120b5c367d73aeecc7ba4f2dbd5bc8127f25829ad5ad9b70480750e84b38d5c27387d065a4bf380cab6c16332dfd501ab8578fe378cf0d17980dc308ca83912a334ac019a25e73a85de718cf99a06c1f44a6dcb0e67936a4726a261127154bdf93b94438441631393c0f59ef75bbfca27016ac7bf4f59cfff753eee96ec48f21246c8c74e2056bbd98f3382725943a904f897c34acb8f037df90d08afd6fe68a89a7a26bf0b2d7bec8aa15b10955958dc855284e764593a1d8056d061319e3e7fd36fea4ec074ea68183200c29a5ae89c73bac87d8741e4bf2299fea47ef42185742f6211d8653b4880c67b54d82c650ae197bdf149058180304042fd4802a4a5acefc7dd9403f12f6b2c9a08ed28542c6b835740f651027fc4eacbe2fd13e35950222e3c92425dcec742813e41926d5eb777d6156a64aab6830b4ccafe3b1417e073df1d89c832859a3da6f3604d8f4cb3df2a327321769522721ebad80bd03a73d4968d4ab0e4b8e46546422a6195d0409cd73911ea901f6d3e46f8e74fb1d5e09197170d2c2eee4d486a13b2f4645c86f8f8a5c78fccbbda659ba246ca9e04778ac585fad468080f8bc44f81f35cc68c3a0650fd4ca4f999f0c6b9413abf88946cbe9dc2f2a9e6e90557652f55da83bfa497703163ca8fbc2199f04fac77839659a6d681a88b07ddae829bce809eb5f2b54425f3af47afa98dd3afbbcd34aeab3f24ff80c087651ed227e497e297afe572e25b953932546998a445576252ed7e7c247b305e5f973b7c49fdca9de517873649b9656bcd573da5a5105df9e9c865bc4e5213ab9a1578d3b3a8c7e777ca0bec3d03071748b11078b052fd1c69b64a2c4f50187a8af9286f71c5e14d0bb9ba9493e4d85c77d0513be7443c61c0b253a367bac3e41d4b852ae76bc47c69fd5352512bd64d6b15bb4d4721b18cfb7dab6e3e2ce8dbc49cd8b564b5a3e92305f476c7153ba580de0cea6f3b5dbdb7e6cdee9fd18abe362af57ffac429467f4b424a3b606c4050b650da526ab067673a2dc0e7b860c0d9b9f497928898c7c3e965c954f853a8fe243a2d9212b4989712758f3aa508670ab2753be319e8b38371f04d11f046aac9e6ca4e0f12fc02bc7e3f97315fc9284661f728f1cf241fa372aa9da4bae56b17fce185daa83c4f597ac34327c0d82a8621b4ccaf0bf80c6a7b134c9b3cdf98a5ec0337964764ecf0412bc427bf9b0b6c778168b7b9bbe5232407805d931a5a1b267783142e9c2a2a86a5aebf747a9126afef46c44ad5860065f92668bdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h94e17ea933643279335a574b98ac74de991ce710e5e3d8268dac253d7640f82d4527d57e128eb68f1bc1a176f48258eaab4f1ebebc705a6f5d5fbf9d71c8b826b2a1e632eec4764ea22a5fb047788e3d48420b4fa5f492e2c5e0b6eb4bbf3562206eb5e9cb4c1aa87c80168e940cb5147a016a742a2a4f13cee16826b9c31ceab781b31ac893afabd1fc3ba38e0130d2b55a179596719912300c0888f490d991ee521976e170586e77eaa9b9fa833e4900d4b476212ff8c6ea0382028033d7251f325cd860e7819d6402fb9705ea59f3c18187cfb7ec86a073e35d489c2f1e1ed96387646aff0908bd66270341a958f7c00b31232934ca4f131ca3702029a6ddab5db7860133b6e597833e7a7e4cd92932209c57a1f8aea894a014f28a55fc3237cd8d8e777488a6265ced87826350e3ed4042ac7f7cfc061fb11c51f9b0e7606316f1b009be814de985a83d1ba4a99865ec7fc4e416ebce8af8278b7944fd0b2702bc759c60297dc339f417a023847aabd8d1a938320e4657e74667196fefcf3f8007212a018a1dfd861ea630c93ed36601babafa261604b16a16e5f1342d4580d0263c3e51ba9fb506d593b2ffb5a0bdfcadc418fbcf449beda12cc1eda62e8f149df9052fd3db60b55b8c7aaa24d451bcb64f3d44b1c7756e6ad62329172416ec067916829ed2ed64d76753b10d2c5ef9a8023b1dc88d7c0cec678efd84f43eef0e0fd36b5d52c5c19ba106d066271609da2ac544c84189c35f037684073a5fe2788414ff5fd6791f5d644e7324b2fb1e831b026b5dbe1674c88bf94a5addfa006aadf4b7d544883c1404034770763081a753d8cf8aac9473d90d141a3ab1d691ca558767a2443cdb9a1ace0e5fd894738f109d7adf3b3a0b7b15609aeb9a670b3a294623d29907e585b52916700268db67cffb17964ba23e8f7cc138460ae5f1465a2bf3a12c2832aa8b7e5d20243e9d7233aa765bc494917c20ec58f7b65f0a8a92a3e4f1a93fc41a8126f048dfaf40b2e8e67c1c26e6e523dde56f391a21b7663e26b22547fdd5b0bad73f0a9c7b9f487c36d006e207ca08409cfe233acd9aa2ef56926e5a83a90f84eb5bf7622ada00d46fd9aa8c275fa8302cc2327122e14c7d28998cfa77c0d57a06760c36725af9723a63ca09467c359220230ee4dad67aa49f970d3065ce37b7bba687dd337d6093fbaac9d07b87a331f258ba2612df019961fbe357e9b234c71029cfde34438e068704eb8f9403e709fcbccba1774479d9ed941668d60e2fc249d05775716a74cb37930168c561626b3c251d8c0043bf50c24ed6912b744b4e86d7ee7b49a8b128a152212cc3c2ef97713b4e061a0fc8be6423158736d7b72e467246133ef41c88276ba0ea50773c4f7ef0d7873a84f7781dc7d116e502b081f48bf124b509f3e05cb318fbe3ad3f0b0cf9039374d079511225445dcf54d7886e7022b08e2d962f7d79122e760f30435c8fb99c65ee906227117aee6b7729bd116fc34fce5501f2ad0c00517736923d50f27c0612f77dfce1f4c287f751affa1b446159d0fb20c34dac5e8c207721b5b77289ba04c1fe9ffac04601941d0ade0353f9e317a6aff3d2600e11eac9dcc74734f6eb0fc44a113244ce8adadf887010f4378ccee693cd9bd53a50d8798090db3e3c0b4d11192db93de397e406e6344756f1488a29f06b59cb9efbca272bb2ba041666008abfa1602d6c3d9387f4f6f48330e5efbcea85434adcfd48364b3137085d7c64fe2eaa485c371dadd3475274a884707602d7682453e179d2646ab8c38ae36c29d19cd73de8c0d0e62ed1ff2ee3ea044ba5b8b1f82d297da33a32ab12c5a5c62a6ccc170e513910b7bdf8412acceff1f42f152e9eb7ff3440ee7b351d516bbb110138d509b26e13cc61c729f4d64e2234d3ad64a642138cfd0baac9c3274eb70831371cad3eaf85285872c0b4a9878c83ad3b62da4ece9d1c8f1bd78ff4d653578bc534323c7a94875d588d9ce33f1d2840644bd49ea2bc690a09a7b0714601223e21f6feecda08da7d8569eee1ca27f31a708b82b3259a83de6c723fa787187aabd034c2755892275ddf9388dd65c5838f29a4f740ea4b0d793a32ac6902f9577d124255832c963d75b910a89568209ee4f1f0973b3cacbc2e72fb962f9730eec1508fd2fb8c134cca4aee0b90e3ef75f384d8a571b25e3d1d87dca6011fa802c8d119ecded0594cb14dfcae24c3144ed2dde120315c4dec7d6c3e29a63b356beda29bf3f443b4dbddb6c28d6589a99ecf045af8f9d14204caa874c4f849c87d7f23eeb212f79f33d11e397d484ca3b7ec00479a3ef5a73ba9496234dfbcb4bc340c62326ea9c54a2f6ae1f0032dc7ec993ba315c10cd4468b3af6051dcff0975ddc4fa90b7436d04731872485f16aa54152dc7d16fd2eeed664b4f62cd9b04a94a034bf48a9cddb08d09303b2bac2c4d054cca7c6fa4a0f7ea2931293c732fcb7f1093dd3e30d4a9271f3ad28d6292957fa9b74dd303220437bb81b2c43e5007ad57008c945f3d2413868633bfd14f4738b9c4455f83b1fa406d74b95c601a8f7c29c0a032150b9fba40f47bb6d81d293cc8de6180ee810444327871b5075be81817a448528c089eb47555177d5806fef1f0f32a15ddc0ee0799e4aa64c7cf742bf8efa4840685c549591092c256c812443eefe209f3c29a8ca3331d0e2ae2f427d8964813b6e8a6b6fc992fde37d735a68a33b6514c7aa39db663ac960cb4421dc4a1a4788f1032a393a81948fc9a3ef142f4125b230c5694ae27a5d72067b37633a3eb4fbed9a11f2e620d34fbf327218117f6b6822a9fcd03c695acc3c11e78069ef7fb86d528c0cb8401312176da36482accb11e7f324e2c2cf263bc0;
        #1
        $finish();
    end
endmodule
