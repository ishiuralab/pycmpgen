module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    compressor_CLA486_16 compressor_CLA486_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA486_16(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [147:0] stage1_0;
   wire [134:0] stage1_1;
   wire [167:0] stage1_2;
   wire [243:0] stage1_3;
   wire [222:0] stage1_4;
   wire [336:0] stage1_5;
   wire [196:0] stage1_6;
   wire [216:0] stage1_7;
   wire [195:0] stage1_8;
   wire [210:0] stage1_9;
   wire [281:0] stage1_10;
   wire [213:0] stage1_11;
   wire [201:0] stage1_12;
   wire [234:0] stage1_13;
   wire [182:0] stage1_14;
   wire [154:0] stage1_15;
   wire [150:0] stage1_16;
   wire [80:0] stage1_17;
   wire [37:0] stage2_0;
   wire [62:0] stage2_1;
   wire [53:0] stage2_2;
   wire [85:0] stage2_3;
   wire [106:0] stage2_4;
   wire [107:0] stage2_5;
   wire [89:0] stage2_6;
   wire [102:0] stage2_7;
   wire [105:0] stage2_8;
   wire [80:0] stage2_9;
   wire [89:0] stage2_10;
   wire [106:0] stage2_11;
   wire [93:0] stage2_12;
   wire [85:0] stage2_13;
   wire [101:0] stage2_14;
   wire [74:0] stage2_15;
   wire [76:0] stage2_16;
   wire [95:0] stage2_17;
   wire [25:0] stage2_18;
   wire [4:0] stage2_19;
   wire [19:0] stage3_0;
   wire [14:0] stage3_1;
   wire [18:0] stage3_2;
   wire [40:0] stage3_3;
   wire [38:0] stage3_4;
   wire [39:0] stage3_5;
   wire [49:0] stage3_6;
   wire [35:0] stage3_7;
   wire [47:0] stage3_8;
   wire [42:0] stage3_9;
   wire [43:0] stage3_10;
   wire [37:0] stage3_11;
   wire [46:0] stage3_12;
   wire [39:0] stage3_13;
   wire [31:0] stage3_14;
   wire [43:0] stage3_15;
   wire [44:0] stage3_16;
   wire [29:0] stage3_17;
   wire [25:0] stage3_18;
   wire [18:0] stage3_19;
   wire [4:0] stage3_20;
   wire [0:0] stage3_21;
   wire [9:0] stage4_0;
   wire [5:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [20:0] stage4_7;
   wire [19:0] stage4_8;
   wire [15:0] stage4_9;
   wire [17:0] stage4_10;
   wire [18:0] stage4_11;
   wire [23:0] stage4_12;
   wire [16:0] stage4_13;
   wire [19:0] stage4_14;
   wire [27:0] stage4_15;
   wire [18:0] stage4_16;
   wire [12:0] stage4_17;
   wire [24:0] stage4_18;
   wire [13:0] stage4_19;
   wire [8:0] stage4_20;
   wire [2:0] stage4_21;
   wire [9:0] stage5_0;
   wire [5:0] stage5_1;
   wire [8:0] stage5_2;
   wire [5:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [8:0] stage5_6;
   wire [8:0] stage5_7;
   wire [13:0] stage5_8;
   wire [8:0] stage5_9;
   wire [7:0] stage5_10;
   wire [6:0] stage5_11;
   wire [6:0] stage5_12;
   wire [9:0] stage5_13;
   wire [7:0] stage5_14;
   wire [9:0] stage5_15;
   wire [9:0] stage5_16;
   wire [7:0] stage5_17;
   wire [6:0] stage5_18;
   wire [10:0] stage5_19;
   wire [11:0] stage5_20;
   wire [3:0] stage5_21;
   wire [0:0] stage5_22;
   wire [5:0] stage6_0;
   wire [3:0] stage6_1;
   wire [4:0] stage6_2;
   wire [2:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [2:0] stage6_6;
   wire [3:0] stage6_7;
   wire [3:0] stage6_8;
   wire [5:0] stage6_9;
   wire [4:0] stage6_10;
   wire [2:0] stage6_11;
   wire [1:0] stage6_12;
   wire [6:0] stage6_13;
   wire [3:0] stage6_14;
   wire [2:0] stage6_15;
   wire [5:0] stage6_16;
   wire [2:0] stage6_17;
   wire [5:0] stage6_18;
   wire [3:0] stage6_19;
   wire [4:0] stage6_20;
   wire [2:0] stage6_21;
   wire [2:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [0:0] stage7_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_2[24]},
      {stage0_3[36]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_2[25]},
      {stage0_3[37]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_2[26]},
      {stage0_3[38]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_2[27]},
      {stage0_3[39]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_2[28]},
      {stage0_3[40]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_2[29]},
      {stage0_3[41]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_2[30]},
      {stage0_3[42]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_2[31]},
      {stage0_3[43]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_2[32]},
      {stage0_3[44]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_2[33]},
      {stage0_3[45]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_2[34]},
      {stage0_3[46]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_2[35]},
      {stage0_3[47]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_2[36]},
      {stage0_3[48]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[0],stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[1],stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[2],stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[3],stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[4],stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[5],stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[6],stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[7],stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[8],stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[9],stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[10],stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[11],stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[12],stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[13],stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[14],stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[15],stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[16],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[17],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[18],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[19],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[20],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[21],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[22],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[23],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[24],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[25],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[26],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[27],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[28],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[29],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[30],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[31],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[32],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[33],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[34],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[35],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[36],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[37],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[38],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[39],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[40],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[41],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[42],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312]},
      {stage1_5[43],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage1_5[44],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324]},
      {stage1_5[45],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage1_5[46],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage1_5[47],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342]},
      {stage1_5[48],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage1_5[49],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[50],stage1_4[135],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[51],stage1_4[136],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[52],stage1_4[137],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[53],stage1_4[138],stage1_3[138],stage1_2[138]}
   );
   gpc615_5 gpc139 (
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_3[349]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[54],stage1_4[139],stage1_3[139],stage1_2[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358]},
      {stage0_3[350]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[55],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363]},
      {stage0_3[351]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[56],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_3[352]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[57],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373]},
      {stage0_3[353]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[58],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage0_3[354]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[59],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_3[355]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[60],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388]},
      {stage0_3[356]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[61],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393]},
      {stage0_3[357]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[62],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage0_3[358]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[63],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403]},
      {stage0_3[359]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[64],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage0_3[360]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[65],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_3[361]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[66],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418]},
      {stage0_3[362]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[67],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423]},
      {stage0_3[363]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[68],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage0_3[364]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[69],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432], stage0_2[433]},
      {stage0_3[365]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[70],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437], stage0_2[438]},
      {stage0_3[366]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[71],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_3[367]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[72],stage1_4[157],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448]},
      {stage0_3[368]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[73],stage1_4[158],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453]},
      {stage0_3[369]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[74],stage1_4[159],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457], stage0_2[458]},
      {stage0_3[370]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[75],stage1_4[160],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462], stage0_2[463]},
      {stage0_3[371]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[76],stage1_4[161],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467], stage0_2[468]},
      {stage0_3[372]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[77],stage1_4[162],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_3[373]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[78],stage1_4[163],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478]},
      {stage0_3[374]},
      {stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179]},
      {stage1_6[29],stage1_5[79],stage1_4[164],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483]},
      {stage0_3[375]},
      {stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185]},
      {stage1_6[30],stage1_5[80],stage1_4[165],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[186]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[31],stage1_5[81],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[187]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[32],stage1_5[82],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[188]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[33],stage1_5[83],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[189]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[34],stage1_5[84],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[190]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[35],stage1_5[85],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[191]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[36],stage1_5[86],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[192]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[37],stage1_5[87],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[193]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[38],stage1_5[88],stage1_4[173],stage1_3[173]}
   );
   gpc606_5 gpc174 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[39],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc175 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[40],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc176 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[41],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc177 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[42],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc178 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[43],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[44],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[45],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[46],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[47],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[48],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[49],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[50],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[51],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[52],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[53],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[54],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[55],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[56],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[57],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[27],stage1_6[58],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[28],stage1_6[59],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[29],stage1_6[60],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[30],stage1_6[61],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[31],stage1_6[62],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[32],stage1_6[63],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[33],stage1_6[64],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[34],stage1_6[65],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[35],stage1_6[66],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[36],stage1_6[67],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[37],stage1_6[68],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[38],stage1_6[69],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[39],stage1_6[70],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[40],stage1_6[71],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[41],stage1_6[72],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[42],stage1_6[73],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[43],stage1_6[74],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[44],stage1_6[75],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[45],stage1_6[76],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[46],stage1_6[77],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[47],stage1_6[78],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[48],stage1_6[79],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[49],stage1_6[80],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[50],stage1_6[81],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[51],stage1_6[82],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[52],stage1_6[83],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[53],stage1_6[84],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[54],stage1_6[85],stage1_5[135],stage1_4[220]}
   );
   gpc615_5 gpc221 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[48]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[55],stage1_6[86],stage1_5[136],stage1_4[221]}
   );
   gpc615_5 gpc222 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485]},
      {stage0_5[49]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[56],stage1_6[87],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[49],stage1_7[57],stage1_6[88],stage1_5[138]}
   );
   gpc606_5 gpc224 (
      {stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[50],stage1_7[58],stage1_6[89],stage1_5[139]}
   );
   gpc606_5 gpc225 (
      {stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[51],stage1_7[59],stage1_6[90],stage1_5[140]}
   );
   gpc606_5 gpc226 (
      {stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[52],stage1_7[60],stage1_6[91],stage1_5[141]}
   );
   gpc606_5 gpc227 (
      {stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[53],stage1_7[61],stage1_6[92],stage1_5[142]}
   );
   gpc606_5 gpc228 (
      {stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[54],stage1_7[62],stage1_6[93],stage1_5[143]}
   );
   gpc606_5 gpc229 (
      {stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[55],stage1_7[63],stage1_6[94],stage1_5[144]}
   );
   gpc606_5 gpc230 (
      {stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[56],stage1_7[64],stage1_6[95],stage1_5[145]}
   );
   gpc606_5 gpc231 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[57],stage1_7[65],stage1_6[96],stage1_5[146]}
   );
   gpc606_5 gpc232 (
      {stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[58],stage1_7[66],stage1_6[97],stage1_5[147]}
   );
   gpc606_5 gpc233 (
      {stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[59],stage1_7[67],stage1_6[98],stage1_5[148]}
   );
   gpc606_5 gpc234 (
      {stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[60],stage1_7[68],stage1_6[99],stage1_5[149]}
   );
   gpc606_5 gpc235 (
      {stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[61],stage1_7[69],stage1_6[100],stage1_5[150]}
   );
   gpc606_5 gpc236 (
      {stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[62],stage1_7[70],stage1_6[101],stage1_5[151]}
   );
   gpc606_5 gpc237 (
      {stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[63],stage1_7[71],stage1_6[102],stage1_5[152]}
   );
   gpc606_5 gpc238 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[64],stage1_7[72],stage1_6[103],stage1_5[153]}
   );
   gpc606_5 gpc239 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[65],stage1_7[73],stage1_6[104],stage1_5[154]}
   );
   gpc606_5 gpc240 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[66],stage1_7[74],stage1_6[105],stage1_5[155]}
   );
   gpc606_5 gpc241 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[67],stage1_7[75],stage1_6[106],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[68],stage1_7[76],stage1_6[107],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[69],stage1_7[77],stage1_6[108],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[70],stage1_7[78],stage1_6[109],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[71],stage1_7[79],stage1_6[110],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[72],stage1_7[80],stage1_6[111],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[73],stage1_7[81],stage1_6[112],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[74],stage1_7[82],stage1_6[113],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[75],stage1_7[83],stage1_6[114],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[76],stage1_7[84],stage1_6[115],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[77],stage1_7[85],stage1_6[116],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[78],stage1_7[86],stage1_6[117],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[79],stage1_7[87],stage1_6[118],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[80],stage1_7[88],stage1_6[119],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[81],stage1_7[89],stage1_6[120],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[82],stage1_7[90],stage1_6[121],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[83],stage1_7[91],stage1_6[122],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[84],stage1_7[92],stage1_6[123],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[85],stage1_7[93],stage1_6[124],stage1_5[174]}
   );
   gpc615_5 gpc260 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_6[294]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[86],stage1_7[94],stage1_6[125],stage1_5[175]}
   );
   gpc615_5 gpc261 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_6[295]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[87],stage1_7[95],stage1_6[126],stage1_5[176]}
   );
   gpc615_5 gpc262 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286]},
      {stage0_6[296]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[88],stage1_7[96],stage1_6[127],stage1_5[177]}
   );
   gpc615_5 gpc263 (
      {stage0_5[287], stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291]},
      {stage0_6[297]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[89],stage1_7[97],stage1_6[128],stage1_5[178]}
   );
   gpc615_5 gpc264 (
      {stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295], stage0_5[296]},
      {stage0_6[298]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[90],stage1_7[98],stage1_6[129],stage1_5[179]}
   );
   gpc615_5 gpc265 (
      {stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_6[299]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[91],stage1_7[99],stage1_6[130],stage1_5[180]}
   );
   gpc615_5 gpc266 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_6[300]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[92],stage1_7[100],stage1_6[131],stage1_5[181]}
   );
   gpc615_5 gpc267 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_6[301]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[93],stage1_7[101],stage1_6[132],stage1_5[182]}
   );
   gpc615_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316]},
      {stage0_6[302]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[94],stage1_7[102],stage1_6[133],stage1_5[183]}
   );
   gpc615_5 gpc269 (
      {stage0_5[317], stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321]},
      {stage0_6[303]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[95],stage1_7[103],stage1_6[134],stage1_5[184]}
   );
   gpc615_5 gpc270 (
      {stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325], stage0_5[326]},
      {stage0_6[304]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[96],stage1_7[104],stage1_6[135],stage1_5[185]}
   );
   gpc615_5 gpc271 (
      {stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_6[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[97],stage1_7[105],stage1_6[136],stage1_5[186]}
   );
   gpc615_5 gpc272 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_6[306]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[98],stage1_7[106],stage1_6[137],stage1_5[187]}
   );
   gpc615_5 gpc273 (
      {stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[99],stage1_7[107],stage1_6[138]}
   );
   gpc615_5 gpc274 (
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[100],stage1_7[108],stage1_6[139]}
   );
   gpc615_5 gpc275 (
      {stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[101],stage1_7[109],stage1_6[140]}
   );
   gpc615_5 gpc276 (
      {stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325], stage0_6[326]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[102],stage1_7[110],stage1_6[141]}
   );
   gpc615_5 gpc277 (
      {stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330], stage0_6[331]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[103],stage1_7[111],stage1_6[142]}
   );
   gpc615_5 gpc278 (
      {stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335], stage0_6[336]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[104],stage1_7[112],stage1_6[143]}
   );
   gpc615_5 gpc279 (
      {stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[105],stage1_7[113],stage1_6[144]}
   );
   gpc615_5 gpc280 (
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[106],stage1_7[114],stage1_6[145]}
   );
   gpc615_5 gpc281 (
      {stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[107],stage1_7[115],stage1_6[146]}
   );
   gpc615_5 gpc282 (
      {stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355], stage0_6[356]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[108],stage1_7[116],stage1_6[147]}
   );
   gpc615_5 gpc283 (
      {stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360], stage0_6[361]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[109],stage1_7[117],stage1_6[148]}
   );
   gpc615_5 gpc284 (
      {stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365], stage0_6[366]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[110],stage1_7[118],stage1_6[149]}
   );
   gpc615_5 gpc285 (
      {stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[111],stage1_7[119],stage1_6[150]}
   );
   gpc615_5 gpc286 (
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[112],stage1_7[120],stage1_6[151]}
   );
   gpc615_5 gpc287 (
      {stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[113],stage1_7[121],stage1_6[152]}
   );
   gpc615_5 gpc288 (
      {stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385], stage0_6[386]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[114],stage1_7[122],stage1_6[153]}
   );
   gpc615_5 gpc289 (
      {stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390], stage0_6[391]},
      {stage0_7[316]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[66],stage1_8[115],stage1_7[123],stage1_6[154]}
   );
   gpc615_5 gpc290 (
      {stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395], stage0_6[396]},
      {stage0_7[317]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[67],stage1_8[116],stage1_7[124],stage1_6[155]}
   );
   gpc615_5 gpc291 (
      {stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage0_7[318]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[68],stage1_8[117],stage1_7[125],stage1_6[156]}
   );
   gpc615_5 gpc292 (
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406]},
      {stage0_7[319]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[69],stage1_8[118],stage1_7[126],stage1_6[157]}
   );
   gpc615_5 gpc293 (
      {stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411]},
      {stage0_7[320]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[70],stage1_8[119],stage1_7[127],stage1_6[158]}
   );
   gpc615_5 gpc294 (
      {stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415], stage0_6[416]},
      {stage0_7[321]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[71],stage1_8[120],stage1_7[128],stage1_6[159]}
   );
   gpc615_5 gpc295 (
      {stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420], stage0_6[421]},
      {stage0_7[322]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[72],stage1_8[121],stage1_7[129],stage1_6[160]}
   );
   gpc615_5 gpc296 (
      {stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425], stage0_6[426]},
      {stage0_7[323]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[73],stage1_8[122],stage1_7[130],stage1_6[161]}
   );
   gpc615_5 gpc297 (
      {stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage0_7[324]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[74],stage1_8[123],stage1_7[131],stage1_6[162]}
   );
   gpc615_5 gpc298 (
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436]},
      {stage0_7[325]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[75],stage1_8[124],stage1_7[132],stage1_6[163]}
   );
   gpc615_5 gpc299 (
      {stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441]},
      {stage0_7[326]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[76],stage1_8[125],stage1_7[133],stage1_6[164]}
   );
   gpc615_5 gpc300 (
      {stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445], stage0_6[446]},
      {stage0_7[327]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[77],stage1_8[126],stage1_7[134],stage1_6[165]}
   );
   gpc615_5 gpc301 (
      {stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450], stage0_6[451]},
      {stage0_7[328]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[78],stage1_8[127],stage1_7[135],stage1_6[166]}
   );
   gpc615_5 gpc302 (
      {stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455], stage0_6[456]},
      {stage0_7[329]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[79],stage1_8[128],stage1_7[136],stage1_6[167]}
   );
   gpc615_5 gpc303 (
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334]},
      {stage0_8[180]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[30],stage1_9[80],stage1_8[129],stage1_7[137]}
   );
   gpc615_5 gpc304 (
      {stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339]},
      {stage0_8[181]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[31],stage1_9[81],stage1_8[130],stage1_7[138]}
   );
   gpc615_5 gpc305 (
      {stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344]},
      {stage0_8[182]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[32],stage1_9[82],stage1_8[131],stage1_7[139]}
   );
   gpc615_5 gpc306 (
      {stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349]},
      {stage0_8[183]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[33],stage1_9[83],stage1_8[132],stage1_7[140]}
   );
   gpc615_5 gpc307 (
      {stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354]},
      {stage0_8[184]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[34],stage1_9[84],stage1_8[133],stage1_7[141]}
   );
   gpc615_5 gpc308 (
      {stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage0_8[185]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[35],stage1_9[85],stage1_8[134],stage1_7[142]}
   );
   gpc615_5 gpc309 (
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_8[186]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[36],stage1_9[86],stage1_8[135],stage1_7[143]}
   );
   gpc615_5 gpc310 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369]},
      {stage0_8[187]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[37],stage1_9[87],stage1_8[136],stage1_7[144]}
   );
   gpc615_5 gpc311 (
      {stage0_7[370], stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374]},
      {stage0_8[188]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[38],stage1_9[88],stage1_8[137],stage1_7[145]}
   );
   gpc615_5 gpc312 (
      {stage0_7[375], stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379]},
      {stage0_8[189]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[39],stage1_9[89],stage1_8[138],stage1_7[146]}
   );
   gpc615_5 gpc313 (
      {stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384]},
      {stage0_8[190]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[40],stage1_9[90],stage1_8[139],stage1_7[147]}
   );
   gpc615_5 gpc314 (
      {stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage0_8[191]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[41],stage1_9[91],stage1_8[140],stage1_7[148]}
   );
   gpc615_5 gpc315 (
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_8[192]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[42],stage1_9[92],stage1_8[141],stage1_7[149]}
   );
   gpc615_5 gpc316 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399]},
      {stage0_8[193]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[43],stage1_9[93],stage1_8[142],stage1_7[150]}
   );
   gpc615_5 gpc317 (
      {stage0_7[400], stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404]},
      {stage0_8[194]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[44],stage1_9[94],stage1_8[143],stage1_7[151]}
   );
   gpc615_5 gpc318 (
      {stage0_7[405], stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409]},
      {stage0_8[195]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[45],stage1_9[95],stage1_8[144],stage1_7[152]}
   );
   gpc615_5 gpc319 (
      {stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414]},
      {stage0_8[196]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[46],stage1_9[96],stage1_8[145],stage1_7[153]}
   );
   gpc615_5 gpc320 (
      {stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage0_8[197]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[47],stage1_9[97],stage1_8[146],stage1_7[154]}
   );
   gpc615_5 gpc321 (
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_8[198]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[48],stage1_9[98],stage1_8[147],stage1_7[155]}
   );
   gpc606_5 gpc322 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[19],stage1_10[49],stage1_9[99],stage1_8[148]}
   );
   gpc606_5 gpc323 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[20],stage1_10[50],stage1_9[100],stage1_8[149]}
   );
   gpc606_5 gpc324 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[21],stage1_10[51],stage1_9[101],stage1_8[150]}
   );
   gpc606_5 gpc325 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[22],stage1_10[52],stage1_9[102],stage1_8[151]}
   );
   gpc606_5 gpc326 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[23],stage1_10[53],stage1_9[103],stage1_8[152]}
   );
   gpc606_5 gpc327 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[24],stage1_10[54],stage1_9[104],stage1_8[153]}
   );
   gpc606_5 gpc328 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[25],stage1_10[55],stage1_9[105],stage1_8[154]}
   );
   gpc606_5 gpc329 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[26],stage1_10[56],stage1_9[106],stage1_8[155]}
   );
   gpc606_5 gpc330 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[27],stage1_10[57],stage1_9[107],stage1_8[156]}
   );
   gpc606_5 gpc331 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[28],stage1_10[58],stage1_9[108],stage1_8[157]}
   );
   gpc606_5 gpc332 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[29],stage1_10[59],stage1_9[109],stage1_8[158]}
   );
   gpc606_5 gpc333 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[30],stage1_10[60],stage1_9[110],stage1_8[159]}
   );
   gpc606_5 gpc334 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[31],stage1_10[61],stage1_9[111],stage1_8[160]}
   );
   gpc606_5 gpc335 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[32],stage1_10[62],stage1_9[112],stage1_8[161]}
   );
   gpc606_5 gpc336 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[33],stage1_10[63],stage1_9[113],stage1_8[162]}
   );
   gpc606_5 gpc337 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[34],stage1_10[64],stage1_9[114],stage1_8[163]}
   );
   gpc606_5 gpc338 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[35],stage1_10[65],stage1_9[115],stage1_8[164]}
   );
   gpc606_5 gpc339 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[36],stage1_10[66],stage1_9[116],stage1_8[165]}
   );
   gpc606_5 gpc340 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[37],stage1_10[67],stage1_9[117],stage1_8[166]}
   );
   gpc606_5 gpc341 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[38],stage1_10[68],stage1_9[118],stage1_8[167]}
   );
   gpc606_5 gpc342 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[39],stage1_10[69],stage1_9[119],stage1_8[168]}
   );
   gpc606_5 gpc343 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[40],stage1_10[70],stage1_9[120],stage1_8[169]}
   );
   gpc606_5 gpc344 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[41],stage1_10[71],stage1_9[121],stage1_8[170]}
   );
   gpc606_5 gpc345 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[42],stage1_10[72],stage1_9[122],stage1_8[171]}
   );
   gpc606_5 gpc346 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[43],stage1_10[73],stage1_9[123],stage1_8[172]}
   );
   gpc606_5 gpc347 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[44],stage1_10[74],stage1_9[124],stage1_8[173]}
   );
   gpc606_5 gpc348 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[45],stage1_10[75],stage1_9[125],stage1_8[174]}
   );
   gpc606_5 gpc349 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[46],stage1_10[76],stage1_9[126],stage1_8[175]}
   );
   gpc606_5 gpc350 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[47],stage1_10[77],stage1_9[127],stage1_8[176]}
   );
   gpc606_5 gpc351 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[48],stage1_10[78],stage1_9[128],stage1_8[177]}
   );
   gpc606_5 gpc352 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[49],stage1_10[79],stage1_9[129],stage1_8[178]}
   );
   gpc606_5 gpc353 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[50],stage1_10[80],stage1_9[130],stage1_8[179]}
   );
   gpc606_5 gpc354 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[51],stage1_10[81],stage1_9[131],stage1_8[180]}
   );
   gpc606_5 gpc355 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[52],stage1_10[82],stage1_9[132],stage1_8[181]}
   );
   gpc606_5 gpc356 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[53],stage1_10[83],stage1_9[133],stage1_8[182]}
   );
   gpc606_5 gpc357 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[54],stage1_10[84],stage1_9[134],stage1_8[183]}
   );
   gpc606_5 gpc358 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[55],stage1_10[85],stage1_9[135],stage1_8[184]}
   );
   gpc606_5 gpc359 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[56],stage1_10[86],stage1_9[136],stage1_8[185]}
   );
   gpc606_5 gpc360 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[57],stage1_10[87],stage1_9[137],stage1_8[186]}
   );
   gpc606_5 gpc361 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[58],stage1_10[88],stage1_9[138],stage1_8[187]}
   );
   gpc606_5 gpc362 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[59],stage1_10[89],stage1_9[139],stage1_8[188]}
   );
   gpc606_5 gpc363 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[60],stage1_10[90],stage1_9[140],stage1_8[189]}
   );
   gpc606_5 gpc364 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[61],stage1_10[91],stage1_9[141],stage1_8[190]}
   );
   gpc606_5 gpc365 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[62],stage1_10[92],stage1_9[142],stage1_8[191]}
   );
   gpc606_5 gpc366 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[63],stage1_10[93],stage1_9[143],stage1_8[192]}
   );
   gpc606_5 gpc367 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[64],stage1_10[94],stage1_9[144],stage1_8[193]}
   );
   gpc606_5 gpc368 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[65],stage1_10[95],stage1_9[145],stage1_8[194]}
   );
   gpc615_5 gpc369 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_9[114]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[66],stage1_10[96],stage1_9[146],stage1_8[195]}
   );
   gpc606_5 gpc370 (
      {stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[48],stage1_11[67],stage1_10[97],stage1_9[147]}
   );
   gpc606_5 gpc371 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[49],stage1_11[68],stage1_10[98],stage1_9[148]}
   );
   gpc606_5 gpc372 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[50],stage1_11[69],stage1_10[99],stage1_9[149]}
   );
   gpc606_5 gpc373 (
      {stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[51],stage1_11[70],stage1_10[100],stage1_9[150]}
   );
   gpc606_5 gpc374 (
      {stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[52],stage1_11[71],stage1_10[101],stage1_9[151]}
   );
   gpc606_5 gpc375 (
      {stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[53],stage1_11[72],stage1_10[102],stage1_9[152]}
   );
   gpc606_5 gpc376 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[54],stage1_11[73],stage1_10[103],stage1_9[153]}
   );
   gpc606_5 gpc377 (
      {stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[55],stage1_11[74],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc378 (
      {stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[56],stage1_11[75],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc379 (
      {stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[57],stage1_11[76],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc380 (
      {stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[58],stage1_11[77],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc381 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[59],stage1_11[78],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc382 (
      {stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[60],stage1_11[79],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc383 (
      {stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[61],stage1_11[80],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc384 (
      {stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[62],stage1_11[81],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc385 (
      {stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[63],stage1_11[82],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc386 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[64],stage1_11[83],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc387 (
      {stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[65],stage1_11[84],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc388 (
      {stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[66],stage1_11[85],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc389 (
      {stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[67],stage1_11[86],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc390 (
      {stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[68],stage1_11[87],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc391 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[69],stage1_11[88],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc392 (
      {stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[70],stage1_11[89],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc393 (
      {stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[71],stage1_11[90],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc394 (
      {stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[72],stage1_11[91],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc395 (
      {stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[73],stage1_11[92],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc396 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[74],stage1_11[93],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc397 (
      {stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[75],stage1_11[94],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc398 (
      {stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[76],stage1_11[95],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc399 (
      {stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[77],stage1_11[96],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc400 (
      {stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[78],stage1_11[97],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc401 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[79],stage1_11[98],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc402 (
      {stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[80],stage1_11[99],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc403 (
      {stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[81],stage1_11[100],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc404 (
      {stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[82],stage1_11[101],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc405 (
      {stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[83],stage1_11[102],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc406 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[84],stage1_11[103],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc407 (
      {stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[85],stage1_11[104],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc408 (
      {stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[86],stage1_11[105],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc409 (
      {stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[87],stage1_11[106],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc410 (
      {stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[88],stage1_11[107],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc411 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[89],stage1_11[108],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc412 (
      {stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[90],stage1_11[109],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc413 (
      {stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[91],stage1_11[110],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc414 (
      {stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[92],stage1_11[111],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc415 (
      {stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[93],stage1_11[112],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc416 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[94],stage1_11[113],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc417 (
      {stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[95],stage1_11[114],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc418 (
      {stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[96],stage1_11[115],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc419 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[97],stage1_11[116],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc420 (
      {stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[98],stage1_11[117],stage1_10[147],stage1_9[197]}
   );
   gpc615_5 gpc421 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[288]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[99],stage1_11[118],stage1_10[148],stage1_9[198]}
   );
   gpc615_5 gpc422 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[289]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[100],stage1_11[119],stage1_10[149],stage1_9[199]}
   );
   gpc615_5 gpc423 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[290]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[101],stage1_11[120],stage1_10[150],stage1_9[200]}
   );
   gpc615_5 gpc424 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[291]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[102],stage1_11[121],stage1_10[151],stage1_9[201]}
   );
   gpc615_5 gpc425 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[292]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[103],stage1_11[122],stage1_10[152],stage1_9[202]}
   );
   gpc615_5 gpc426 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[293]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[104],stage1_11[123],stage1_10[153],stage1_9[203]}
   );
   gpc615_5 gpc427 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[294]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[105],stage1_11[124],stage1_10[154],stage1_9[204]}
   );
   gpc615_5 gpc428 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[295]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[106],stage1_11[125],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc429 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[296]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[107],stage1_11[126],stage1_10[156],stage1_9[206]}
   );
   gpc615_5 gpc430 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[297]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[108],stage1_11[127],stage1_10[157],stage1_9[207]}
   );
   gpc615_5 gpc431 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[298]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[109],stage1_11[128],stage1_10[158],stage1_9[208]}
   );
   gpc615_5 gpc432 (
      {stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479], stage0_9[480]},
      {stage0_10[299]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[110],stage1_11[129],stage1_10[159],stage1_9[209]}
   );
   gpc615_5 gpc433 (
      {stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_10[300]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[111],stage1_11[130],stage1_10[160],stage1_9[210]}
   );
   gpc615_5 gpc434 (
      {stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage0_11[384]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[64],stage1_12[112],stage1_11[131],stage1_10[161]}
   );
   gpc615_5 gpc435 (
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310]},
      {stage0_11[385]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[65],stage1_12[113],stage1_11[132],stage1_10[162]}
   );
   gpc615_5 gpc436 (
      {stage0_10[311], stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315]},
      {stage0_11[386]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[66],stage1_12[114],stage1_11[133],stage1_10[163]}
   );
   gpc615_5 gpc437 (
      {stage0_10[316], stage0_10[317], stage0_10[318], stage0_10[319], stage0_10[320]},
      {stage0_11[387]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[67],stage1_12[115],stage1_11[134],stage1_10[164]}
   );
   gpc615_5 gpc438 (
      {stage0_10[321], stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325]},
      {stage0_11[388]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[68],stage1_12[116],stage1_11[135],stage1_10[165]}
   );
   gpc615_5 gpc439 (
      {stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329], stage0_10[330]},
      {stage0_11[389]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[69],stage1_12[117],stage1_11[136],stage1_10[166]}
   );
   gpc615_5 gpc440 (
      {stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[70],stage1_12[118],stage1_11[137],stage1_10[167]}
   );
   gpc615_5 gpc441 (
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[71],stage1_12[119],stage1_11[138],stage1_10[168]}
   );
   gpc615_5 gpc442 (
      {stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[72],stage1_12[120],stage1_11[139],stage1_10[169]}
   );
   gpc615_5 gpc443 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[73],stage1_12[121],stage1_11[140],stage1_10[170]}
   );
   gpc615_5 gpc444 (
      {stage0_10[351], stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[74],stage1_12[122],stage1_11[141],stage1_10[171]}
   );
   gpc615_5 gpc445 (
      {stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359], stage0_10[360]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[75],stage1_12[123],stage1_11[142],stage1_10[172]}
   );
   gpc615_5 gpc446 (
      {stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[76],stage1_12[124],stage1_11[143],stage1_10[173]}
   );
   gpc615_5 gpc447 (
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[77],stage1_12[125],stage1_11[144],stage1_10[174]}
   );
   gpc615_5 gpc448 (
      {stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[78],stage1_12[126],stage1_11[145],stage1_10[175]}
   );
   gpc615_5 gpc449 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[79],stage1_12[127],stage1_11[146],stage1_10[176]}
   );
   gpc2135_5 gpc450 (
      {stage0_11[400], stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404]},
      {stage0_12[96], stage0_12[97], stage0_12[98]},
      {stage0_13[0]},
      {stage0_14[0], stage0_14[1]},
      {stage1_15[0],stage1_14[16],stage1_13[80],stage1_12[128],stage1_11[147]}
   );
   gpc606_5 gpc451 (
      {stage0_11[405], stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5], stage0_13[6]},
      {stage1_15[1],stage1_14[17],stage1_13[81],stage1_12[129],stage1_11[148]}
   );
   gpc606_5 gpc452 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416]},
      {stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage1_15[2],stage1_14[18],stage1_13[82],stage1_12[130],stage1_11[149]}
   );
   gpc606_5 gpc453 (
      {stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422]},
      {stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18]},
      {stage1_15[3],stage1_14[19],stage1_13[83],stage1_12[131],stage1_11[150]}
   );
   gpc606_5 gpc454 (
      {stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7]},
      {stage1_16[0],stage1_15[4],stage1_14[20],stage1_13[84],stage1_12[132]}
   );
   gpc606_5 gpc455 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110]},
      {stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13]},
      {stage1_16[1],stage1_15[5],stage1_14[21],stage1_13[85],stage1_12[133]}
   );
   gpc606_5 gpc456 (
      {stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116]},
      {stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19]},
      {stage1_16[2],stage1_15[6],stage1_14[22],stage1_13[86],stage1_12[134]}
   );
   gpc606_5 gpc457 (
      {stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25]},
      {stage1_16[3],stage1_15[7],stage1_14[23],stage1_13[87],stage1_12[135]}
   );
   gpc606_5 gpc458 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128]},
      {stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31]},
      {stage1_16[4],stage1_15[8],stage1_14[24],stage1_13[88],stage1_12[136]}
   );
   gpc606_5 gpc459 (
      {stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134]},
      {stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36], stage0_14[37]},
      {stage1_16[5],stage1_15[9],stage1_14[25],stage1_13[89],stage1_12[137]}
   );
   gpc606_5 gpc460 (
      {stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140]},
      {stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42], stage0_14[43]},
      {stage1_16[6],stage1_15[10],stage1_14[26],stage1_13[90],stage1_12[138]}
   );
   gpc606_5 gpc461 (
      {stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49]},
      {stage1_16[7],stage1_15[11],stage1_14[27],stage1_13[91],stage1_12[139]}
   );
   gpc606_5 gpc462 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152]},
      {stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage1_16[8],stage1_15[12],stage1_14[28],stage1_13[92],stage1_12[140]}
   );
   gpc606_5 gpc463 (
      {stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158]},
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60], stage0_14[61]},
      {stage1_16[9],stage1_15[13],stage1_14[29],stage1_13[93],stage1_12[141]}
   );
   gpc606_5 gpc464 (
      {stage0_12[159], stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164]},
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67]},
      {stage1_16[10],stage1_15[14],stage1_14[30],stage1_13[94],stage1_12[142]}
   );
   gpc606_5 gpc465 (
      {stage0_12[165], stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169], stage0_12[170]},
      {stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73]},
      {stage1_16[11],stage1_15[15],stage1_14[31],stage1_13[95],stage1_12[143]}
   );
   gpc606_5 gpc466 (
      {stage0_12[171], stage0_12[172], stage0_12[173], stage0_12[174], stage0_12[175], stage0_12[176]},
      {stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79]},
      {stage1_16[12],stage1_15[16],stage1_14[32],stage1_13[96],stage1_12[144]}
   );
   gpc606_5 gpc467 (
      {stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182]},
      {stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83], stage0_14[84], stage0_14[85]},
      {stage1_16[13],stage1_15[17],stage1_14[33],stage1_13[97],stage1_12[145]}
   );
   gpc606_5 gpc468 (
      {stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89], stage0_14[90], stage0_14[91]},
      {stage1_16[14],stage1_15[18],stage1_14[34],stage1_13[98],stage1_12[146]}
   );
   gpc606_5 gpc469 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194]},
      {stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95], stage0_14[96], stage0_14[97]},
      {stage1_16[15],stage1_15[19],stage1_14[35],stage1_13[99],stage1_12[147]}
   );
   gpc606_5 gpc470 (
      {stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199], stage0_12[200]},
      {stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102], stage0_14[103]},
      {stage1_16[16],stage1_15[20],stage1_14[36],stage1_13[100],stage1_12[148]}
   );
   gpc606_5 gpc471 (
      {stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205], stage0_12[206]},
      {stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108], stage0_14[109]},
      {stage1_16[17],stage1_15[21],stage1_14[37],stage1_13[101],stage1_12[149]}
   );
   gpc606_5 gpc472 (
      {stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212]},
      {stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114], stage0_14[115]},
      {stage1_16[18],stage1_15[22],stage1_14[38],stage1_13[102],stage1_12[150]}
   );
   gpc606_5 gpc473 (
      {stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121]},
      {stage1_16[19],stage1_15[23],stage1_14[39],stage1_13[103],stage1_12[151]}
   );
   gpc606_5 gpc474 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223], stage0_12[224]},
      {stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage1_16[20],stage1_15[24],stage1_14[40],stage1_13[104],stage1_12[152]}
   );
   gpc606_5 gpc475 (
      {stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229], stage0_12[230]},
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132], stage0_14[133]},
      {stage1_16[21],stage1_15[25],stage1_14[41],stage1_13[105],stage1_12[153]}
   );
   gpc606_5 gpc476 (
      {stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236]},
      {stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage1_16[22],stage1_15[26],stage1_14[42],stage1_13[106],stage1_12[154]}
   );
   gpc606_5 gpc477 (
      {stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242]},
      {stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144], stage0_14[145]},
      {stage1_16[23],stage1_15[27],stage1_14[43],stage1_13[107],stage1_12[155]}
   );
   gpc606_5 gpc478 (
      {stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151]},
      {stage1_16[24],stage1_15[28],stage1_14[44],stage1_13[108],stage1_12[156]}
   );
   gpc606_5 gpc479 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254]},
      {stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage1_16[25],stage1_15[29],stage1_14[45],stage1_13[109],stage1_12[157]}
   );
   gpc606_5 gpc480 (
      {stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260]},
      {stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162], stage0_14[163]},
      {stage1_16[26],stage1_15[30],stage1_14[46],stage1_13[110],stage1_12[158]}
   );
   gpc606_5 gpc481 (
      {stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266]},
      {stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168], stage0_14[169]},
      {stage1_16[27],stage1_15[31],stage1_14[47],stage1_13[111],stage1_12[159]}
   );
   gpc606_5 gpc482 (
      {stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272]},
      {stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174], stage0_14[175]},
      {stage1_16[28],stage1_15[32],stage1_14[48],stage1_13[112],stage1_12[160]}
   );
   gpc606_5 gpc483 (
      {stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180], stage0_14[181]},
      {stage1_16[29],stage1_15[33],stage1_14[49],stage1_13[113],stage1_12[161]}
   );
   gpc606_5 gpc484 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284]},
      {stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186], stage0_14[187]},
      {stage1_16[30],stage1_15[34],stage1_14[50],stage1_13[114],stage1_12[162]}
   );
   gpc606_5 gpc485 (
      {stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290]},
      {stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192], stage0_14[193]},
      {stage1_16[31],stage1_15[35],stage1_14[51],stage1_13[115],stage1_12[163]}
   );
   gpc606_5 gpc486 (
      {stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296]},
      {stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198], stage0_14[199]},
      {stage1_16[32],stage1_15[36],stage1_14[52],stage1_13[116],stage1_12[164]}
   );
   gpc606_5 gpc487 (
      {stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302]},
      {stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204], stage0_14[205]},
      {stage1_16[33],stage1_15[37],stage1_14[53],stage1_13[117],stage1_12[165]}
   );
   gpc606_5 gpc488 (
      {stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210], stage0_14[211]},
      {stage1_16[34],stage1_15[38],stage1_14[54],stage1_13[118],stage1_12[166]}
   );
   gpc606_5 gpc489 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314]},
      {stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216], stage0_14[217]},
      {stage1_16[35],stage1_15[39],stage1_14[55],stage1_13[119],stage1_12[167]}
   );
   gpc606_5 gpc490 (
      {stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320]},
      {stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222], stage0_14[223]},
      {stage1_16[36],stage1_15[40],stage1_14[56],stage1_13[120],stage1_12[168]}
   );
   gpc615_5 gpc491 (
      {stage0_12[321], stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325]},
      {stage0_13[19]},
      {stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228], stage0_14[229]},
      {stage1_16[37],stage1_15[41],stage1_14[57],stage1_13[121],stage1_12[169]}
   );
   gpc615_5 gpc492 (
      {stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330]},
      {stage0_13[20]},
      {stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234], stage0_14[235]},
      {stage1_16[38],stage1_15[42],stage1_14[58],stage1_13[122],stage1_12[170]}
   );
   gpc615_5 gpc493 (
      {stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_13[21]},
      {stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239], stage0_14[240], stage0_14[241]},
      {stage1_16[39],stage1_15[43],stage1_14[59],stage1_13[123],stage1_12[171]}
   );
   gpc615_5 gpc494 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340]},
      {stage0_13[22]},
      {stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245], stage0_14[246], stage0_14[247]},
      {stage1_16[40],stage1_15[44],stage1_14[60],stage1_13[124],stage1_12[172]}
   );
   gpc615_5 gpc495 (
      {stage0_12[341], stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345]},
      {stage0_13[23]},
      {stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251], stage0_14[252], stage0_14[253]},
      {stage1_16[41],stage1_15[45],stage1_14[61],stage1_13[125],stage1_12[173]}
   );
   gpc615_5 gpc496 (
      {stage0_12[346], stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350]},
      {stage0_13[24]},
      {stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257], stage0_14[258], stage0_14[259]},
      {stage1_16[42],stage1_15[46],stage1_14[62],stage1_13[126],stage1_12[174]}
   );
   gpc615_5 gpc497 (
      {stage0_12[351], stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355]},
      {stage0_13[25]},
      {stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265]},
      {stage1_16[43],stage1_15[47],stage1_14[63],stage1_13[127],stage1_12[175]}
   );
   gpc615_5 gpc498 (
      {stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360]},
      {stage0_13[26]},
      {stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271]},
      {stage1_16[44],stage1_15[48],stage1_14[64],stage1_13[128],stage1_12[176]}
   );
   gpc615_5 gpc499 (
      {stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_13[27]},
      {stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277]},
      {stage1_16[45],stage1_15[49],stage1_14[65],stage1_13[129],stage1_12[177]}
   );
   gpc615_5 gpc500 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370]},
      {stage0_13[28]},
      {stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283]},
      {stage1_16[46],stage1_15[50],stage1_14[66],stage1_13[130],stage1_12[178]}
   );
   gpc615_5 gpc501 (
      {stage0_12[371], stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375]},
      {stage0_13[29]},
      {stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289]},
      {stage1_16[47],stage1_15[51],stage1_14[67],stage1_13[131],stage1_12[179]}
   );
   gpc615_5 gpc502 (
      {stage0_12[376], stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380]},
      {stage0_13[30]},
      {stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295]},
      {stage1_16[48],stage1_15[52],stage1_14[68],stage1_13[132],stage1_12[180]}
   );
   gpc615_5 gpc503 (
      {stage0_12[381], stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385]},
      {stage0_13[31]},
      {stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301]},
      {stage1_16[49],stage1_15[53],stage1_14[69],stage1_13[133],stage1_12[181]}
   );
   gpc615_5 gpc504 (
      {stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390]},
      {stage0_13[32]},
      {stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307]},
      {stage1_16[50],stage1_15[54],stage1_14[70],stage1_13[134],stage1_12[182]}
   );
   gpc615_5 gpc505 (
      {stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_13[33]},
      {stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage1_16[51],stage1_15[55],stage1_14[71],stage1_13[135],stage1_12[183]}
   );
   gpc615_5 gpc506 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400]},
      {stage0_13[34]},
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318], stage0_14[319]},
      {stage1_16[52],stage1_15[56],stage1_14[72],stage1_13[136],stage1_12[184]}
   );
   gpc615_5 gpc507 (
      {stage0_12[401], stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405]},
      {stage0_13[35]},
      {stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323], stage0_14[324], stage0_14[325]},
      {stage1_16[53],stage1_15[57],stage1_14[73],stage1_13[137],stage1_12[185]}
   );
   gpc615_5 gpc508 (
      {stage0_12[406], stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410]},
      {stage0_13[36]},
      {stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329], stage0_14[330], stage0_14[331]},
      {stage1_16[54],stage1_15[58],stage1_14[74],stage1_13[138],stage1_12[186]}
   );
   gpc615_5 gpc509 (
      {stage0_12[411], stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415]},
      {stage0_13[37]},
      {stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337]},
      {stage1_16[55],stage1_15[59],stage1_14[75],stage1_13[139],stage1_12[187]}
   );
   gpc615_5 gpc510 (
      {stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420]},
      {stage0_13[38]},
      {stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage1_16[56],stage1_15[60],stage1_14[76],stage1_13[140],stage1_12[188]}
   );
   gpc615_5 gpc511 (
      {stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_13[39]},
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348], stage0_14[349]},
      {stage1_16[57],stage1_15[61],stage1_14[77],stage1_13[141],stage1_12[189]}
   );
   gpc615_5 gpc512 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430]},
      {stage0_13[40]},
      {stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353], stage0_14[354], stage0_14[355]},
      {stage1_16[58],stage1_15[62],stage1_14[78],stage1_13[142],stage1_12[190]}
   );
   gpc615_5 gpc513 (
      {stage0_12[431], stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435]},
      {stage0_13[41]},
      {stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359], stage0_14[360], stage0_14[361]},
      {stage1_16[59],stage1_15[63],stage1_14[79],stage1_13[143],stage1_12[191]}
   );
   gpc615_5 gpc514 (
      {stage0_12[436], stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440]},
      {stage0_13[42]},
      {stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365], stage0_14[366], stage0_14[367]},
      {stage1_16[60],stage1_15[64],stage1_14[80],stage1_13[144],stage1_12[192]}
   );
   gpc615_5 gpc515 (
      {stage0_12[441], stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445]},
      {stage0_13[43]},
      {stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371], stage0_14[372], stage0_14[373]},
      {stage1_16[61],stage1_15[65],stage1_14[81],stage1_13[145],stage1_12[193]}
   );
   gpc615_5 gpc516 (
      {stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450]},
      {stage0_13[44]},
      {stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377], stage0_14[378], stage0_14[379]},
      {stage1_16[62],stage1_15[66],stage1_14[82],stage1_13[146],stage1_12[194]}
   );
   gpc615_5 gpc517 (
      {stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_13[45]},
      {stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383], stage0_14[384], stage0_14[385]},
      {stage1_16[63],stage1_15[67],stage1_14[83],stage1_13[147],stage1_12[195]}
   );
   gpc615_5 gpc518 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460]},
      {stage0_13[46]},
      {stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389], stage0_14[390], stage0_14[391]},
      {stage1_16[64],stage1_15[68],stage1_14[84],stage1_13[148],stage1_12[196]}
   );
   gpc615_5 gpc519 (
      {stage0_12[461], stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465]},
      {stage0_13[47]},
      {stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397]},
      {stage1_16[65],stage1_15[69],stage1_14[85],stage1_13[149],stage1_12[197]}
   );
   gpc615_5 gpc520 (
      {stage0_12[466], stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470]},
      {stage0_13[48]},
      {stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage1_16[66],stage1_15[70],stage1_14[86],stage1_13[150],stage1_12[198]}
   );
   gpc615_5 gpc521 (
      {stage0_12[471], stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475]},
      {stage0_13[49]},
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408], stage0_14[409]},
      {stage1_16[67],stage1_15[71],stage1_14[87],stage1_13[151],stage1_12[199]}
   );
   gpc615_5 gpc522 (
      {stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480]},
      {stage0_13[50]},
      {stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413], stage0_14[414], stage0_14[415]},
      {stage1_16[68],stage1_15[72],stage1_14[88],stage1_13[152],stage1_12[200]}
   );
   gpc615_5 gpc523 (
      {stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_13[51]},
      {stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419], stage0_14[420], stage0_14[421]},
      {stage1_16[69],stage1_15[73],stage1_14[89],stage1_13[153],stage1_12[201]}
   );
   gpc606_5 gpc524 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[70],stage1_15[74],stage1_14[90],stage1_13[154]}
   );
   gpc606_5 gpc525 (
      {stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[71],stage1_15[75],stage1_14[91],stage1_13[155]}
   );
   gpc606_5 gpc526 (
      {stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[72],stage1_15[76],stage1_14[92],stage1_13[156]}
   );
   gpc606_5 gpc527 (
      {stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[73],stage1_15[77],stage1_14[93],stage1_13[157]}
   );
   gpc606_5 gpc528 (
      {stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[74],stage1_15[78],stage1_14[94],stage1_13[158]}
   );
   gpc606_5 gpc529 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[75],stage1_15[79],stage1_14[95],stage1_13[159]}
   );
   gpc606_5 gpc530 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[76],stage1_15[80],stage1_14[96],stage1_13[160]}
   );
   gpc606_5 gpc531 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[77],stage1_15[81],stage1_14[97],stage1_13[161]}
   );
   gpc606_5 gpc532 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[78],stage1_15[82],stage1_14[98],stage1_13[162]}
   );
   gpc606_5 gpc533 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[79],stage1_15[83],stage1_14[99],stage1_13[163]}
   );
   gpc606_5 gpc534 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[80],stage1_15[84],stage1_14[100],stage1_13[164]}
   );
   gpc606_5 gpc535 (
      {stage0_13[118], stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[81],stage1_15[85],stage1_14[101],stage1_13[165]}
   );
   gpc606_5 gpc536 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[82],stage1_15[86],stage1_14[102],stage1_13[166]}
   );
   gpc606_5 gpc537 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[83],stage1_15[87],stage1_14[103],stage1_13[167]}
   );
   gpc606_5 gpc538 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[84],stage1_15[88],stage1_14[104],stage1_13[168]}
   );
   gpc606_5 gpc539 (
      {stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[85],stage1_15[89],stage1_14[105],stage1_13[169]}
   );
   gpc606_5 gpc540 (
      {stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[86],stage1_15[90],stage1_14[106],stage1_13[170]}
   );
   gpc606_5 gpc541 (
      {stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[87],stage1_15[91],stage1_14[107],stage1_13[171]}
   );
   gpc606_5 gpc542 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[88],stage1_15[92],stage1_14[108],stage1_13[172]}
   );
   gpc606_5 gpc543 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[89],stage1_15[93],stage1_14[109],stage1_13[173]}
   );
   gpc606_5 gpc544 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[90],stage1_15[94],stage1_14[110],stage1_13[174]}
   );
   gpc606_5 gpc545 (
      {stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[91],stage1_15[95],stage1_14[111],stage1_13[175]}
   );
   gpc606_5 gpc546 (
      {stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[92],stage1_15[96],stage1_14[112],stage1_13[176]}
   );
   gpc606_5 gpc547 (
      {stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[93],stage1_15[97],stage1_14[113],stage1_13[177]}
   );
   gpc606_5 gpc548 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[94],stage1_15[98],stage1_14[114],stage1_13[178]}
   );
   gpc606_5 gpc549 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[95],stage1_15[99],stage1_14[115],stage1_13[179]}
   );
   gpc606_5 gpc550 (
      {stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[96],stage1_15[100],stage1_14[116],stage1_13[180]}
   );
   gpc606_5 gpc551 (
      {stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[97],stage1_15[101],stage1_14[117],stage1_13[181]}
   );
   gpc606_5 gpc552 (
      {stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[98],stage1_15[102],stage1_14[118],stage1_13[182]}
   );
   gpc615_5 gpc553 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[422]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[99],stage1_15[103],stage1_14[119],stage1_13[183]}
   );
   gpc615_5 gpc554 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[423]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[100],stage1_15[104],stage1_14[120],stage1_13[184]}
   );
   gpc615_5 gpc555 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[424]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[101],stage1_15[105],stage1_14[121],stage1_13[185]}
   );
   gpc615_5 gpc556 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[425]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[102],stage1_15[106],stage1_14[122],stage1_13[186]}
   );
   gpc615_5 gpc557 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[426]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[103],stage1_15[107],stage1_14[123],stage1_13[187]}
   );
   gpc615_5 gpc558 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[427]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[104],stage1_15[108],stage1_14[124],stage1_13[188]}
   );
   gpc615_5 gpc559 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[428]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[105],stage1_15[109],stage1_14[125],stage1_13[189]}
   );
   gpc615_5 gpc560 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[429]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[106],stage1_15[110],stage1_14[126],stage1_13[190]}
   );
   gpc615_5 gpc561 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[430]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[107],stage1_15[111],stage1_14[127],stage1_13[191]}
   );
   gpc615_5 gpc562 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[431]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[108],stage1_15[112],stage1_14[128],stage1_13[192]}
   );
   gpc615_5 gpc563 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[432]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[109],stage1_15[113],stage1_14[129],stage1_13[193]}
   );
   gpc615_5 gpc564 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[433]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[110],stage1_15[114],stage1_14[130],stage1_13[194]}
   );
   gpc615_5 gpc565 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[434]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[111],stage1_15[115],stage1_14[131],stage1_13[195]}
   );
   gpc615_5 gpc566 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[435]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[112],stage1_15[116],stage1_14[132],stage1_13[196]}
   );
   gpc615_5 gpc567 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[436]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[113],stage1_15[117],stage1_14[133],stage1_13[197]}
   );
   gpc615_5 gpc568 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[437]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[114],stage1_15[118],stage1_14[134],stage1_13[198]}
   );
   gpc615_5 gpc569 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[438]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[115],stage1_15[119],stage1_14[135],stage1_13[199]}
   );
   gpc615_5 gpc570 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[439]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[116],stage1_15[120],stage1_14[136],stage1_13[200]}
   );
   gpc615_5 gpc571 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[440]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[117],stage1_15[121],stage1_14[137],stage1_13[201]}
   );
   gpc615_5 gpc572 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[441]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[118],stage1_15[122],stage1_14[138],stage1_13[202]}
   );
   gpc615_5 gpc573 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[442]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[119],stage1_15[123],stage1_14[139],stage1_13[203]}
   );
   gpc615_5 gpc574 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[443]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[120],stage1_15[124],stage1_14[140],stage1_13[204]}
   );
   gpc615_5 gpc575 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[444]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[121],stage1_15[125],stage1_14[141],stage1_13[205]}
   );
   gpc615_5 gpc576 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[445]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[122],stage1_15[126],stage1_14[142],stage1_13[206]}
   );
   gpc615_5 gpc577 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[446]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[123],stage1_15[127],stage1_14[143],stage1_13[207]}
   );
   gpc615_5 gpc578 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[447]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[124],stage1_15[128],stage1_14[144],stage1_13[208]}
   );
   gpc615_5 gpc579 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[448]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[125],stage1_15[129],stage1_14[145],stage1_13[209]}
   );
   gpc615_5 gpc580 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[449]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[126],stage1_15[130],stage1_14[146],stage1_13[210]}
   );
   gpc615_5 gpc581 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[450]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[127],stage1_15[131],stage1_14[147],stage1_13[211]}
   );
   gpc615_5 gpc582 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[451]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[128],stage1_15[132],stage1_14[148],stage1_13[212]}
   );
   gpc615_5 gpc583 (
      {stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_14[452]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[129],stage1_15[133],stage1_14[149],stage1_13[213]}
   );
   gpc615_5 gpc584 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385]},
      {stage0_14[453]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[130],stage1_15[134],stage1_14[150],stage1_13[214]}
   );
   gpc615_5 gpc585 (
      {stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390]},
      {stage0_14[454]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[131],stage1_15[135],stage1_14[151],stage1_13[215]}
   );
   gpc615_5 gpc586 (
      {stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_14[455]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[132],stage1_15[136],stage1_14[152],stage1_13[216]}
   );
   gpc615_5 gpc587 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400]},
      {stage0_14[456]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[133],stage1_15[137],stage1_14[153],stage1_13[217]}
   );
   gpc615_5 gpc588 (
      {stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405]},
      {stage0_14[457]},
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage1_17[64],stage1_16[134],stage1_15[138],stage1_14[154],stage1_13[218]}
   );
   gpc615_5 gpc589 (
      {stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_14[458]},
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage1_17[65],stage1_16[135],stage1_15[139],stage1_14[155],stage1_13[219]}
   );
   gpc615_5 gpc590 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415]},
      {stage0_14[459]},
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage1_17[66],stage1_16[136],stage1_15[140],stage1_14[156],stage1_13[220]}
   );
   gpc615_5 gpc591 (
      {stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420]},
      {stage0_14[460]},
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407]},
      {stage1_17[67],stage1_16[137],stage1_15[141],stage1_14[157],stage1_13[221]}
   );
   gpc615_5 gpc592 (
      {stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_14[461]},
      {stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage1_17[68],stage1_16[138],stage1_15[142],stage1_14[158],stage1_13[222]}
   );
   gpc615_5 gpc593 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430]},
      {stage0_14[462]},
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage1_17[69],stage1_16[139],stage1_15[143],stage1_14[159],stage1_13[223]}
   );
   gpc615_5 gpc594 (
      {stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435]},
      {stage0_14[463]},
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage1_17[70],stage1_16[140],stage1_15[144],stage1_14[160],stage1_13[224]}
   );
   gpc615_5 gpc595 (
      {stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_14[464]},
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage1_17[71],stage1_16[141],stage1_15[145],stage1_14[161],stage1_13[225]}
   );
   gpc615_5 gpc596 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445]},
      {stage0_14[465]},
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437]},
      {stage1_17[72],stage1_16[142],stage1_15[146],stage1_14[162],stage1_13[226]}
   );
   gpc615_5 gpc597 (
      {stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450]},
      {stage0_14[466]},
      {stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage1_17[73],stage1_16[143],stage1_15[147],stage1_14[163],stage1_13[227]}
   );
   gpc615_5 gpc598 (
      {stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_14[467]},
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage1_17[74],stage1_16[144],stage1_15[148],stage1_14[164],stage1_13[228]}
   );
   gpc615_5 gpc599 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[468]},
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage1_17[75],stage1_16[145],stage1_15[149],stage1_14[165],stage1_13[229]}
   );
   gpc615_5 gpc600 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[469]},
      {stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459], stage0_15[460], stage0_15[461]},
      {stage1_17[76],stage1_16[146],stage1_15[150],stage1_14[166],stage1_13[230]}
   );
   gpc615_5 gpc601 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[470]},
      {stage0_15[462], stage0_15[463], stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467]},
      {stage1_17[77],stage1_16[147],stage1_15[151],stage1_14[167],stage1_13[231]}
   );
   gpc615_5 gpc602 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[471]},
      {stage0_15[468], stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage1_17[78],stage1_16[148],stage1_15[152],stage1_14[168],stage1_13[232]}
   );
   gpc615_5 gpc603 (
      {stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480]},
      {stage0_14[472]},
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage1_17[79],stage1_16[149],stage1_15[153],stage1_14[169],stage1_13[233]}
   );
   gpc615_5 gpc604 (
      {stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_14[473]},
      {stage0_15[480], stage0_15[481], stage0_15[482], stage0_15[483], stage0_15[484], stage0_15[485]},
      {stage1_17[80],stage1_16[150],stage1_15[154],stage1_14[170],stage1_13[234]}
   );
   gpc1_1 gpc605 (
      {stage0_0[423]},
      {stage1_0[85]}
   );
   gpc1_1 gpc606 (
      {stage0_0[424]},
      {stage1_0[86]}
   );
   gpc1_1 gpc607 (
      {stage0_0[425]},
      {stage1_0[87]}
   );
   gpc1_1 gpc608 (
      {stage0_0[426]},
      {stage1_0[88]}
   );
   gpc1_1 gpc609 (
      {stage0_0[427]},
      {stage1_0[89]}
   );
   gpc1_1 gpc610 (
      {stage0_0[428]},
      {stage1_0[90]}
   );
   gpc1_1 gpc611 (
      {stage0_0[429]},
      {stage1_0[91]}
   );
   gpc1_1 gpc612 (
      {stage0_0[430]},
      {stage1_0[92]}
   );
   gpc1_1 gpc613 (
      {stage0_0[431]},
      {stage1_0[93]}
   );
   gpc1_1 gpc614 (
      {stage0_0[432]},
      {stage1_0[94]}
   );
   gpc1_1 gpc615 (
      {stage0_0[433]},
      {stage1_0[95]}
   );
   gpc1_1 gpc616 (
      {stage0_0[434]},
      {stage1_0[96]}
   );
   gpc1_1 gpc617 (
      {stage0_0[435]},
      {stage1_0[97]}
   );
   gpc1_1 gpc618 (
      {stage0_0[436]},
      {stage1_0[98]}
   );
   gpc1_1 gpc619 (
      {stage0_0[437]},
      {stage1_0[99]}
   );
   gpc1_1 gpc620 (
      {stage0_0[438]},
      {stage1_0[100]}
   );
   gpc1_1 gpc621 (
      {stage0_0[439]},
      {stage1_0[101]}
   );
   gpc1_1 gpc622 (
      {stage0_0[440]},
      {stage1_0[102]}
   );
   gpc1_1 gpc623 (
      {stage0_0[441]},
      {stage1_0[103]}
   );
   gpc1_1 gpc624 (
      {stage0_0[442]},
      {stage1_0[104]}
   );
   gpc1_1 gpc625 (
      {stage0_0[443]},
      {stage1_0[105]}
   );
   gpc1_1 gpc626 (
      {stage0_0[444]},
      {stage1_0[106]}
   );
   gpc1_1 gpc627 (
      {stage0_0[445]},
      {stage1_0[107]}
   );
   gpc1_1 gpc628 (
      {stage0_0[446]},
      {stage1_0[108]}
   );
   gpc1_1 gpc629 (
      {stage0_0[447]},
      {stage1_0[109]}
   );
   gpc1_1 gpc630 (
      {stage0_0[448]},
      {stage1_0[110]}
   );
   gpc1_1 gpc631 (
      {stage0_0[449]},
      {stage1_0[111]}
   );
   gpc1_1 gpc632 (
      {stage0_0[450]},
      {stage1_0[112]}
   );
   gpc1_1 gpc633 (
      {stage0_0[451]},
      {stage1_0[113]}
   );
   gpc1_1 gpc634 (
      {stage0_0[452]},
      {stage1_0[114]}
   );
   gpc1_1 gpc635 (
      {stage0_0[453]},
      {stage1_0[115]}
   );
   gpc1_1 gpc636 (
      {stage0_0[454]},
      {stage1_0[116]}
   );
   gpc1_1 gpc637 (
      {stage0_0[455]},
      {stage1_0[117]}
   );
   gpc1_1 gpc638 (
      {stage0_0[456]},
      {stage1_0[118]}
   );
   gpc1_1 gpc639 (
      {stage0_0[457]},
      {stage1_0[119]}
   );
   gpc1_1 gpc640 (
      {stage0_0[458]},
      {stage1_0[120]}
   );
   gpc1_1 gpc641 (
      {stage0_0[459]},
      {stage1_0[121]}
   );
   gpc1_1 gpc642 (
      {stage0_0[460]},
      {stage1_0[122]}
   );
   gpc1_1 gpc643 (
      {stage0_0[461]},
      {stage1_0[123]}
   );
   gpc1_1 gpc644 (
      {stage0_0[462]},
      {stage1_0[124]}
   );
   gpc1_1 gpc645 (
      {stage0_0[463]},
      {stage1_0[125]}
   );
   gpc1_1 gpc646 (
      {stage0_0[464]},
      {stage1_0[126]}
   );
   gpc1_1 gpc647 (
      {stage0_0[465]},
      {stage1_0[127]}
   );
   gpc1_1 gpc648 (
      {stage0_0[466]},
      {stage1_0[128]}
   );
   gpc1_1 gpc649 (
      {stage0_0[467]},
      {stage1_0[129]}
   );
   gpc1_1 gpc650 (
      {stage0_0[468]},
      {stage1_0[130]}
   );
   gpc1_1 gpc651 (
      {stage0_0[469]},
      {stage1_0[131]}
   );
   gpc1_1 gpc652 (
      {stage0_0[470]},
      {stage1_0[132]}
   );
   gpc1_1 gpc653 (
      {stage0_0[471]},
      {stage1_0[133]}
   );
   gpc1_1 gpc654 (
      {stage0_0[472]},
      {stage1_0[134]}
   );
   gpc1_1 gpc655 (
      {stage0_0[473]},
      {stage1_0[135]}
   );
   gpc1_1 gpc656 (
      {stage0_0[474]},
      {stage1_0[136]}
   );
   gpc1_1 gpc657 (
      {stage0_0[475]},
      {stage1_0[137]}
   );
   gpc1_1 gpc658 (
      {stage0_0[476]},
      {stage1_0[138]}
   );
   gpc1_1 gpc659 (
      {stage0_0[477]},
      {stage1_0[139]}
   );
   gpc1_1 gpc660 (
      {stage0_0[478]},
      {stage1_0[140]}
   );
   gpc1_1 gpc661 (
      {stage0_0[479]},
      {stage1_0[141]}
   );
   gpc1_1 gpc662 (
      {stage0_0[480]},
      {stage1_0[142]}
   );
   gpc1_1 gpc663 (
      {stage0_0[481]},
      {stage1_0[143]}
   );
   gpc1_1 gpc664 (
      {stage0_0[482]},
      {stage1_0[144]}
   );
   gpc1_1 gpc665 (
      {stage0_0[483]},
      {stage1_0[145]}
   );
   gpc1_1 gpc666 (
      {stage0_0[484]},
      {stage1_0[146]}
   );
   gpc1_1 gpc667 (
      {stage0_0[485]},
      {stage1_0[147]}
   );
   gpc1_1 gpc668 (
      {stage0_2[484]},
      {stage1_2[166]}
   );
   gpc1_1 gpc669 (
      {stage0_2[485]},
      {stage1_2[167]}
   );
   gpc1_1 gpc670 (
      {stage0_3[416]},
      {stage1_3[174]}
   );
   gpc1_1 gpc671 (
      {stage0_3[417]},
      {stage1_3[175]}
   );
   gpc1_1 gpc672 (
      {stage0_3[418]},
      {stage1_3[176]}
   );
   gpc1_1 gpc673 (
      {stage0_3[419]},
      {stage1_3[177]}
   );
   gpc1_1 gpc674 (
      {stage0_3[420]},
      {stage1_3[178]}
   );
   gpc1_1 gpc675 (
      {stage0_3[421]},
      {stage1_3[179]}
   );
   gpc1_1 gpc676 (
      {stage0_3[422]},
      {stage1_3[180]}
   );
   gpc1_1 gpc677 (
      {stage0_3[423]},
      {stage1_3[181]}
   );
   gpc1_1 gpc678 (
      {stage0_3[424]},
      {stage1_3[182]}
   );
   gpc1_1 gpc679 (
      {stage0_3[425]},
      {stage1_3[183]}
   );
   gpc1_1 gpc680 (
      {stage0_3[426]},
      {stage1_3[184]}
   );
   gpc1_1 gpc681 (
      {stage0_3[427]},
      {stage1_3[185]}
   );
   gpc1_1 gpc682 (
      {stage0_3[428]},
      {stage1_3[186]}
   );
   gpc1_1 gpc683 (
      {stage0_3[429]},
      {stage1_3[187]}
   );
   gpc1_1 gpc684 (
      {stage0_3[430]},
      {stage1_3[188]}
   );
   gpc1_1 gpc685 (
      {stage0_3[431]},
      {stage1_3[189]}
   );
   gpc1_1 gpc686 (
      {stage0_3[432]},
      {stage1_3[190]}
   );
   gpc1_1 gpc687 (
      {stage0_3[433]},
      {stage1_3[191]}
   );
   gpc1_1 gpc688 (
      {stage0_3[434]},
      {stage1_3[192]}
   );
   gpc1_1 gpc689 (
      {stage0_3[435]},
      {stage1_3[193]}
   );
   gpc1_1 gpc690 (
      {stage0_3[436]},
      {stage1_3[194]}
   );
   gpc1_1 gpc691 (
      {stage0_3[437]},
      {stage1_3[195]}
   );
   gpc1_1 gpc692 (
      {stage0_3[438]},
      {stage1_3[196]}
   );
   gpc1_1 gpc693 (
      {stage0_3[439]},
      {stage1_3[197]}
   );
   gpc1_1 gpc694 (
      {stage0_3[440]},
      {stage1_3[198]}
   );
   gpc1_1 gpc695 (
      {stage0_3[441]},
      {stage1_3[199]}
   );
   gpc1_1 gpc696 (
      {stage0_3[442]},
      {stage1_3[200]}
   );
   gpc1_1 gpc697 (
      {stage0_3[443]},
      {stage1_3[201]}
   );
   gpc1_1 gpc698 (
      {stage0_3[444]},
      {stage1_3[202]}
   );
   gpc1_1 gpc699 (
      {stage0_3[445]},
      {stage1_3[203]}
   );
   gpc1_1 gpc700 (
      {stage0_3[446]},
      {stage1_3[204]}
   );
   gpc1_1 gpc701 (
      {stage0_3[447]},
      {stage1_3[205]}
   );
   gpc1_1 gpc702 (
      {stage0_3[448]},
      {stage1_3[206]}
   );
   gpc1_1 gpc703 (
      {stage0_3[449]},
      {stage1_3[207]}
   );
   gpc1_1 gpc704 (
      {stage0_3[450]},
      {stage1_3[208]}
   );
   gpc1_1 gpc705 (
      {stage0_3[451]},
      {stage1_3[209]}
   );
   gpc1_1 gpc706 (
      {stage0_3[452]},
      {stage1_3[210]}
   );
   gpc1_1 gpc707 (
      {stage0_3[453]},
      {stage1_3[211]}
   );
   gpc1_1 gpc708 (
      {stage0_3[454]},
      {stage1_3[212]}
   );
   gpc1_1 gpc709 (
      {stage0_3[455]},
      {stage1_3[213]}
   );
   gpc1_1 gpc710 (
      {stage0_3[456]},
      {stage1_3[214]}
   );
   gpc1_1 gpc711 (
      {stage0_3[457]},
      {stage1_3[215]}
   );
   gpc1_1 gpc712 (
      {stage0_3[458]},
      {stage1_3[216]}
   );
   gpc1_1 gpc713 (
      {stage0_3[459]},
      {stage1_3[217]}
   );
   gpc1_1 gpc714 (
      {stage0_3[460]},
      {stage1_3[218]}
   );
   gpc1_1 gpc715 (
      {stage0_3[461]},
      {stage1_3[219]}
   );
   gpc1_1 gpc716 (
      {stage0_3[462]},
      {stage1_3[220]}
   );
   gpc1_1 gpc717 (
      {stage0_3[463]},
      {stage1_3[221]}
   );
   gpc1_1 gpc718 (
      {stage0_3[464]},
      {stage1_3[222]}
   );
   gpc1_1 gpc719 (
      {stage0_3[465]},
      {stage1_3[223]}
   );
   gpc1_1 gpc720 (
      {stage0_3[466]},
      {stage1_3[224]}
   );
   gpc1_1 gpc721 (
      {stage0_3[467]},
      {stage1_3[225]}
   );
   gpc1_1 gpc722 (
      {stage0_3[468]},
      {stage1_3[226]}
   );
   gpc1_1 gpc723 (
      {stage0_3[469]},
      {stage1_3[227]}
   );
   gpc1_1 gpc724 (
      {stage0_3[470]},
      {stage1_3[228]}
   );
   gpc1_1 gpc725 (
      {stage0_3[471]},
      {stage1_3[229]}
   );
   gpc1_1 gpc726 (
      {stage0_3[472]},
      {stage1_3[230]}
   );
   gpc1_1 gpc727 (
      {stage0_3[473]},
      {stage1_3[231]}
   );
   gpc1_1 gpc728 (
      {stage0_3[474]},
      {stage1_3[232]}
   );
   gpc1_1 gpc729 (
      {stage0_3[475]},
      {stage1_3[233]}
   );
   gpc1_1 gpc730 (
      {stage0_3[476]},
      {stage1_3[234]}
   );
   gpc1_1 gpc731 (
      {stage0_3[477]},
      {stage1_3[235]}
   );
   gpc1_1 gpc732 (
      {stage0_3[478]},
      {stage1_3[236]}
   );
   gpc1_1 gpc733 (
      {stage0_3[479]},
      {stage1_3[237]}
   );
   gpc1_1 gpc734 (
      {stage0_3[480]},
      {stage1_3[238]}
   );
   gpc1_1 gpc735 (
      {stage0_3[481]},
      {stage1_3[239]}
   );
   gpc1_1 gpc736 (
      {stage0_3[482]},
      {stage1_3[240]}
   );
   gpc1_1 gpc737 (
      {stage0_3[483]},
      {stage1_3[241]}
   );
   gpc1_1 gpc738 (
      {stage0_3[484]},
      {stage1_3[242]}
   );
   gpc1_1 gpc739 (
      {stage0_3[485]},
      {stage1_3[243]}
   );
   gpc1_1 gpc740 (
      {stage0_5[337]},
      {stage1_5[188]}
   );
   gpc1_1 gpc741 (
      {stage0_5[338]},
      {stage1_5[189]}
   );
   gpc1_1 gpc742 (
      {stage0_5[339]},
      {stage1_5[190]}
   );
   gpc1_1 gpc743 (
      {stage0_5[340]},
      {stage1_5[191]}
   );
   gpc1_1 gpc744 (
      {stage0_5[341]},
      {stage1_5[192]}
   );
   gpc1_1 gpc745 (
      {stage0_5[342]},
      {stage1_5[193]}
   );
   gpc1_1 gpc746 (
      {stage0_5[343]},
      {stage1_5[194]}
   );
   gpc1_1 gpc747 (
      {stage0_5[344]},
      {stage1_5[195]}
   );
   gpc1_1 gpc748 (
      {stage0_5[345]},
      {stage1_5[196]}
   );
   gpc1_1 gpc749 (
      {stage0_5[346]},
      {stage1_5[197]}
   );
   gpc1_1 gpc750 (
      {stage0_5[347]},
      {stage1_5[198]}
   );
   gpc1_1 gpc751 (
      {stage0_5[348]},
      {stage1_5[199]}
   );
   gpc1_1 gpc752 (
      {stage0_5[349]},
      {stage1_5[200]}
   );
   gpc1_1 gpc753 (
      {stage0_5[350]},
      {stage1_5[201]}
   );
   gpc1_1 gpc754 (
      {stage0_5[351]},
      {stage1_5[202]}
   );
   gpc1_1 gpc755 (
      {stage0_5[352]},
      {stage1_5[203]}
   );
   gpc1_1 gpc756 (
      {stage0_5[353]},
      {stage1_5[204]}
   );
   gpc1_1 gpc757 (
      {stage0_5[354]},
      {stage1_5[205]}
   );
   gpc1_1 gpc758 (
      {stage0_5[355]},
      {stage1_5[206]}
   );
   gpc1_1 gpc759 (
      {stage0_5[356]},
      {stage1_5[207]}
   );
   gpc1_1 gpc760 (
      {stage0_5[357]},
      {stage1_5[208]}
   );
   gpc1_1 gpc761 (
      {stage0_5[358]},
      {stage1_5[209]}
   );
   gpc1_1 gpc762 (
      {stage0_5[359]},
      {stage1_5[210]}
   );
   gpc1_1 gpc763 (
      {stage0_5[360]},
      {stage1_5[211]}
   );
   gpc1_1 gpc764 (
      {stage0_5[361]},
      {stage1_5[212]}
   );
   gpc1_1 gpc765 (
      {stage0_5[362]},
      {stage1_5[213]}
   );
   gpc1_1 gpc766 (
      {stage0_5[363]},
      {stage1_5[214]}
   );
   gpc1_1 gpc767 (
      {stage0_5[364]},
      {stage1_5[215]}
   );
   gpc1_1 gpc768 (
      {stage0_5[365]},
      {stage1_5[216]}
   );
   gpc1_1 gpc769 (
      {stage0_5[366]},
      {stage1_5[217]}
   );
   gpc1_1 gpc770 (
      {stage0_5[367]},
      {stage1_5[218]}
   );
   gpc1_1 gpc771 (
      {stage0_5[368]},
      {stage1_5[219]}
   );
   gpc1_1 gpc772 (
      {stage0_5[369]},
      {stage1_5[220]}
   );
   gpc1_1 gpc773 (
      {stage0_5[370]},
      {stage1_5[221]}
   );
   gpc1_1 gpc774 (
      {stage0_5[371]},
      {stage1_5[222]}
   );
   gpc1_1 gpc775 (
      {stage0_5[372]},
      {stage1_5[223]}
   );
   gpc1_1 gpc776 (
      {stage0_5[373]},
      {stage1_5[224]}
   );
   gpc1_1 gpc777 (
      {stage0_5[374]},
      {stage1_5[225]}
   );
   gpc1_1 gpc778 (
      {stage0_5[375]},
      {stage1_5[226]}
   );
   gpc1_1 gpc779 (
      {stage0_5[376]},
      {stage1_5[227]}
   );
   gpc1_1 gpc780 (
      {stage0_5[377]},
      {stage1_5[228]}
   );
   gpc1_1 gpc781 (
      {stage0_5[378]},
      {stage1_5[229]}
   );
   gpc1_1 gpc782 (
      {stage0_5[379]},
      {stage1_5[230]}
   );
   gpc1_1 gpc783 (
      {stage0_5[380]},
      {stage1_5[231]}
   );
   gpc1_1 gpc784 (
      {stage0_5[381]},
      {stage1_5[232]}
   );
   gpc1_1 gpc785 (
      {stage0_5[382]},
      {stage1_5[233]}
   );
   gpc1_1 gpc786 (
      {stage0_5[383]},
      {stage1_5[234]}
   );
   gpc1_1 gpc787 (
      {stage0_5[384]},
      {stage1_5[235]}
   );
   gpc1_1 gpc788 (
      {stage0_5[385]},
      {stage1_5[236]}
   );
   gpc1_1 gpc789 (
      {stage0_5[386]},
      {stage1_5[237]}
   );
   gpc1_1 gpc790 (
      {stage0_5[387]},
      {stage1_5[238]}
   );
   gpc1_1 gpc791 (
      {stage0_5[388]},
      {stage1_5[239]}
   );
   gpc1_1 gpc792 (
      {stage0_5[389]},
      {stage1_5[240]}
   );
   gpc1_1 gpc793 (
      {stage0_5[390]},
      {stage1_5[241]}
   );
   gpc1_1 gpc794 (
      {stage0_5[391]},
      {stage1_5[242]}
   );
   gpc1_1 gpc795 (
      {stage0_5[392]},
      {stage1_5[243]}
   );
   gpc1_1 gpc796 (
      {stage0_5[393]},
      {stage1_5[244]}
   );
   gpc1_1 gpc797 (
      {stage0_5[394]},
      {stage1_5[245]}
   );
   gpc1_1 gpc798 (
      {stage0_5[395]},
      {stage1_5[246]}
   );
   gpc1_1 gpc799 (
      {stage0_5[396]},
      {stage1_5[247]}
   );
   gpc1_1 gpc800 (
      {stage0_5[397]},
      {stage1_5[248]}
   );
   gpc1_1 gpc801 (
      {stage0_5[398]},
      {stage1_5[249]}
   );
   gpc1_1 gpc802 (
      {stage0_5[399]},
      {stage1_5[250]}
   );
   gpc1_1 gpc803 (
      {stage0_5[400]},
      {stage1_5[251]}
   );
   gpc1_1 gpc804 (
      {stage0_5[401]},
      {stage1_5[252]}
   );
   gpc1_1 gpc805 (
      {stage0_5[402]},
      {stage1_5[253]}
   );
   gpc1_1 gpc806 (
      {stage0_5[403]},
      {stage1_5[254]}
   );
   gpc1_1 gpc807 (
      {stage0_5[404]},
      {stage1_5[255]}
   );
   gpc1_1 gpc808 (
      {stage0_5[405]},
      {stage1_5[256]}
   );
   gpc1_1 gpc809 (
      {stage0_5[406]},
      {stage1_5[257]}
   );
   gpc1_1 gpc810 (
      {stage0_5[407]},
      {stage1_5[258]}
   );
   gpc1_1 gpc811 (
      {stage0_5[408]},
      {stage1_5[259]}
   );
   gpc1_1 gpc812 (
      {stage0_5[409]},
      {stage1_5[260]}
   );
   gpc1_1 gpc813 (
      {stage0_5[410]},
      {stage1_5[261]}
   );
   gpc1_1 gpc814 (
      {stage0_5[411]},
      {stage1_5[262]}
   );
   gpc1_1 gpc815 (
      {stage0_5[412]},
      {stage1_5[263]}
   );
   gpc1_1 gpc816 (
      {stage0_5[413]},
      {stage1_5[264]}
   );
   gpc1_1 gpc817 (
      {stage0_5[414]},
      {stage1_5[265]}
   );
   gpc1_1 gpc818 (
      {stage0_5[415]},
      {stage1_5[266]}
   );
   gpc1_1 gpc819 (
      {stage0_5[416]},
      {stage1_5[267]}
   );
   gpc1_1 gpc820 (
      {stage0_5[417]},
      {stage1_5[268]}
   );
   gpc1_1 gpc821 (
      {stage0_5[418]},
      {stage1_5[269]}
   );
   gpc1_1 gpc822 (
      {stage0_5[419]},
      {stage1_5[270]}
   );
   gpc1_1 gpc823 (
      {stage0_5[420]},
      {stage1_5[271]}
   );
   gpc1_1 gpc824 (
      {stage0_5[421]},
      {stage1_5[272]}
   );
   gpc1_1 gpc825 (
      {stage0_5[422]},
      {stage1_5[273]}
   );
   gpc1_1 gpc826 (
      {stage0_5[423]},
      {stage1_5[274]}
   );
   gpc1_1 gpc827 (
      {stage0_5[424]},
      {stage1_5[275]}
   );
   gpc1_1 gpc828 (
      {stage0_5[425]},
      {stage1_5[276]}
   );
   gpc1_1 gpc829 (
      {stage0_5[426]},
      {stage1_5[277]}
   );
   gpc1_1 gpc830 (
      {stage0_5[427]},
      {stage1_5[278]}
   );
   gpc1_1 gpc831 (
      {stage0_5[428]},
      {stage1_5[279]}
   );
   gpc1_1 gpc832 (
      {stage0_5[429]},
      {stage1_5[280]}
   );
   gpc1_1 gpc833 (
      {stage0_5[430]},
      {stage1_5[281]}
   );
   gpc1_1 gpc834 (
      {stage0_5[431]},
      {stage1_5[282]}
   );
   gpc1_1 gpc835 (
      {stage0_5[432]},
      {stage1_5[283]}
   );
   gpc1_1 gpc836 (
      {stage0_5[433]},
      {stage1_5[284]}
   );
   gpc1_1 gpc837 (
      {stage0_5[434]},
      {stage1_5[285]}
   );
   gpc1_1 gpc838 (
      {stage0_5[435]},
      {stage1_5[286]}
   );
   gpc1_1 gpc839 (
      {stage0_5[436]},
      {stage1_5[287]}
   );
   gpc1_1 gpc840 (
      {stage0_5[437]},
      {stage1_5[288]}
   );
   gpc1_1 gpc841 (
      {stage0_5[438]},
      {stage1_5[289]}
   );
   gpc1_1 gpc842 (
      {stage0_5[439]},
      {stage1_5[290]}
   );
   gpc1_1 gpc843 (
      {stage0_5[440]},
      {stage1_5[291]}
   );
   gpc1_1 gpc844 (
      {stage0_5[441]},
      {stage1_5[292]}
   );
   gpc1_1 gpc845 (
      {stage0_5[442]},
      {stage1_5[293]}
   );
   gpc1_1 gpc846 (
      {stage0_5[443]},
      {stage1_5[294]}
   );
   gpc1_1 gpc847 (
      {stage0_5[444]},
      {stage1_5[295]}
   );
   gpc1_1 gpc848 (
      {stage0_5[445]},
      {stage1_5[296]}
   );
   gpc1_1 gpc849 (
      {stage0_5[446]},
      {stage1_5[297]}
   );
   gpc1_1 gpc850 (
      {stage0_5[447]},
      {stage1_5[298]}
   );
   gpc1_1 gpc851 (
      {stage0_5[448]},
      {stage1_5[299]}
   );
   gpc1_1 gpc852 (
      {stage0_5[449]},
      {stage1_5[300]}
   );
   gpc1_1 gpc853 (
      {stage0_5[450]},
      {stage1_5[301]}
   );
   gpc1_1 gpc854 (
      {stage0_5[451]},
      {stage1_5[302]}
   );
   gpc1_1 gpc855 (
      {stage0_5[452]},
      {stage1_5[303]}
   );
   gpc1_1 gpc856 (
      {stage0_5[453]},
      {stage1_5[304]}
   );
   gpc1_1 gpc857 (
      {stage0_5[454]},
      {stage1_5[305]}
   );
   gpc1_1 gpc858 (
      {stage0_5[455]},
      {stage1_5[306]}
   );
   gpc1_1 gpc859 (
      {stage0_5[456]},
      {stage1_5[307]}
   );
   gpc1_1 gpc860 (
      {stage0_5[457]},
      {stage1_5[308]}
   );
   gpc1_1 gpc861 (
      {stage0_5[458]},
      {stage1_5[309]}
   );
   gpc1_1 gpc862 (
      {stage0_5[459]},
      {stage1_5[310]}
   );
   gpc1_1 gpc863 (
      {stage0_5[460]},
      {stage1_5[311]}
   );
   gpc1_1 gpc864 (
      {stage0_5[461]},
      {stage1_5[312]}
   );
   gpc1_1 gpc865 (
      {stage0_5[462]},
      {stage1_5[313]}
   );
   gpc1_1 gpc866 (
      {stage0_5[463]},
      {stage1_5[314]}
   );
   gpc1_1 gpc867 (
      {stage0_5[464]},
      {stage1_5[315]}
   );
   gpc1_1 gpc868 (
      {stage0_5[465]},
      {stage1_5[316]}
   );
   gpc1_1 gpc869 (
      {stage0_5[466]},
      {stage1_5[317]}
   );
   gpc1_1 gpc870 (
      {stage0_5[467]},
      {stage1_5[318]}
   );
   gpc1_1 gpc871 (
      {stage0_5[468]},
      {stage1_5[319]}
   );
   gpc1_1 gpc872 (
      {stage0_5[469]},
      {stage1_5[320]}
   );
   gpc1_1 gpc873 (
      {stage0_5[470]},
      {stage1_5[321]}
   );
   gpc1_1 gpc874 (
      {stage0_5[471]},
      {stage1_5[322]}
   );
   gpc1_1 gpc875 (
      {stage0_5[472]},
      {stage1_5[323]}
   );
   gpc1_1 gpc876 (
      {stage0_5[473]},
      {stage1_5[324]}
   );
   gpc1_1 gpc877 (
      {stage0_5[474]},
      {stage1_5[325]}
   );
   gpc1_1 gpc878 (
      {stage0_5[475]},
      {stage1_5[326]}
   );
   gpc1_1 gpc879 (
      {stage0_5[476]},
      {stage1_5[327]}
   );
   gpc1_1 gpc880 (
      {stage0_5[477]},
      {stage1_5[328]}
   );
   gpc1_1 gpc881 (
      {stage0_5[478]},
      {stage1_5[329]}
   );
   gpc1_1 gpc882 (
      {stage0_5[479]},
      {stage1_5[330]}
   );
   gpc1_1 gpc883 (
      {stage0_5[480]},
      {stage1_5[331]}
   );
   gpc1_1 gpc884 (
      {stage0_5[481]},
      {stage1_5[332]}
   );
   gpc1_1 gpc885 (
      {stage0_5[482]},
      {stage1_5[333]}
   );
   gpc1_1 gpc886 (
      {stage0_5[483]},
      {stage1_5[334]}
   );
   gpc1_1 gpc887 (
      {stage0_5[484]},
      {stage1_5[335]}
   );
   gpc1_1 gpc888 (
      {stage0_5[485]},
      {stage1_5[336]}
   );
   gpc1_1 gpc889 (
      {stage0_6[457]},
      {stage1_6[168]}
   );
   gpc1_1 gpc890 (
      {stage0_6[458]},
      {stage1_6[169]}
   );
   gpc1_1 gpc891 (
      {stage0_6[459]},
      {stage1_6[170]}
   );
   gpc1_1 gpc892 (
      {stage0_6[460]},
      {stage1_6[171]}
   );
   gpc1_1 gpc893 (
      {stage0_6[461]},
      {stage1_6[172]}
   );
   gpc1_1 gpc894 (
      {stage0_6[462]},
      {stage1_6[173]}
   );
   gpc1_1 gpc895 (
      {stage0_6[463]},
      {stage1_6[174]}
   );
   gpc1_1 gpc896 (
      {stage0_6[464]},
      {stage1_6[175]}
   );
   gpc1_1 gpc897 (
      {stage0_6[465]},
      {stage1_6[176]}
   );
   gpc1_1 gpc898 (
      {stage0_6[466]},
      {stage1_6[177]}
   );
   gpc1_1 gpc899 (
      {stage0_6[467]},
      {stage1_6[178]}
   );
   gpc1_1 gpc900 (
      {stage0_6[468]},
      {stage1_6[179]}
   );
   gpc1_1 gpc901 (
      {stage0_6[469]},
      {stage1_6[180]}
   );
   gpc1_1 gpc902 (
      {stage0_6[470]},
      {stage1_6[181]}
   );
   gpc1_1 gpc903 (
      {stage0_6[471]},
      {stage1_6[182]}
   );
   gpc1_1 gpc904 (
      {stage0_6[472]},
      {stage1_6[183]}
   );
   gpc1_1 gpc905 (
      {stage0_6[473]},
      {stage1_6[184]}
   );
   gpc1_1 gpc906 (
      {stage0_6[474]},
      {stage1_6[185]}
   );
   gpc1_1 gpc907 (
      {stage0_6[475]},
      {stage1_6[186]}
   );
   gpc1_1 gpc908 (
      {stage0_6[476]},
      {stage1_6[187]}
   );
   gpc1_1 gpc909 (
      {stage0_6[477]},
      {stage1_6[188]}
   );
   gpc1_1 gpc910 (
      {stage0_6[478]},
      {stage1_6[189]}
   );
   gpc1_1 gpc911 (
      {stage0_6[479]},
      {stage1_6[190]}
   );
   gpc1_1 gpc912 (
      {stage0_6[480]},
      {stage1_6[191]}
   );
   gpc1_1 gpc913 (
      {stage0_6[481]},
      {stage1_6[192]}
   );
   gpc1_1 gpc914 (
      {stage0_6[482]},
      {stage1_6[193]}
   );
   gpc1_1 gpc915 (
      {stage0_6[483]},
      {stage1_6[194]}
   );
   gpc1_1 gpc916 (
      {stage0_6[484]},
      {stage1_6[195]}
   );
   gpc1_1 gpc917 (
      {stage0_6[485]},
      {stage1_6[196]}
   );
   gpc1_1 gpc918 (
      {stage0_7[425]},
      {stage1_7[156]}
   );
   gpc1_1 gpc919 (
      {stage0_7[426]},
      {stage1_7[157]}
   );
   gpc1_1 gpc920 (
      {stage0_7[427]},
      {stage1_7[158]}
   );
   gpc1_1 gpc921 (
      {stage0_7[428]},
      {stage1_7[159]}
   );
   gpc1_1 gpc922 (
      {stage0_7[429]},
      {stage1_7[160]}
   );
   gpc1_1 gpc923 (
      {stage0_7[430]},
      {stage1_7[161]}
   );
   gpc1_1 gpc924 (
      {stage0_7[431]},
      {stage1_7[162]}
   );
   gpc1_1 gpc925 (
      {stage0_7[432]},
      {stage1_7[163]}
   );
   gpc1_1 gpc926 (
      {stage0_7[433]},
      {stage1_7[164]}
   );
   gpc1_1 gpc927 (
      {stage0_7[434]},
      {stage1_7[165]}
   );
   gpc1_1 gpc928 (
      {stage0_7[435]},
      {stage1_7[166]}
   );
   gpc1_1 gpc929 (
      {stage0_7[436]},
      {stage1_7[167]}
   );
   gpc1_1 gpc930 (
      {stage0_7[437]},
      {stage1_7[168]}
   );
   gpc1_1 gpc931 (
      {stage0_7[438]},
      {stage1_7[169]}
   );
   gpc1_1 gpc932 (
      {stage0_7[439]},
      {stage1_7[170]}
   );
   gpc1_1 gpc933 (
      {stage0_7[440]},
      {stage1_7[171]}
   );
   gpc1_1 gpc934 (
      {stage0_7[441]},
      {stage1_7[172]}
   );
   gpc1_1 gpc935 (
      {stage0_7[442]},
      {stage1_7[173]}
   );
   gpc1_1 gpc936 (
      {stage0_7[443]},
      {stage1_7[174]}
   );
   gpc1_1 gpc937 (
      {stage0_7[444]},
      {stage1_7[175]}
   );
   gpc1_1 gpc938 (
      {stage0_7[445]},
      {stage1_7[176]}
   );
   gpc1_1 gpc939 (
      {stage0_7[446]},
      {stage1_7[177]}
   );
   gpc1_1 gpc940 (
      {stage0_7[447]},
      {stage1_7[178]}
   );
   gpc1_1 gpc941 (
      {stage0_7[448]},
      {stage1_7[179]}
   );
   gpc1_1 gpc942 (
      {stage0_7[449]},
      {stage1_7[180]}
   );
   gpc1_1 gpc943 (
      {stage0_7[450]},
      {stage1_7[181]}
   );
   gpc1_1 gpc944 (
      {stage0_7[451]},
      {stage1_7[182]}
   );
   gpc1_1 gpc945 (
      {stage0_7[452]},
      {stage1_7[183]}
   );
   gpc1_1 gpc946 (
      {stage0_7[453]},
      {stage1_7[184]}
   );
   gpc1_1 gpc947 (
      {stage0_7[454]},
      {stage1_7[185]}
   );
   gpc1_1 gpc948 (
      {stage0_7[455]},
      {stage1_7[186]}
   );
   gpc1_1 gpc949 (
      {stage0_7[456]},
      {stage1_7[187]}
   );
   gpc1_1 gpc950 (
      {stage0_7[457]},
      {stage1_7[188]}
   );
   gpc1_1 gpc951 (
      {stage0_7[458]},
      {stage1_7[189]}
   );
   gpc1_1 gpc952 (
      {stage0_7[459]},
      {stage1_7[190]}
   );
   gpc1_1 gpc953 (
      {stage0_7[460]},
      {stage1_7[191]}
   );
   gpc1_1 gpc954 (
      {stage0_7[461]},
      {stage1_7[192]}
   );
   gpc1_1 gpc955 (
      {stage0_7[462]},
      {stage1_7[193]}
   );
   gpc1_1 gpc956 (
      {stage0_7[463]},
      {stage1_7[194]}
   );
   gpc1_1 gpc957 (
      {stage0_7[464]},
      {stage1_7[195]}
   );
   gpc1_1 gpc958 (
      {stage0_7[465]},
      {stage1_7[196]}
   );
   gpc1_1 gpc959 (
      {stage0_7[466]},
      {stage1_7[197]}
   );
   gpc1_1 gpc960 (
      {stage0_7[467]},
      {stage1_7[198]}
   );
   gpc1_1 gpc961 (
      {stage0_7[468]},
      {stage1_7[199]}
   );
   gpc1_1 gpc962 (
      {stage0_7[469]},
      {stage1_7[200]}
   );
   gpc1_1 gpc963 (
      {stage0_7[470]},
      {stage1_7[201]}
   );
   gpc1_1 gpc964 (
      {stage0_7[471]},
      {stage1_7[202]}
   );
   gpc1_1 gpc965 (
      {stage0_7[472]},
      {stage1_7[203]}
   );
   gpc1_1 gpc966 (
      {stage0_7[473]},
      {stage1_7[204]}
   );
   gpc1_1 gpc967 (
      {stage0_7[474]},
      {stage1_7[205]}
   );
   gpc1_1 gpc968 (
      {stage0_7[475]},
      {stage1_7[206]}
   );
   gpc1_1 gpc969 (
      {stage0_7[476]},
      {stage1_7[207]}
   );
   gpc1_1 gpc970 (
      {stage0_7[477]},
      {stage1_7[208]}
   );
   gpc1_1 gpc971 (
      {stage0_7[478]},
      {stage1_7[209]}
   );
   gpc1_1 gpc972 (
      {stage0_7[479]},
      {stage1_7[210]}
   );
   gpc1_1 gpc973 (
      {stage0_7[480]},
      {stage1_7[211]}
   );
   gpc1_1 gpc974 (
      {stage0_7[481]},
      {stage1_7[212]}
   );
   gpc1_1 gpc975 (
      {stage0_7[482]},
      {stage1_7[213]}
   );
   gpc1_1 gpc976 (
      {stage0_7[483]},
      {stage1_7[214]}
   );
   gpc1_1 gpc977 (
      {stage0_7[484]},
      {stage1_7[215]}
   );
   gpc1_1 gpc978 (
      {stage0_7[485]},
      {stage1_7[216]}
   );
   gpc1_1 gpc979 (
      {stage0_10[381]},
      {stage1_10[177]}
   );
   gpc1_1 gpc980 (
      {stage0_10[382]},
      {stage1_10[178]}
   );
   gpc1_1 gpc981 (
      {stage0_10[383]},
      {stage1_10[179]}
   );
   gpc1_1 gpc982 (
      {stage0_10[384]},
      {stage1_10[180]}
   );
   gpc1_1 gpc983 (
      {stage0_10[385]},
      {stage1_10[181]}
   );
   gpc1_1 gpc984 (
      {stage0_10[386]},
      {stage1_10[182]}
   );
   gpc1_1 gpc985 (
      {stage0_10[387]},
      {stage1_10[183]}
   );
   gpc1_1 gpc986 (
      {stage0_10[388]},
      {stage1_10[184]}
   );
   gpc1_1 gpc987 (
      {stage0_10[389]},
      {stage1_10[185]}
   );
   gpc1_1 gpc988 (
      {stage0_10[390]},
      {stage1_10[186]}
   );
   gpc1_1 gpc989 (
      {stage0_10[391]},
      {stage1_10[187]}
   );
   gpc1_1 gpc990 (
      {stage0_10[392]},
      {stage1_10[188]}
   );
   gpc1_1 gpc991 (
      {stage0_10[393]},
      {stage1_10[189]}
   );
   gpc1_1 gpc992 (
      {stage0_10[394]},
      {stage1_10[190]}
   );
   gpc1_1 gpc993 (
      {stage0_10[395]},
      {stage1_10[191]}
   );
   gpc1_1 gpc994 (
      {stage0_10[396]},
      {stage1_10[192]}
   );
   gpc1_1 gpc995 (
      {stage0_10[397]},
      {stage1_10[193]}
   );
   gpc1_1 gpc996 (
      {stage0_10[398]},
      {stage1_10[194]}
   );
   gpc1_1 gpc997 (
      {stage0_10[399]},
      {stage1_10[195]}
   );
   gpc1_1 gpc998 (
      {stage0_10[400]},
      {stage1_10[196]}
   );
   gpc1_1 gpc999 (
      {stage0_10[401]},
      {stage1_10[197]}
   );
   gpc1_1 gpc1000 (
      {stage0_10[402]},
      {stage1_10[198]}
   );
   gpc1_1 gpc1001 (
      {stage0_10[403]},
      {stage1_10[199]}
   );
   gpc1_1 gpc1002 (
      {stage0_10[404]},
      {stage1_10[200]}
   );
   gpc1_1 gpc1003 (
      {stage0_10[405]},
      {stage1_10[201]}
   );
   gpc1_1 gpc1004 (
      {stage0_10[406]},
      {stage1_10[202]}
   );
   gpc1_1 gpc1005 (
      {stage0_10[407]},
      {stage1_10[203]}
   );
   gpc1_1 gpc1006 (
      {stage0_10[408]},
      {stage1_10[204]}
   );
   gpc1_1 gpc1007 (
      {stage0_10[409]},
      {stage1_10[205]}
   );
   gpc1_1 gpc1008 (
      {stage0_10[410]},
      {stage1_10[206]}
   );
   gpc1_1 gpc1009 (
      {stage0_10[411]},
      {stage1_10[207]}
   );
   gpc1_1 gpc1010 (
      {stage0_10[412]},
      {stage1_10[208]}
   );
   gpc1_1 gpc1011 (
      {stage0_10[413]},
      {stage1_10[209]}
   );
   gpc1_1 gpc1012 (
      {stage0_10[414]},
      {stage1_10[210]}
   );
   gpc1_1 gpc1013 (
      {stage0_10[415]},
      {stage1_10[211]}
   );
   gpc1_1 gpc1014 (
      {stage0_10[416]},
      {stage1_10[212]}
   );
   gpc1_1 gpc1015 (
      {stage0_10[417]},
      {stage1_10[213]}
   );
   gpc1_1 gpc1016 (
      {stage0_10[418]},
      {stage1_10[214]}
   );
   gpc1_1 gpc1017 (
      {stage0_10[419]},
      {stage1_10[215]}
   );
   gpc1_1 gpc1018 (
      {stage0_10[420]},
      {stage1_10[216]}
   );
   gpc1_1 gpc1019 (
      {stage0_10[421]},
      {stage1_10[217]}
   );
   gpc1_1 gpc1020 (
      {stage0_10[422]},
      {stage1_10[218]}
   );
   gpc1_1 gpc1021 (
      {stage0_10[423]},
      {stage1_10[219]}
   );
   gpc1_1 gpc1022 (
      {stage0_10[424]},
      {stage1_10[220]}
   );
   gpc1_1 gpc1023 (
      {stage0_10[425]},
      {stage1_10[221]}
   );
   gpc1_1 gpc1024 (
      {stage0_10[426]},
      {stage1_10[222]}
   );
   gpc1_1 gpc1025 (
      {stage0_10[427]},
      {stage1_10[223]}
   );
   gpc1_1 gpc1026 (
      {stage0_10[428]},
      {stage1_10[224]}
   );
   gpc1_1 gpc1027 (
      {stage0_10[429]},
      {stage1_10[225]}
   );
   gpc1_1 gpc1028 (
      {stage0_10[430]},
      {stage1_10[226]}
   );
   gpc1_1 gpc1029 (
      {stage0_10[431]},
      {stage1_10[227]}
   );
   gpc1_1 gpc1030 (
      {stage0_10[432]},
      {stage1_10[228]}
   );
   gpc1_1 gpc1031 (
      {stage0_10[433]},
      {stage1_10[229]}
   );
   gpc1_1 gpc1032 (
      {stage0_10[434]},
      {stage1_10[230]}
   );
   gpc1_1 gpc1033 (
      {stage0_10[435]},
      {stage1_10[231]}
   );
   gpc1_1 gpc1034 (
      {stage0_10[436]},
      {stage1_10[232]}
   );
   gpc1_1 gpc1035 (
      {stage0_10[437]},
      {stage1_10[233]}
   );
   gpc1_1 gpc1036 (
      {stage0_10[438]},
      {stage1_10[234]}
   );
   gpc1_1 gpc1037 (
      {stage0_10[439]},
      {stage1_10[235]}
   );
   gpc1_1 gpc1038 (
      {stage0_10[440]},
      {stage1_10[236]}
   );
   gpc1_1 gpc1039 (
      {stage0_10[441]},
      {stage1_10[237]}
   );
   gpc1_1 gpc1040 (
      {stage0_10[442]},
      {stage1_10[238]}
   );
   gpc1_1 gpc1041 (
      {stage0_10[443]},
      {stage1_10[239]}
   );
   gpc1_1 gpc1042 (
      {stage0_10[444]},
      {stage1_10[240]}
   );
   gpc1_1 gpc1043 (
      {stage0_10[445]},
      {stage1_10[241]}
   );
   gpc1_1 gpc1044 (
      {stage0_10[446]},
      {stage1_10[242]}
   );
   gpc1_1 gpc1045 (
      {stage0_10[447]},
      {stage1_10[243]}
   );
   gpc1_1 gpc1046 (
      {stage0_10[448]},
      {stage1_10[244]}
   );
   gpc1_1 gpc1047 (
      {stage0_10[449]},
      {stage1_10[245]}
   );
   gpc1_1 gpc1048 (
      {stage0_10[450]},
      {stage1_10[246]}
   );
   gpc1_1 gpc1049 (
      {stage0_10[451]},
      {stage1_10[247]}
   );
   gpc1_1 gpc1050 (
      {stage0_10[452]},
      {stage1_10[248]}
   );
   gpc1_1 gpc1051 (
      {stage0_10[453]},
      {stage1_10[249]}
   );
   gpc1_1 gpc1052 (
      {stage0_10[454]},
      {stage1_10[250]}
   );
   gpc1_1 gpc1053 (
      {stage0_10[455]},
      {stage1_10[251]}
   );
   gpc1_1 gpc1054 (
      {stage0_10[456]},
      {stage1_10[252]}
   );
   gpc1_1 gpc1055 (
      {stage0_10[457]},
      {stage1_10[253]}
   );
   gpc1_1 gpc1056 (
      {stage0_10[458]},
      {stage1_10[254]}
   );
   gpc1_1 gpc1057 (
      {stage0_10[459]},
      {stage1_10[255]}
   );
   gpc1_1 gpc1058 (
      {stage0_10[460]},
      {stage1_10[256]}
   );
   gpc1_1 gpc1059 (
      {stage0_10[461]},
      {stage1_10[257]}
   );
   gpc1_1 gpc1060 (
      {stage0_10[462]},
      {stage1_10[258]}
   );
   gpc1_1 gpc1061 (
      {stage0_10[463]},
      {stage1_10[259]}
   );
   gpc1_1 gpc1062 (
      {stage0_10[464]},
      {stage1_10[260]}
   );
   gpc1_1 gpc1063 (
      {stage0_10[465]},
      {stage1_10[261]}
   );
   gpc1_1 gpc1064 (
      {stage0_10[466]},
      {stage1_10[262]}
   );
   gpc1_1 gpc1065 (
      {stage0_10[467]},
      {stage1_10[263]}
   );
   gpc1_1 gpc1066 (
      {stage0_10[468]},
      {stage1_10[264]}
   );
   gpc1_1 gpc1067 (
      {stage0_10[469]},
      {stage1_10[265]}
   );
   gpc1_1 gpc1068 (
      {stage0_10[470]},
      {stage1_10[266]}
   );
   gpc1_1 gpc1069 (
      {stage0_10[471]},
      {stage1_10[267]}
   );
   gpc1_1 gpc1070 (
      {stage0_10[472]},
      {stage1_10[268]}
   );
   gpc1_1 gpc1071 (
      {stage0_10[473]},
      {stage1_10[269]}
   );
   gpc1_1 gpc1072 (
      {stage0_10[474]},
      {stage1_10[270]}
   );
   gpc1_1 gpc1073 (
      {stage0_10[475]},
      {stage1_10[271]}
   );
   gpc1_1 gpc1074 (
      {stage0_10[476]},
      {stage1_10[272]}
   );
   gpc1_1 gpc1075 (
      {stage0_10[477]},
      {stage1_10[273]}
   );
   gpc1_1 gpc1076 (
      {stage0_10[478]},
      {stage1_10[274]}
   );
   gpc1_1 gpc1077 (
      {stage0_10[479]},
      {stage1_10[275]}
   );
   gpc1_1 gpc1078 (
      {stage0_10[480]},
      {stage1_10[276]}
   );
   gpc1_1 gpc1079 (
      {stage0_10[481]},
      {stage1_10[277]}
   );
   gpc1_1 gpc1080 (
      {stage0_10[482]},
      {stage1_10[278]}
   );
   gpc1_1 gpc1081 (
      {stage0_10[483]},
      {stage1_10[279]}
   );
   gpc1_1 gpc1082 (
      {stage0_10[484]},
      {stage1_10[280]}
   );
   gpc1_1 gpc1083 (
      {stage0_10[485]},
      {stage1_10[281]}
   );
   gpc1_1 gpc1084 (
      {stage0_11[423]},
      {stage1_11[151]}
   );
   gpc1_1 gpc1085 (
      {stage0_11[424]},
      {stage1_11[152]}
   );
   gpc1_1 gpc1086 (
      {stage0_11[425]},
      {stage1_11[153]}
   );
   gpc1_1 gpc1087 (
      {stage0_11[426]},
      {stage1_11[154]}
   );
   gpc1_1 gpc1088 (
      {stage0_11[427]},
      {stage1_11[155]}
   );
   gpc1_1 gpc1089 (
      {stage0_11[428]},
      {stage1_11[156]}
   );
   gpc1_1 gpc1090 (
      {stage0_11[429]},
      {stage1_11[157]}
   );
   gpc1_1 gpc1091 (
      {stage0_11[430]},
      {stage1_11[158]}
   );
   gpc1_1 gpc1092 (
      {stage0_11[431]},
      {stage1_11[159]}
   );
   gpc1_1 gpc1093 (
      {stage0_11[432]},
      {stage1_11[160]}
   );
   gpc1_1 gpc1094 (
      {stage0_11[433]},
      {stage1_11[161]}
   );
   gpc1_1 gpc1095 (
      {stage0_11[434]},
      {stage1_11[162]}
   );
   gpc1_1 gpc1096 (
      {stage0_11[435]},
      {stage1_11[163]}
   );
   gpc1_1 gpc1097 (
      {stage0_11[436]},
      {stage1_11[164]}
   );
   gpc1_1 gpc1098 (
      {stage0_11[437]},
      {stage1_11[165]}
   );
   gpc1_1 gpc1099 (
      {stage0_11[438]},
      {stage1_11[166]}
   );
   gpc1_1 gpc1100 (
      {stage0_11[439]},
      {stage1_11[167]}
   );
   gpc1_1 gpc1101 (
      {stage0_11[440]},
      {stage1_11[168]}
   );
   gpc1_1 gpc1102 (
      {stage0_11[441]},
      {stage1_11[169]}
   );
   gpc1_1 gpc1103 (
      {stage0_11[442]},
      {stage1_11[170]}
   );
   gpc1_1 gpc1104 (
      {stage0_11[443]},
      {stage1_11[171]}
   );
   gpc1_1 gpc1105 (
      {stage0_11[444]},
      {stage1_11[172]}
   );
   gpc1_1 gpc1106 (
      {stage0_11[445]},
      {stage1_11[173]}
   );
   gpc1_1 gpc1107 (
      {stage0_11[446]},
      {stage1_11[174]}
   );
   gpc1_1 gpc1108 (
      {stage0_11[447]},
      {stage1_11[175]}
   );
   gpc1_1 gpc1109 (
      {stage0_11[448]},
      {stage1_11[176]}
   );
   gpc1_1 gpc1110 (
      {stage0_11[449]},
      {stage1_11[177]}
   );
   gpc1_1 gpc1111 (
      {stage0_11[450]},
      {stage1_11[178]}
   );
   gpc1_1 gpc1112 (
      {stage0_11[451]},
      {stage1_11[179]}
   );
   gpc1_1 gpc1113 (
      {stage0_11[452]},
      {stage1_11[180]}
   );
   gpc1_1 gpc1114 (
      {stage0_11[453]},
      {stage1_11[181]}
   );
   gpc1_1 gpc1115 (
      {stage0_11[454]},
      {stage1_11[182]}
   );
   gpc1_1 gpc1116 (
      {stage0_11[455]},
      {stage1_11[183]}
   );
   gpc1_1 gpc1117 (
      {stage0_11[456]},
      {stage1_11[184]}
   );
   gpc1_1 gpc1118 (
      {stage0_11[457]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1119 (
      {stage0_11[458]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1120 (
      {stage0_11[459]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1121 (
      {stage0_11[460]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1122 (
      {stage0_11[461]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1123 (
      {stage0_11[462]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1124 (
      {stage0_11[463]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1125 (
      {stage0_11[464]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1126 (
      {stage0_11[465]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1127 (
      {stage0_11[466]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1128 (
      {stage0_11[467]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1129 (
      {stage0_11[468]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1130 (
      {stage0_11[469]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1131 (
      {stage0_11[470]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1132 (
      {stage0_11[471]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1133 (
      {stage0_11[472]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1134 (
      {stage0_11[473]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1135 (
      {stage0_11[474]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1136 (
      {stage0_11[475]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1137 (
      {stage0_11[476]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1138 (
      {stage0_11[477]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1139 (
      {stage0_11[478]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1140 (
      {stage0_11[479]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1141 (
      {stage0_11[480]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1142 (
      {stage0_11[481]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1143 (
      {stage0_11[482]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1144 (
      {stage0_11[483]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1145 (
      {stage0_11[484]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1146 (
      {stage0_11[485]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1147 (
      {stage0_14[474]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1148 (
      {stage0_14[475]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1149 (
      {stage0_14[476]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1150 (
      {stage0_14[477]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1151 (
      {stage0_14[478]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1152 (
      {stage0_14[479]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1153 (
      {stage0_14[480]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1154 (
      {stage0_14[481]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1155 (
      {stage0_14[482]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1156 (
      {stage0_14[483]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1157 (
      {stage0_14[484]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1158 (
      {stage0_14[485]},
      {stage1_14[182]}
   );
   gpc1163_5 gpc1159 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1160 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1161 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1162 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1163 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1164 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1165 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1166 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1167 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1168 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc1169 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc1170 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1171 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1172 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1173 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1174 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1175 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1176 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1177 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1178 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1179 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1180 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc1181 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1182 (
      {stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111], stage1_0[112], stage1_0[113]},
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc1183 (
      {stage1_0[114], stage1_0[115], stage1_0[116], stage1_0[117], stage1_0[118], stage1_0[119]},
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc606_5 gpc1184 (
      {stage1_0[120], stage1_0[121], stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125]},
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc606_5 gpc1185 (
      {stage1_0[126], stage1_0[127], stage1_0[128], stage1_0[129], stage1_0[130], stage1_0[131]},
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc1186 (
      {stage1_0[132], stage1_0[133], stage1_0[134], stage1_0[135], stage1_0[136], stage1_0[137]},
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27],stage2_0[27]}
   );
   gpc606_5 gpc1187 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage2_5[0],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1188 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[1],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1189 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[2],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1190 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[3],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1191 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[4],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1192 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[5],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1193 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[6],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1194 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[7],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc615_5 gpc1195 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[58]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[8],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc1196 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[59]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[9],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc1197 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[60]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[10],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc1198 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[11],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc1199 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[62]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[12],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc1200 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[63]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[13],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1201 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[64]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[14],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1202 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[15],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1203 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[16],stage2_4[44],stage2_3[44]}
   );
   gpc615_5 gpc1204 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[17],stage2_4[45],stage2_3[45]}
   );
   gpc615_5 gpc1205 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[18],stage2_4[46],stage2_3[46]}
   );
   gpc615_5 gpc1206 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[19],stage2_4[47],stage2_3[47]}
   );
   gpc615_5 gpc1207 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[20],stage2_4[48],stage2_3[48]}
   );
   gpc615_5 gpc1208 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[21],stage2_4[49],stage2_3[49]}
   );
   gpc615_5 gpc1209 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[22],stage2_4[50],stage2_3[50]}
   );
   gpc615_5 gpc1210 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[23],stage2_4[51],stage2_3[51]}
   );
   gpc615_5 gpc1211 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[56]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[16],stage2_5[24],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc1212 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[57]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[17],stage2_5[25],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc1213 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[58]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[18],stage2_5[26],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc1214 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[59]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[19],stage2_5[27],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc1215 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[60]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[20],stage2_5[28],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc1216 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[61]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[21],stage2_5[29],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc1217 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[62]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[22],stage2_5[30],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc1218 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[63]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[23],stage2_5[31],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc1219 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[64]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[24],stage2_5[32],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1220 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[65]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[25],stage2_5[33],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1221 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[66]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[26],stage2_5[34],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1222 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[67]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[27],stage2_5[35],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1223 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[68]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[28],stage2_5[36],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1224 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[69]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[29],stage2_5[37],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1225 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[70]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[30],stage2_5[38],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1226 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[71]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[31],stage2_5[39],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1227 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[72]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[32],stage2_5[40],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1228 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[73]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[33],stage2_5[41],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1229 (
      {stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199], stage1_3[200]},
      {stage1_4[74]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[34],stage2_5[42],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1230 (
      {stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204], stage1_3[205]},
      {stage1_4[75]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[35],stage2_5[43],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1231 (
      {stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209], stage1_3[210]},
      {stage1_4[76]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[36],stage2_5[44],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1232 (
      {stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214], stage1_3[215]},
      {stage1_4[77]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[37],stage2_5[45],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1233 (
      {stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219], stage1_3[220]},
      {stage1_4[78]},
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage2_7[30],stage2_6[38],stage2_5[46],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1234 (
      {stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224], stage1_3[225]},
      {stage1_4[79]},
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage2_7[31],stage2_6[39],stage2_5[47],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc1235 (
      {stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229], stage1_3[230]},
      {stage1_4[80]},
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage2_7[32],stage2_6[40],stage2_5[48],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc1236 (
      {stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234], stage1_3[235]},
      {stage1_4[81]},
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage2_7[33],stage2_6[41],stage2_5[49],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc1237 (
      {stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_5[204]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[34],stage2_6[42],stage2_5[50],stage2_4[78]}
   );
   gpc615_5 gpc1238 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_5[205]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[35],stage2_6[43],stage2_5[51],stage2_4[79]}
   );
   gpc615_5 gpc1239 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96]},
      {stage1_5[206]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[36],stage2_6[44],stage2_5[52],stage2_4[80]}
   );
   gpc615_5 gpc1240 (
      {stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_5[207]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[37],stage2_6[45],stage2_5[53],stage2_4[81]}
   );
   gpc615_5 gpc1241 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_5[208]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[38],stage2_6[46],stage2_5[54],stage2_4[82]}
   );
   gpc615_5 gpc1242 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111]},
      {stage1_5[209]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[39],stage2_6[47],stage2_5[55],stage2_4[83]}
   );
   gpc615_5 gpc1243 (
      {stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_5[210]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[40],stage2_6[48],stage2_5[56],stage2_4[84]}
   );
   gpc615_5 gpc1244 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_5[211]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[41],stage2_6[49],stage2_5[57],stage2_4[85]}
   );
   gpc615_5 gpc1245 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126]},
      {stage1_5[212]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[42],stage2_6[50],stage2_5[58],stage2_4[86]}
   );
   gpc615_5 gpc1246 (
      {stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage1_5[213]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[43],stage2_6[51],stage2_5[59],stage2_4[87]}
   );
   gpc615_5 gpc1247 (
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136]},
      {stage1_5[214]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[44],stage2_6[52],stage2_5[60],stage2_4[88]}
   );
   gpc615_5 gpc1248 (
      {stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_5[215]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[45],stage2_6[53],stage2_5[61],stage2_4[89]}
   );
   gpc615_5 gpc1249 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_5[216]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[46],stage2_6[54],stage2_5[62],stage2_4[90]}
   );
   gpc615_5 gpc1250 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151]},
      {stage1_5[217]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[47],stage2_6[55],stage2_5[63],stage2_4[91]}
   );
   gpc615_5 gpc1251 (
      {stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_5[218]},
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage2_8[14],stage2_7[48],stage2_6[56],stage2_5[64],stage2_4[92]}
   );
   gpc615_5 gpc1252 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage1_5[219]},
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage2_8[15],stage2_7[49],stage2_6[57],stage2_5[65],stage2_4[93]}
   );
   gpc615_5 gpc1253 (
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166]},
      {stage1_5[220]},
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage2_8[16],stage2_7[50],stage2_6[58],stage2_5[66],stage2_4[94]}
   );
   gpc615_5 gpc1254 (
      {stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_5[221]},
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage2_8[17],stage2_7[51],stage2_6[59],stage2_5[67],stage2_4[95]}
   );
   gpc615_5 gpc1255 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_5[222]},
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage2_8[18],stage2_7[52],stage2_6[60],stage2_5[68],stage2_4[96]}
   );
   gpc615_5 gpc1256 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181]},
      {stage1_5[223]},
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage2_8[19],stage2_7[53],stage2_6[61],stage2_5[69],stage2_4[97]}
   );
   gpc615_5 gpc1257 (
      {stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_5[224]},
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage2_8[20],stage2_7[54],stage2_6[62],stage2_5[70],stage2_4[98]}
   );
   gpc615_5 gpc1258 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191]},
      {stage1_5[225]},
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage2_8[21],stage2_7[55],stage2_6[63],stage2_5[71],stage2_4[99]}
   );
   gpc615_5 gpc1259 (
      {stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196]},
      {stage1_5[226]},
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage2_8[22],stage2_7[56],stage2_6[64],stage2_5[72],stage2_4[100]}
   );
   gpc615_5 gpc1260 (
      {stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_5[227]},
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage2_8[23],stage2_7[57],stage2_6[65],stage2_5[73],stage2_4[101]}
   );
   gpc615_5 gpc1261 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_5[228]},
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage2_8[24],stage2_7[58],stage2_6[66],stage2_5[74],stage2_4[102]}
   );
   gpc615_5 gpc1262 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[229]},
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage2_8[25],stage2_7[59],stage2_6[67],stage2_5[75],stage2_4[103]}
   );
   gpc615_5 gpc1263 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[230]},
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage2_8[26],stage2_7[60],stage2_6[68],stage2_5[76],stage2_4[104]}
   );
   gpc615_5 gpc1264 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_5[231]},
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage2_8[27],stage2_7[61],stage2_6[69],stage2_5[77],stage2_4[105]}
   );
   gpc606_5 gpc1265 (
      {stage1_5[232], stage1_5[233], stage1_5[234], stage1_5[235], stage1_5[236], stage1_5[237]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[28],stage2_7[62],stage2_6[70],stage2_5[78]}
   );
   gpc606_5 gpc1266 (
      {stage1_5[238], stage1_5[239], stage1_5[240], stage1_5[241], stage1_5[242], stage1_5[243]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[29],stage2_7[63],stage2_6[71],stage2_5[79]}
   );
   gpc606_5 gpc1267 (
      {stage1_5[244], stage1_5[245], stage1_5[246], stage1_5[247], stage1_5[248], stage1_5[249]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[30],stage2_7[64],stage2_6[72],stage2_5[80]}
   );
   gpc606_5 gpc1268 (
      {stage1_5[250], stage1_5[251], stage1_5[252], stage1_5[253], stage1_5[254], stage1_5[255]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[31],stage2_7[65],stage2_6[73],stage2_5[81]}
   );
   gpc606_5 gpc1269 (
      {stage1_5[256], stage1_5[257], stage1_5[258], stage1_5[259], stage1_5[260], stage1_5[261]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[32],stage2_7[66],stage2_6[74],stage2_5[82]}
   );
   gpc606_5 gpc1270 (
      {stage1_5[262], stage1_5[263], stage1_5[264], stage1_5[265], stage1_5[266], stage1_5[267]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[33],stage2_7[67],stage2_6[75],stage2_5[83]}
   );
   gpc606_5 gpc1271 (
      {stage1_5[268], stage1_5[269], stage1_5[270], stage1_5[271], stage1_5[272], stage1_5[273]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[34],stage2_7[68],stage2_6[76],stage2_5[84]}
   );
   gpc606_5 gpc1272 (
      {stage1_5[274], stage1_5[275], stage1_5[276], stage1_5[277], stage1_5[278], stage1_5[279]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[35],stage2_7[69],stage2_6[77],stage2_5[85]}
   );
   gpc606_5 gpc1273 (
      {stage1_5[280], stage1_5[281], stage1_5[282], stage1_5[283], stage1_5[284], stage1_5[285]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[36],stage2_7[70],stage2_6[78],stage2_5[86]}
   );
   gpc606_5 gpc1274 (
      {stage1_5[286], stage1_5[287], stage1_5[288], stage1_5[289], stage1_5[290], stage1_5[291]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[37],stage2_7[71],stage2_6[79],stage2_5[87]}
   );
   gpc606_5 gpc1275 (
      {stage1_5[292], stage1_5[293], stage1_5[294], stage1_5[295], stage1_5[296], stage1_5[297]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[38],stage2_7[72],stage2_6[80],stage2_5[88]}
   );
   gpc606_5 gpc1276 (
      {stage1_5[298], stage1_5[299], stage1_5[300], stage1_5[301], stage1_5[302], stage1_5[303]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[39],stage2_7[73],stage2_6[81],stage2_5[89]}
   );
   gpc606_5 gpc1277 (
      {stage1_5[304], stage1_5[305], stage1_5[306], stage1_5[307], stage1_5[308], stage1_5[309]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[40],stage2_7[74],stage2_6[82],stage2_5[90]}
   );
   gpc606_5 gpc1278 (
      {stage1_5[310], stage1_5[311], stage1_5[312], stage1_5[313], stage1_5[314], stage1_5[315]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[41],stage2_7[75],stage2_6[83],stage2_5[91]}
   );
   gpc606_5 gpc1279 (
      {stage1_5[316], stage1_5[317], stage1_5[318], stage1_5[319], stage1_5[320], stage1_5[321]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[42],stage2_7[76],stage2_6[84],stage2_5[92]}
   );
   gpc606_5 gpc1280 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[43],stage2_7[77],stage2_6[85]}
   );
   gpc606_5 gpc1281 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[44],stage2_7[78],stage2_6[86]}
   );
   gpc606_5 gpc1282 (
      {stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[45],stage2_7[79],stage2_6[87]}
   );
   gpc606_5 gpc1283 (
      {stage1_6[186], stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[46],stage2_7[80],stage2_6[88]}
   );
   gpc615_5 gpc1284 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[90]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[47],stage2_7[81],stage2_6[89]}
   );
   gpc606_5 gpc1285 (
      {stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[20],stage2_8[48],stage2_7[82]}
   );
   gpc606_5 gpc1286 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[21],stage2_8[49],stage2_7[83]}
   );
   gpc606_5 gpc1287 (
      {stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[22],stage2_8[50],stage2_7[84]}
   );
   gpc606_5 gpc1288 (
      {stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[23],stage2_8[51],stage2_7[85]}
   );
   gpc606_5 gpc1289 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[24],stage2_8[52],stage2_7[86]}
   );
   gpc606_5 gpc1290 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[25],stage2_8[53],stage2_7[87]}
   );
   gpc606_5 gpc1291 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131], stage1_7[132]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[26],stage2_8[54],stage2_7[88]}
   );
   gpc606_5 gpc1292 (
      {stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[27],stage2_8[55],stage2_7[89]}
   );
   gpc606_5 gpc1293 (
      {stage1_7[139], stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[28],stage2_8[56],stage2_7[90]}
   );
   gpc606_5 gpc1294 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[29],stage2_8[57],stage2_7[91]}
   );
   gpc606_5 gpc1295 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[30],stage2_8[58],stage2_7[92]}
   );
   gpc606_5 gpc1296 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161], stage1_7[162]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[31],stage2_8[59],stage2_7[93]}
   );
   gpc606_5 gpc1297 (
      {stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[32],stage2_8[60],stage2_7[94]}
   );
   gpc606_5 gpc1298 (
      {stage1_7[169], stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[33],stage2_8[61],stage2_7[95]}
   );
   gpc606_5 gpc1299 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[34],stage2_8[62],stage2_7[96]}
   );
   gpc606_5 gpc1300 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[35],stage2_8[63],stage2_7[97]}
   );
   gpc606_5 gpc1301 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191], stage1_7[192]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[36],stage2_8[64],stage2_7[98]}
   );
   gpc606_5 gpc1302 (
      {stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[37],stage2_8[65],stage2_7[99]}
   );
   gpc606_5 gpc1303 (
      {stage1_7[199], stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[38],stage2_8[66],stage2_7[100]}
   );
   gpc606_5 gpc1304 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[39],stage2_8[67],stage2_7[101]}
   );
   gpc606_5 gpc1305 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[40],stage2_8[68],stage2_7[102]}
   );
   gpc606_5 gpc1306 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[21],stage2_10[26],stage2_9[41],stage2_8[69]}
   );
   gpc606_5 gpc1307 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[22],stage2_10[27],stage2_9[42],stage2_8[70]}
   );
   gpc606_5 gpc1308 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[23],stage2_10[28],stage2_9[43],stage2_8[71]}
   );
   gpc606_5 gpc1309 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[24],stage2_10[29],stage2_9[44],stage2_8[72]}
   );
   gpc606_5 gpc1310 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[25],stage2_10[30],stage2_9[45],stage2_8[73]}
   );
   gpc606_5 gpc1311 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[26],stage2_10[31],stage2_9[46],stage2_8[74]}
   );
   gpc606_5 gpc1312 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[27],stage2_10[32],stage2_9[47],stage2_8[75]}
   );
   gpc606_5 gpc1313 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[28],stage2_10[33],stage2_9[48],stage2_8[76]}
   );
   gpc606_5 gpc1314 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[29],stage2_10[34],stage2_9[49],stage2_8[77]}
   );
   gpc606_5 gpc1315 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[30],stage2_10[35],stage2_9[50],stage2_8[78]}
   );
   gpc606_5 gpc1316 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[31],stage2_10[36],stage2_9[51],stage2_8[79]}
   );
   gpc606_5 gpc1317 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[32],stage2_10[37],stage2_9[52],stage2_8[80]}
   );
   gpc606_5 gpc1318 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[33],stage2_10[38],stage2_9[53],stage2_8[81]}
   );
   gpc606_5 gpc1319 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[34],stage2_10[39],stage2_9[54],stage2_8[82]}
   );
   gpc606_5 gpc1320 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[35],stage2_10[40],stage2_9[55],stage2_8[83]}
   );
   gpc606_5 gpc1321 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[36],stage2_10[41],stage2_9[56],stage2_8[84]}
   );
   gpc606_5 gpc1322 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[37],stage2_10[42],stage2_9[57],stage2_8[85]}
   );
   gpc606_5 gpc1323 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[38],stage2_10[43],stage2_9[58],stage2_8[86]}
   );
   gpc606_5 gpc1324 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[39],stage2_10[44],stage2_9[59],stage2_8[87]}
   );
   gpc606_5 gpc1325 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[40],stage2_10[45],stage2_9[60],stage2_8[88]}
   );
   gpc606_5 gpc1326 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[41],stage2_10[46],stage2_9[61],stage2_8[89]}
   );
   gpc606_5 gpc1327 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[42],stage2_10[47],stage2_9[62],stage2_8[90]}
   );
   gpc606_5 gpc1328 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[43],stage2_10[48],stage2_9[63],stage2_8[91]}
   );
   gpc606_5 gpc1329 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[44],stage2_10[49],stage2_9[64],stage2_8[92]}
   );
   gpc606_5 gpc1330 (
      {stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177], stage1_8[178], stage1_8[179]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[45],stage2_10[50],stage2_9[65],stage2_8[93]}
   );
   gpc615_5 gpc1331 (
      {stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183], stage1_8[184]},
      {stage1_9[126]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[46],stage2_10[51],stage2_9[66],stage2_8[94]}
   );
   gpc606_5 gpc1332 (
      {stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131], stage1_9[132]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[26],stage2_11[47],stage2_10[52],stage2_9[67]}
   );
   gpc606_5 gpc1333 (
      {stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137], stage1_9[138]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[27],stage2_11[48],stage2_10[53],stage2_9[68]}
   );
   gpc606_5 gpc1334 (
      {stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143], stage1_9[144]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[28],stage2_11[49],stage2_10[54],stage2_9[69]}
   );
   gpc606_5 gpc1335 (
      {stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149], stage1_9[150]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[29],stage2_11[50],stage2_10[55],stage2_9[70]}
   );
   gpc606_5 gpc1336 (
      {stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155], stage1_9[156]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[30],stage2_11[51],stage2_10[56],stage2_9[71]}
   );
   gpc606_5 gpc1337 (
      {stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161], stage1_9[162]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[31],stage2_11[52],stage2_10[57],stage2_9[72]}
   );
   gpc606_5 gpc1338 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[32],stage2_11[53],stage2_10[58],stage2_9[73]}
   );
   gpc606_5 gpc1339 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[33],stage2_11[54],stage2_10[59],stage2_9[74]}
   );
   gpc606_5 gpc1340 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[34],stage2_11[55],stage2_10[60],stage2_9[75]}
   );
   gpc606_5 gpc1341 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185], stage1_9[186]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[35],stage2_11[56],stage2_10[61],stage2_9[76]}
   );
   gpc606_5 gpc1342 (
      {stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[36],stage2_11[57],stage2_10[62],stage2_9[77]}
   );
   gpc606_5 gpc1343 (
      {stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[37],stage2_11[58],stage2_10[63],stage2_9[78]}
   );
   gpc606_5 gpc1344 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[38],stage2_11[59],stage2_10[64],stage2_9[79]}
   );
   gpc606_5 gpc1345 (
      {stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[39],stage2_11[60],stage2_10[65],stage2_9[80]}
   );
   gpc606_5 gpc1346 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[14],stage2_12[40],stage2_11[61],stage2_10[66]}
   );
   gpc606_5 gpc1347 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[15],stage2_12[41],stage2_11[62],stage2_10[67]}
   );
   gpc606_5 gpc1348 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[16],stage2_12[42],stage2_11[63],stage2_10[68]}
   );
   gpc606_5 gpc1349 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[17],stage2_12[43],stage2_11[64],stage2_10[69]}
   );
   gpc606_5 gpc1350 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[18],stage2_12[44],stage2_11[65],stage2_10[70]}
   );
   gpc606_5 gpc1351 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[19],stage2_12[45],stage2_11[66],stage2_10[71]}
   );
   gpc606_5 gpc1352 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[20],stage2_12[46],stage2_11[67],stage2_10[72]}
   );
   gpc606_5 gpc1353 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[21],stage2_12[47],stage2_11[68],stage2_10[73]}
   );
   gpc606_5 gpc1354 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[22],stage2_12[48],stage2_11[69],stage2_10[74]}
   );
   gpc606_5 gpc1355 (
      {stage1_10[210], stage1_10[211], stage1_10[212], stage1_10[213], stage1_10[214], stage1_10[215]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[23],stage2_12[49],stage2_11[70],stage2_10[75]}
   );
   gpc615_5 gpc1356 (
      {stage1_10[216], stage1_10[217], stage1_10[218], stage1_10[219], stage1_10[220]},
      {stage1_11[84]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[24],stage2_12[50],stage2_11[71],stage2_10[76]}
   );
   gpc615_5 gpc1357 (
      {stage1_10[221], stage1_10[222], stage1_10[223], stage1_10[224], stage1_10[225]},
      {stage1_11[85]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[25],stage2_12[51],stage2_11[72],stage2_10[77]}
   );
   gpc615_5 gpc1358 (
      {stage1_10[226], stage1_10[227], stage1_10[228], stage1_10[229], stage1_10[230]},
      {stage1_11[86]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[26],stage2_12[52],stage2_11[73],stage2_10[78]}
   );
   gpc615_5 gpc1359 (
      {stage1_10[231], stage1_10[232], stage1_10[233], stage1_10[234], stage1_10[235]},
      {stage1_11[87]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[27],stage2_12[53],stage2_11[74],stage2_10[79]}
   );
   gpc615_5 gpc1360 (
      {stage1_10[236], stage1_10[237], stage1_10[238], stage1_10[239], stage1_10[240]},
      {stage1_11[88]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[28],stage2_12[54],stage2_11[75],stage2_10[80]}
   );
   gpc615_5 gpc1361 (
      {stage1_10[241], stage1_10[242], stage1_10[243], stage1_10[244], stage1_10[245]},
      {stage1_11[89]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[29],stage2_12[55],stage2_11[76],stage2_10[81]}
   );
   gpc615_5 gpc1362 (
      {stage1_10[246], stage1_10[247], stage1_10[248], stage1_10[249], stage1_10[250]},
      {stage1_11[90]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[30],stage2_12[56],stage2_11[77],stage2_10[82]}
   );
   gpc615_5 gpc1363 (
      {stage1_10[251], stage1_10[252], stage1_10[253], stage1_10[254], stage1_10[255]},
      {stage1_11[91]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage2_14[17],stage2_13[31],stage2_12[57],stage2_11[78],stage2_10[83]}
   );
   gpc615_5 gpc1364 (
      {stage1_10[256], stage1_10[257], stage1_10[258], stage1_10[259], stage1_10[260]},
      {stage1_11[92]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage2_14[18],stage2_13[32],stage2_12[58],stage2_11[79],stage2_10[84]}
   );
   gpc615_5 gpc1365 (
      {stage1_10[261], stage1_10[262], stage1_10[263], stage1_10[264], stage1_10[265]},
      {stage1_11[93]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage2_14[19],stage2_13[33],stage2_12[59],stage2_11[80],stage2_10[85]}
   );
   gpc615_5 gpc1366 (
      {stage1_10[266], stage1_10[267], stage1_10[268], stage1_10[269], stage1_10[270]},
      {stage1_11[94]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage2_14[20],stage2_13[34],stage2_12[60],stage2_11[81],stage2_10[86]}
   );
   gpc615_5 gpc1367 (
      {stage1_10[271], stage1_10[272], stage1_10[273], stage1_10[274], stage1_10[275]},
      {stage1_11[95]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage2_14[21],stage2_13[35],stage2_12[61],stage2_11[82],stage2_10[87]}
   );
   gpc615_5 gpc1368 (
      {stage1_10[276], stage1_10[277], stage1_10[278], stage1_10[279], stage1_10[280]},
      {stage1_11[96]},
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage2_14[22],stage2_13[36],stage2_12[62],stage2_11[83],stage2_10[88]}
   );
   gpc606_5 gpc1369 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[23],stage2_13[37],stage2_12[63],stage2_11[84]}
   );
   gpc606_5 gpc1370 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[24],stage2_13[38],stage2_12[64],stage2_11[85]}
   );
   gpc615_5 gpc1371 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage1_12[138]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[25],stage2_13[39],stage2_12[65],stage2_11[86]}
   );
   gpc615_5 gpc1372 (
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118]},
      {stage1_12[139]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[26],stage2_13[40],stage2_12[66],stage2_11[87]}
   );
   gpc615_5 gpc1373 (
      {stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[140]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[27],stage2_13[41],stage2_12[67],stage2_11[88]}
   );
   gpc615_5 gpc1374 (
      {stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128]},
      {stage1_12[141]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[28],stage2_13[42],stage2_12[68],stage2_11[89]}
   );
   gpc615_5 gpc1375 (
      {stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133]},
      {stage1_12[142]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[29],stage2_13[43],stage2_12[69],stage2_11[90]}
   );
   gpc615_5 gpc1376 (
      {stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[143]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[30],stage2_13[44],stage2_12[70],stage2_11[91]}
   );
   gpc615_5 gpc1377 (
      {stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143]},
      {stage1_12[144]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[31],stage2_13[45],stage2_12[71],stage2_11[92]}
   );
   gpc615_5 gpc1378 (
      {stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148]},
      {stage1_12[145]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[32],stage2_13[46],stage2_12[72],stage2_11[93]}
   );
   gpc615_5 gpc1379 (
      {stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[146]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[33],stage2_13[47],stage2_12[73],stage2_11[94]}
   );
   gpc615_5 gpc1380 (
      {stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158]},
      {stage1_12[147]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[34],stage2_13[48],stage2_12[74],stage2_11[95]}
   );
   gpc615_5 gpc1381 (
      {stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163]},
      {stage1_12[148]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[35],stage2_13[49],stage2_12[75],stage2_11[96]}
   );
   gpc615_5 gpc1382 (
      {stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[149]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[36],stage2_13[50],stage2_12[76],stage2_11[97]}
   );
   gpc615_5 gpc1383 (
      {stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173]},
      {stage1_12[150]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[37],stage2_13[51],stage2_12[77],stage2_11[98]}
   );
   gpc615_5 gpc1384 (
      {stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178]},
      {stage1_12[151]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[38],stage2_13[52],stage2_12[78],stage2_11[99]}
   );
   gpc615_5 gpc1385 (
      {stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183]},
      {stage1_12[152]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[39],stage2_13[53],stage2_12[79],stage2_11[100]}
   );
   gpc615_5 gpc1386 (
      {stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188]},
      {stage1_12[153]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[40],stage2_13[54],stage2_12[80],stage2_11[101]}
   );
   gpc615_5 gpc1387 (
      {stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193]},
      {stage1_12[154]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[41],stage2_13[55],stage2_12[81],stage2_11[102]}
   );
   gpc615_5 gpc1388 (
      {stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198]},
      {stage1_12[155]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[42],stage2_13[56],stage2_12[82],stage2_11[103]}
   );
   gpc615_5 gpc1389 (
      {stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203]},
      {stage1_12[156]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[43],stage2_13[57],stage2_12[83],stage2_11[104]}
   );
   gpc615_5 gpc1390 (
      {stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208]},
      {stage1_12[157]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[44],stage2_13[58],stage2_12[84],stage2_11[105]}
   );
   gpc615_5 gpc1391 (
      {stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213]},
      {stage1_12[158]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[45],stage2_13[59],stage2_12[85],stage2_11[106]}
   );
   gpc606_5 gpc1392 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[23],stage2_14[46],stage2_13[60],stage2_12[86]}
   );
   gpc606_5 gpc1393 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[24],stage2_14[47],stage2_13[61],stage2_12[87]}
   );
   gpc606_5 gpc1394 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[25],stage2_14[48],stage2_13[62],stage2_12[88]}
   );
   gpc606_5 gpc1395 (
      {stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180], stage1_12[181], stage1_12[182]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[26],stage2_14[49],stage2_13[63],stage2_12[89]}
   );
   gpc606_5 gpc1396 (
      {stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[27],stage2_14[50],stage2_13[64],stage2_12[90]}
   );
   gpc606_5 gpc1397 (
      {stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[28],stage2_14[51],stage2_13[65],stage2_12[91]}
   );
   gpc606_5 gpc1398 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199], stage1_12[200]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[29],stage2_14[52],stage2_13[66],stage2_12[92]}
   );
   gpc606_5 gpc1399 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[30],stage2_14[53],stage2_13[67]}
   );
   gpc606_5 gpc1400 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[8],stage2_15[31],stage2_14[54],stage2_13[68]}
   );
   gpc615_5 gpc1401 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154]},
      {stage1_14[42]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[9],stage2_15[32],stage2_14[55],stage2_13[69]}
   );
   gpc615_5 gpc1402 (
      {stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159]},
      {stage1_14[43]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[10],stage2_15[33],stage2_14[56],stage2_13[70]}
   );
   gpc615_5 gpc1403 (
      {stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage1_14[44]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[11],stage2_15[34],stage2_14[57],stage2_13[71]}
   );
   gpc615_5 gpc1404 (
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169]},
      {stage1_14[45]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[12],stage2_15[35],stage2_14[58],stage2_13[72]}
   );
   gpc615_5 gpc1405 (
      {stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174]},
      {stage1_14[46]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[13],stage2_15[36],stage2_14[59],stage2_13[73]}
   );
   gpc615_5 gpc1406 (
      {stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_14[47]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[14],stage2_15[37],stage2_14[60],stage2_13[74]}
   );
   gpc615_5 gpc1407 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[48]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[15],stage2_15[38],stage2_14[61],stage2_13[75]}
   );
   gpc615_5 gpc1408 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[49]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[16],stage2_15[39],stage2_14[62],stage2_13[76]}
   );
   gpc615_5 gpc1409 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[50]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[17],stage2_15[40],stage2_14[63],stage2_13[77]}
   );
   gpc615_5 gpc1410 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[51]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[18],stage2_15[41],stage2_14[64],stage2_13[78]}
   );
   gpc615_5 gpc1411 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[52]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[19],stage2_15[42],stage2_14[65],stage2_13[79]}
   );
   gpc615_5 gpc1412 (
      {stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage1_14[53]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[20],stage2_15[43],stage2_14[66],stage2_13[80]}
   );
   gpc615_5 gpc1413 (
      {stage1_13[210], stage1_13[211], stage1_13[212], stage1_13[213], stage1_13[214]},
      {stage1_14[54]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[21],stage2_15[44],stage2_14[67],stage2_13[81]}
   );
   gpc615_5 gpc1414 (
      {stage1_13[215], stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219]},
      {stage1_14[55]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[22],stage2_15[45],stage2_14[68],stage2_13[82]}
   );
   gpc615_5 gpc1415 (
      {stage1_13[220], stage1_13[221], stage1_13[222], stage1_13[223], stage1_13[224]},
      {stage1_14[56]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[23],stage2_15[46],stage2_14[69],stage2_13[83]}
   );
   gpc615_5 gpc1416 (
      {stage1_13[225], stage1_13[226], stage1_13[227], stage1_13[228], stage1_13[229]},
      {stage1_14[57]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[24],stage2_15[47],stage2_14[70],stage2_13[84]}
   );
   gpc615_5 gpc1417 (
      {stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233], stage1_13[234]},
      {stage1_14[58]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[25],stage2_15[48],stage2_14[71],stage2_13[85]}
   );
   gpc606_5 gpc1418 (
      {stage1_14[59], stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[19],stage2_16[26],stage2_15[49],stage2_14[72]}
   );
   gpc606_5 gpc1419 (
      {stage1_14[65], stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[20],stage2_16[27],stage2_15[50],stage2_14[73]}
   );
   gpc606_5 gpc1420 (
      {stage1_14[71], stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[21],stage2_16[28],stage2_15[51],stage2_14[74]}
   );
   gpc606_5 gpc1421 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[22],stage2_16[29],stage2_15[52],stage2_14[75]}
   );
   gpc606_5 gpc1422 (
      {stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[23],stage2_16[30],stage2_15[53],stage2_14[76]}
   );
   gpc606_5 gpc1423 (
      {stage1_14[89], stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[24],stage2_16[31],stage2_15[54],stage2_14[77]}
   );
   gpc606_5 gpc1424 (
      {stage1_14[95], stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[25],stage2_16[32],stage2_15[55],stage2_14[78]}
   );
   gpc606_5 gpc1425 (
      {stage1_14[101], stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[26],stage2_16[33],stage2_15[56],stage2_14[79]}
   );
   gpc606_5 gpc1426 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[27],stage2_16[34],stage2_15[57],stage2_14[80]}
   );
   gpc606_5 gpc1427 (
      {stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[28],stage2_16[35],stage2_15[58],stage2_14[81]}
   );
   gpc615_5 gpc1428 (
      {stage1_14[119], stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123]},
      {stage1_15[114]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[29],stage2_16[36],stage2_15[59],stage2_14[82]}
   );
   gpc615_5 gpc1429 (
      {stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[115]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[30],stage2_16[37],stage2_15[60],stage2_14[83]}
   );
   gpc615_5 gpc1430 (
      {stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_15[116]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[31],stage2_16[38],stage2_15[61],stage2_14[84]}
   );
   gpc615_5 gpc1431 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138]},
      {stage1_15[117]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[32],stage2_16[39],stage2_15[62],stage2_14[85]}
   );
   gpc615_5 gpc1432 (
      {stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage1_15[118]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[33],stage2_16[40],stage2_15[63],stage2_14[86]}
   );
   gpc615_5 gpc1433 (
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148]},
      {stage1_15[119]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[34],stage2_16[41],stage2_15[64],stage2_14[87]}
   );
   gpc615_5 gpc1434 (
      {stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153]},
      {stage1_15[120]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[35],stage2_16[42],stage2_15[65],stage2_14[88]}
   );
   gpc615_5 gpc1435 (
      {stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_15[121]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[36],stage2_16[43],stage2_15[66],stage2_14[89]}
   );
   gpc615_5 gpc1436 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_15[122]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[37],stage2_16[44],stage2_15[67],stage2_14[90]}
   );
   gpc615_5 gpc1437 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168]},
      {stage1_15[123]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[38],stage2_16[45],stage2_15[68],stage2_14[91]}
   );
   gpc615_5 gpc1438 (
      {stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage1_15[124]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[39],stage2_16[46],stage2_15[69],stage2_14[92]}
   );
   gpc606_5 gpc1439 (
      {stage1_15[125], stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[21],stage2_17[40],stage2_16[47],stage2_15[70]}
   );
   gpc606_5 gpc1440 (
      {stage1_15[131], stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[22],stage2_17[41],stage2_16[48],stage2_15[71]}
   );
   gpc606_5 gpc1441 (
      {stage1_15[137], stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[23],stage2_17[42],stage2_16[49],stage2_15[72]}
   );
   gpc606_5 gpc1442 (
      {stage1_15[143], stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[24],stage2_17[43],stage2_16[50],stage2_15[73]}
   );
   gpc606_5 gpc1443 (
      {stage1_15[149], stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[25],stage2_17[44],stage2_16[51],stage2_15[74]}
   );
   gpc1_1 gpc1444 (
      {stage1_0[138]},
      {stage2_0[28]}
   );
   gpc1_1 gpc1445 (
      {stage1_0[139]},
      {stage2_0[29]}
   );
   gpc1_1 gpc1446 (
      {stage1_0[140]},
      {stage2_0[30]}
   );
   gpc1_1 gpc1447 (
      {stage1_0[141]},
      {stage2_0[31]}
   );
   gpc1_1 gpc1448 (
      {stage1_0[142]},
      {stage2_0[32]}
   );
   gpc1_1 gpc1449 (
      {stage1_0[143]},
      {stage2_0[33]}
   );
   gpc1_1 gpc1450 (
      {stage1_0[144]},
      {stage2_0[34]}
   );
   gpc1_1 gpc1451 (
      {stage1_0[145]},
      {stage2_0[35]}
   );
   gpc1_1 gpc1452 (
      {stage1_0[146]},
      {stage2_0[36]}
   );
   gpc1_1 gpc1453 (
      {stage1_0[147]},
      {stage2_0[37]}
   );
   gpc1_1 gpc1454 (
      {stage1_1[108]},
      {stage2_1[36]}
   );
   gpc1_1 gpc1455 (
      {stage1_1[109]},
      {stage2_1[37]}
   );
   gpc1_1 gpc1456 (
      {stage1_1[110]},
      {stage2_1[38]}
   );
   gpc1_1 gpc1457 (
      {stage1_1[111]},
      {stage2_1[39]}
   );
   gpc1_1 gpc1458 (
      {stage1_1[112]},
      {stage2_1[40]}
   );
   gpc1_1 gpc1459 (
      {stage1_1[113]},
      {stage2_1[41]}
   );
   gpc1_1 gpc1460 (
      {stage1_1[114]},
      {stage2_1[42]}
   );
   gpc1_1 gpc1461 (
      {stage1_1[115]},
      {stage2_1[43]}
   );
   gpc1_1 gpc1462 (
      {stage1_1[116]},
      {stage2_1[44]}
   );
   gpc1_1 gpc1463 (
      {stage1_1[117]},
      {stage2_1[45]}
   );
   gpc1_1 gpc1464 (
      {stage1_1[118]},
      {stage2_1[46]}
   );
   gpc1_1 gpc1465 (
      {stage1_1[119]},
      {stage2_1[47]}
   );
   gpc1_1 gpc1466 (
      {stage1_1[120]},
      {stage2_1[48]}
   );
   gpc1_1 gpc1467 (
      {stage1_1[121]},
      {stage2_1[49]}
   );
   gpc1_1 gpc1468 (
      {stage1_1[122]},
      {stage2_1[50]}
   );
   gpc1_1 gpc1469 (
      {stage1_1[123]},
      {stage2_1[51]}
   );
   gpc1_1 gpc1470 (
      {stage1_1[124]},
      {stage2_1[52]}
   );
   gpc1_1 gpc1471 (
      {stage1_1[125]},
      {stage2_1[53]}
   );
   gpc1_1 gpc1472 (
      {stage1_1[126]},
      {stage2_1[54]}
   );
   gpc1_1 gpc1473 (
      {stage1_1[127]},
      {stage2_1[55]}
   );
   gpc1_1 gpc1474 (
      {stage1_1[128]},
      {stage2_1[56]}
   );
   gpc1_1 gpc1475 (
      {stage1_1[129]},
      {stage2_1[57]}
   );
   gpc1_1 gpc1476 (
      {stage1_1[130]},
      {stage2_1[58]}
   );
   gpc1_1 gpc1477 (
      {stage1_1[131]},
      {stage2_1[59]}
   );
   gpc1_1 gpc1478 (
      {stage1_1[132]},
      {stage2_1[60]}
   );
   gpc1_1 gpc1479 (
      {stage1_1[133]},
      {stage2_1[61]}
   );
   gpc1_1 gpc1480 (
      {stage1_1[134]},
      {stage2_1[62]}
   );
   gpc1_1 gpc1481 (
      {stage1_2[158]},
      {stage2_2[44]}
   );
   gpc1_1 gpc1482 (
      {stage1_2[159]},
      {stage2_2[45]}
   );
   gpc1_1 gpc1483 (
      {stage1_2[160]},
      {stage2_2[46]}
   );
   gpc1_1 gpc1484 (
      {stage1_2[161]},
      {stage2_2[47]}
   );
   gpc1_1 gpc1485 (
      {stage1_2[162]},
      {stage2_2[48]}
   );
   gpc1_1 gpc1486 (
      {stage1_2[163]},
      {stage2_2[49]}
   );
   gpc1_1 gpc1487 (
      {stage1_2[164]},
      {stage2_2[50]}
   );
   gpc1_1 gpc1488 (
      {stage1_2[165]},
      {stage2_2[51]}
   );
   gpc1_1 gpc1489 (
      {stage1_2[166]},
      {stage2_2[52]}
   );
   gpc1_1 gpc1490 (
      {stage1_2[167]},
      {stage2_2[53]}
   );
   gpc1_1 gpc1491 (
      {stage1_3[236]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1492 (
      {stage1_3[237]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1493 (
      {stage1_3[238]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1494 (
      {stage1_3[239]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1495 (
      {stage1_3[240]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1496 (
      {stage1_3[241]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1497 (
      {stage1_3[242]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1498 (
      {stage1_3[243]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1499 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1500 (
      {stage1_5[322]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1501 (
      {stage1_5[323]},
      {stage2_5[94]}
   );
   gpc1_1 gpc1502 (
      {stage1_5[324]},
      {stage2_5[95]}
   );
   gpc1_1 gpc1503 (
      {stage1_5[325]},
      {stage2_5[96]}
   );
   gpc1_1 gpc1504 (
      {stage1_5[326]},
      {stage2_5[97]}
   );
   gpc1_1 gpc1505 (
      {stage1_5[327]},
      {stage2_5[98]}
   );
   gpc1_1 gpc1506 (
      {stage1_5[328]},
      {stage2_5[99]}
   );
   gpc1_1 gpc1507 (
      {stage1_5[329]},
      {stage2_5[100]}
   );
   gpc1_1 gpc1508 (
      {stage1_5[330]},
      {stage2_5[101]}
   );
   gpc1_1 gpc1509 (
      {stage1_5[331]},
      {stage2_5[102]}
   );
   gpc1_1 gpc1510 (
      {stage1_5[332]},
      {stage2_5[103]}
   );
   gpc1_1 gpc1511 (
      {stage1_5[333]},
      {stage2_5[104]}
   );
   gpc1_1 gpc1512 (
      {stage1_5[334]},
      {stage2_5[105]}
   );
   gpc1_1 gpc1513 (
      {stage1_5[335]},
      {stage2_5[106]}
   );
   gpc1_1 gpc1514 (
      {stage1_5[336]},
      {stage2_5[107]}
   );
   gpc1_1 gpc1515 (
      {stage1_8[185]},
      {stage2_8[95]}
   );
   gpc1_1 gpc1516 (
      {stage1_8[186]},
      {stage2_8[96]}
   );
   gpc1_1 gpc1517 (
      {stage1_8[187]},
      {stage2_8[97]}
   );
   gpc1_1 gpc1518 (
      {stage1_8[188]},
      {stage2_8[98]}
   );
   gpc1_1 gpc1519 (
      {stage1_8[189]},
      {stage2_8[99]}
   );
   gpc1_1 gpc1520 (
      {stage1_8[190]},
      {stage2_8[100]}
   );
   gpc1_1 gpc1521 (
      {stage1_8[191]},
      {stage2_8[101]}
   );
   gpc1_1 gpc1522 (
      {stage1_8[192]},
      {stage2_8[102]}
   );
   gpc1_1 gpc1523 (
      {stage1_8[193]},
      {stage2_8[103]}
   );
   gpc1_1 gpc1524 (
      {stage1_8[194]},
      {stage2_8[104]}
   );
   gpc1_1 gpc1525 (
      {stage1_8[195]},
      {stage2_8[105]}
   );
   gpc1_1 gpc1526 (
      {stage1_10[281]},
      {stage2_10[89]}
   );
   gpc1_1 gpc1527 (
      {stage1_12[201]},
      {stage2_12[93]}
   );
   gpc1_1 gpc1528 (
      {stage1_14[174]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1529 (
      {stage1_14[175]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1530 (
      {stage1_14[176]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1531 (
      {stage1_14[177]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1532 (
      {stage1_14[178]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1533 (
      {stage1_14[179]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1534 (
      {stage1_14[180]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1535 (
      {stage1_14[181]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1536 (
      {stage1_14[182]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1537 (
      {stage1_16[126]},
      {stage2_16[52]}
   );
   gpc1_1 gpc1538 (
      {stage1_16[127]},
      {stage2_16[53]}
   );
   gpc1_1 gpc1539 (
      {stage1_16[128]},
      {stage2_16[54]}
   );
   gpc1_1 gpc1540 (
      {stage1_16[129]},
      {stage2_16[55]}
   );
   gpc1_1 gpc1541 (
      {stage1_16[130]},
      {stage2_16[56]}
   );
   gpc1_1 gpc1542 (
      {stage1_16[131]},
      {stage2_16[57]}
   );
   gpc1_1 gpc1543 (
      {stage1_16[132]},
      {stage2_16[58]}
   );
   gpc1_1 gpc1544 (
      {stage1_16[133]},
      {stage2_16[59]}
   );
   gpc1_1 gpc1545 (
      {stage1_16[134]},
      {stage2_16[60]}
   );
   gpc1_1 gpc1546 (
      {stage1_16[135]},
      {stage2_16[61]}
   );
   gpc1_1 gpc1547 (
      {stage1_16[136]},
      {stage2_16[62]}
   );
   gpc1_1 gpc1548 (
      {stage1_16[137]},
      {stage2_16[63]}
   );
   gpc1_1 gpc1549 (
      {stage1_16[138]},
      {stage2_16[64]}
   );
   gpc1_1 gpc1550 (
      {stage1_16[139]},
      {stage2_16[65]}
   );
   gpc1_1 gpc1551 (
      {stage1_16[140]},
      {stage2_16[66]}
   );
   gpc1_1 gpc1552 (
      {stage1_16[141]},
      {stage2_16[67]}
   );
   gpc1_1 gpc1553 (
      {stage1_16[142]},
      {stage2_16[68]}
   );
   gpc1_1 gpc1554 (
      {stage1_16[143]},
      {stage2_16[69]}
   );
   gpc1_1 gpc1555 (
      {stage1_16[144]},
      {stage2_16[70]}
   );
   gpc1_1 gpc1556 (
      {stage1_16[145]},
      {stage2_16[71]}
   );
   gpc1_1 gpc1557 (
      {stage1_16[146]},
      {stage2_16[72]}
   );
   gpc1_1 gpc1558 (
      {stage1_16[147]},
      {stage2_16[73]}
   );
   gpc1_1 gpc1559 (
      {stage1_16[148]},
      {stage2_16[74]}
   );
   gpc1_1 gpc1560 (
      {stage1_16[149]},
      {stage2_16[75]}
   );
   gpc1_1 gpc1561 (
      {stage1_16[150]},
      {stage2_16[76]}
   );
   gpc1_1 gpc1562 (
      {stage1_17[30]},
      {stage2_17[45]}
   );
   gpc1_1 gpc1563 (
      {stage1_17[31]},
      {stage2_17[46]}
   );
   gpc1_1 gpc1564 (
      {stage1_17[32]},
      {stage2_17[47]}
   );
   gpc1_1 gpc1565 (
      {stage1_17[33]},
      {stage2_17[48]}
   );
   gpc1_1 gpc1566 (
      {stage1_17[34]},
      {stage2_17[49]}
   );
   gpc1_1 gpc1567 (
      {stage1_17[35]},
      {stage2_17[50]}
   );
   gpc1_1 gpc1568 (
      {stage1_17[36]},
      {stage2_17[51]}
   );
   gpc1_1 gpc1569 (
      {stage1_17[37]},
      {stage2_17[52]}
   );
   gpc1_1 gpc1570 (
      {stage1_17[38]},
      {stage2_17[53]}
   );
   gpc1_1 gpc1571 (
      {stage1_17[39]},
      {stage2_17[54]}
   );
   gpc1_1 gpc1572 (
      {stage1_17[40]},
      {stage2_17[55]}
   );
   gpc1_1 gpc1573 (
      {stage1_17[41]},
      {stage2_17[56]}
   );
   gpc1_1 gpc1574 (
      {stage1_17[42]},
      {stage2_17[57]}
   );
   gpc1_1 gpc1575 (
      {stage1_17[43]},
      {stage2_17[58]}
   );
   gpc1_1 gpc1576 (
      {stage1_17[44]},
      {stage2_17[59]}
   );
   gpc1_1 gpc1577 (
      {stage1_17[45]},
      {stage2_17[60]}
   );
   gpc1_1 gpc1578 (
      {stage1_17[46]},
      {stage2_17[61]}
   );
   gpc1_1 gpc1579 (
      {stage1_17[47]},
      {stage2_17[62]}
   );
   gpc1_1 gpc1580 (
      {stage1_17[48]},
      {stage2_17[63]}
   );
   gpc1_1 gpc1581 (
      {stage1_17[49]},
      {stage2_17[64]}
   );
   gpc1_1 gpc1582 (
      {stage1_17[50]},
      {stage2_17[65]}
   );
   gpc1_1 gpc1583 (
      {stage1_17[51]},
      {stage2_17[66]}
   );
   gpc1_1 gpc1584 (
      {stage1_17[52]},
      {stage2_17[67]}
   );
   gpc1_1 gpc1585 (
      {stage1_17[53]},
      {stage2_17[68]}
   );
   gpc1_1 gpc1586 (
      {stage1_17[54]},
      {stage2_17[69]}
   );
   gpc1_1 gpc1587 (
      {stage1_17[55]},
      {stage2_17[70]}
   );
   gpc1_1 gpc1588 (
      {stage1_17[56]},
      {stage2_17[71]}
   );
   gpc1_1 gpc1589 (
      {stage1_17[57]},
      {stage2_17[72]}
   );
   gpc1_1 gpc1590 (
      {stage1_17[58]},
      {stage2_17[73]}
   );
   gpc1_1 gpc1591 (
      {stage1_17[59]},
      {stage2_17[74]}
   );
   gpc1_1 gpc1592 (
      {stage1_17[60]},
      {stage2_17[75]}
   );
   gpc1_1 gpc1593 (
      {stage1_17[61]},
      {stage2_17[76]}
   );
   gpc1_1 gpc1594 (
      {stage1_17[62]},
      {stage2_17[77]}
   );
   gpc1_1 gpc1595 (
      {stage1_17[63]},
      {stage2_17[78]}
   );
   gpc1_1 gpc1596 (
      {stage1_17[64]},
      {stage2_17[79]}
   );
   gpc1_1 gpc1597 (
      {stage1_17[65]},
      {stage2_17[80]}
   );
   gpc1_1 gpc1598 (
      {stage1_17[66]},
      {stage2_17[81]}
   );
   gpc1_1 gpc1599 (
      {stage1_17[67]},
      {stage2_17[82]}
   );
   gpc1_1 gpc1600 (
      {stage1_17[68]},
      {stage2_17[83]}
   );
   gpc1_1 gpc1601 (
      {stage1_17[69]},
      {stage2_17[84]}
   );
   gpc1_1 gpc1602 (
      {stage1_17[70]},
      {stage2_17[85]}
   );
   gpc1_1 gpc1603 (
      {stage1_17[71]},
      {stage2_17[86]}
   );
   gpc1_1 gpc1604 (
      {stage1_17[72]},
      {stage2_17[87]}
   );
   gpc1_1 gpc1605 (
      {stage1_17[73]},
      {stage2_17[88]}
   );
   gpc1_1 gpc1606 (
      {stage1_17[74]},
      {stage2_17[89]}
   );
   gpc1_1 gpc1607 (
      {stage1_17[75]},
      {stage2_17[90]}
   );
   gpc1_1 gpc1608 (
      {stage1_17[76]},
      {stage2_17[91]}
   );
   gpc1_1 gpc1609 (
      {stage1_17[77]},
      {stage2_17[92]}
   );
   gpc1_1 gpc1610 (
      {stage1_17[78]},
      {stage2_17[93]}
   );
   gpc1_1 gpc1611 (
      {stage1_17[79]},
      {stage2_17[94]}
   );
   gpc1_1 gpc1612 (
      {stage1_17[80]},
      {stage2_17[95]}
   );
   gpc1163_5 gpc1613 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc1614 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc1615 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc1616 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1617 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc1618 (
      {stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc1619 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1620 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1621 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1622 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1623 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc1624 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc1625 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc1626 (
      {stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc1627 (
      {stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1628 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1629 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc1630 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[17],stage3_3[17],stage3_2[17]}
   );
   gpc615_5 gpc1631 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc1632 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1633 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1634 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1635 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1636 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc606_5 gpc1637 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[24]}
   );
   gpc606_5 gpc1638 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[25]}
   );
   gpc606_5 gpc1639 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[26]}
   );
   gpc606_5 gpc1640 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[27]}
   );
   gpc606_5 gpc1641 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[28]}
   );
   gpc606_5 gpc1642 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[29]}
   );
   gpc606_5 gpc1643 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[30]}
   );
   gpc606_5 gpc1644 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[31]}
   );
   gpc606_5 gpc1645 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[32]}
   );
   gpc606_5 gpc1646 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[9],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc1647 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[10],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc606_5 gpc1648 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[11],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc606_5 gpc1649 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[12],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc606_5 gpc1650 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[13],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc606_5 gpc1651 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[14],stage3_7[19],stage3_6[26],stage3_5[32]}
   );
   gpc606_5 gpc1652 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[15],stage3_7[20],stage3_6[27],stage3_5[33]}
   );
   gpc606_5 gpc1653 (
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[16],stage3_7[21],stage3_6[28],stage3_5[34]}
   );
   gpc606_5 gpc1654 (
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51], stage2_7[52], stage2_7[53]},
      {stage3_9[8],stage3_8[17],stage3_7[22],stage3_6[29],stage3_5[35]}
   );
   gpc606_5 gpc1655 (
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage3_9[9],stage3_8[18],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc606_5 gpc1656 (
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65]},
      {stage3_9[10],stage3_8[19],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1657 (
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage3_9[11],stage3_8[20],stage3_7[25],stage3_6[32],stage3_5[38]}
   );
   gpc606_5 gpc1658 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77]},
      {stage3_9[12],stage3_8[21],stage3_7[26],stage3_6[33],stage3_5[39]}
   );
   gpc615_5 gpc1659 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[78]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[13],stage3_8[22],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc1660 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[14],stage3_8[23],stage3_7[28],stage3_6[35]}
   );
   gpc615_5 gpc1661 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[80]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[15],stage3_8[24],stage3_7[29],stage3_6[36]}
   );
   gpc615_5 gpc1662 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[81]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[16],stage3_8[25],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1663 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[82]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[17],stage3_8[26],stage3_7[31],stage3_6[38]}
   );
   gpc615_5 gpc1664 (
      {stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87]},
      {stage2_8[30]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[5],stage3_9[18],stage3_8[27],stage3_7[32]}
   );
   gpc615_5 gpc1665 (
      {stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91], stage2_7[92]},
      {stage2_8[31]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[6],stage3_9[19],stage3_8[28],stage3_7[33]}
   );
   gpc615_5 gpc1666 (
      {stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96], stage2_7[97]},
      {stage2_8[32]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[7],stage3_9[20],stage3_8[29],stage3_7[34]}
   );
   gpc615_5 gpc1667 (
      {stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101], stage2_7[102]},
      {stage2_8[33]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[8],stage3_9[21],stage3_8[30],stage3_7[35]}
   );
   gpc606_5 gpc1668 (
      {stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[9],stage3_9[22],stage3_8[31]}
   );
   gpc606_5 gpc1669 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[10],stage3_9[23],stage3_8[32]}
   );
   gpc606_5 gpc1670 (
      {stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[11],stage3_9[24],stage3_8[33]}
   );
   gpc606_5 gpc1671 (
      {stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[12],stage3_9[25],stage3_8[34]}
   );
   gpc606_5 gpc1672 (
      {stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[13],stage3_9[26],stage3_8[35]}
   );
   gpc606_5 gpc1673 (
      {stage2_8[64], stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[14],stage3_9[27],stage3_8[36]}
   );
   gpc606_5 gpc1674 (
      {stage2_8[70], stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[10],stage3_10[15],stage3_9[28],stage3_8[37]}
   );
   gpc606_5 gpc1675 (
      {stage2_8[76], stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[11],stage3_10[16],stage3_9[29],stage3_8[38]}
   );
   gpc606_5 gpc1676 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[12],stage3_10[17],stage3_9[30],stage3_8[39]}
   );
   gpc606_5 gpc1677 (
      {stage2_8[88], stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[13],stage3_10[18],stage3_9[31],stage3_8[40]}
   );
   gpc606_5 gpc1678 (
      {stage2_8[94], stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[14],stage3_10[19],stage3_9[32],stage3_8[41]}
   );
   gpc207_4 gpc1679 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30]},
      {stage2_11[0], stage2_11[1]},
      {stage3_12[11],stage3_11[15],stage3_10[20],stage3_9[33]}
   );
   gpc207_4 gpc1680 (
      {stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37]},
      {stage2_11[2], stage2_11[3]},
      {stage3_12[12],stage3_11[16],stage3_10[21],stage3_9[34]}
   );
   gpc606_5 gpc1681 (
      {stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[0],stage3_12[13],stage3_11[17],stage3_10[22],stage3_9[35]}
   );
   gpc606_5 gpc1682 (
      {stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[1],stage3_12[14],stage3_11[18],stage3_10[23],stage3_9[36]}
   );
   gpc606_5 gpc1683 (
      {stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[2],stage3_12[15],stage3_11[19],stage3_10[24],stage3_9[37]}
   );
   gpc606_5 gpc1684 (
      {stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61]},
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage3_13[3],stage3_12[16],stage3_11[20],stage3_10[25],stage3_9[38]}
   );
   gpc606_5 gpc1685 (
      {stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67]},
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage3_13[4],stage3_12[17],stage3_11[21],stage3_10[26],stage3_9[39]}
   );
   gpc606_5 gpc1686 (
      {stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73]},
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage3_13[5],stage3_12[18],stage3_11[22],stage3_10[27],stage3_9[40]}
   );
   gpc606_5 gpc1687 (
      {stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79]},
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage3_13[6],stage3_12[19],stage3_11[23],stage3_10[28],stage3_9[41]}
   );
   gpc606_5 gpc1688 (
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[7],stage3_12[20],stage3_11[24],stage3_10[29]}
   );
   gpc615_5 gpc1689 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[46]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[8],stage3_12[21],stage3_11[25],stage3_10[30]}
   );
   gpc615_5 gpc1690 (
      {stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_12[12]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[9],stage3_12[22],stage3_11[26]}
   );
   gpc615_5 gpc1691 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_12[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[10],stage3_12[23],stage3_11[27]}
   );
   gpc615_5 gpc1692 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_12[14]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[11],stage3_12[24],stage3_11[28]}
   );
   gpc615_5 gpc1693 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66]},
      {stage2_12[15]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[12],stage3_12[25],stage3_11[29]}
   );
   gpc615_5 gpc1694 (
      {stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage2_12[16]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[6],stage3_13[13],stage3_12[26],stage3_11[30]}
   );
   gpc615_5 gpc1695 (
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76]},
      {stage2_12[17]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[7],stage3_13[14],stage3_12[27],stage3_11[31]}
   );
   gpc615_5 gpc1696 (
      {stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81]},
      {stage2_12[18]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[8],stage3_13[15],stage3_12[28],stage3_11[32]}
   );
   gpc615_5 gpc1697 (
      {stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_12[19]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[9],stage3_13[16],stage3_12[29],stage3_11[33]}
   );
   gpc615_5 gpc1698 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91]},
      {stage2_12[20]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[10],stage3_13[17],stage3_12[30],stage3_11[34]}
   );
   gpc615_5 gpc1699 (
      {stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_12[21]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[11],stage3_13[18],stage3_12[31],stage3_11[35]}
   );
   gpc615_5 gpc1700 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage2_12[22]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[12],stage3_13[19],stage3_12[32],stage3_11[36]}
   );
   gpc615_5 gpc1701 (
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106]},
      {stage2_12[23]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[13],stage3_13[20],stage3_12[33],stage3_11[37]}
   );
   gpc606_5 gpc1702 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[12],stage3_14[14],stage3_13[21],stage3_12[34]}
   );
   gpc606_5 gpc1703 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[13],stage3_14[15],stage3_13[22],stage3_12[35]}
   );
   gpc606_5 gpc1704 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[14],stage3_14[16],stage3_13[23],stage3_12[36]}
   );
   gpc606_5 gpc1705 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[15],stage3_14[17],stage3_13[24],stage3_12[37]}
   );
   gpc606_5 gpc1706 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[16],stage3_14[18],stage3_13[25],stage3_12[38]}
   );
   gpc615_5 gpc1707 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58]},
      {stage2_13[72]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[17],stage3_14[19],stage3_13[26],stage3_12[39]}
   );
   gpc615_5 gpc1708 (
      {stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage2_13[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[18],stage3_14[20],stage3_13[27],stage3_12[40]}
   );
   gpc615_5 gpc1709 (
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68]},
      {stage2_13[74]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[19],stage3_14[21],stage3_13[28],stage3_12[41]}
   );
   gpc615_5 gpc1710 (
      {stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_13[75]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[20],stage3_14[22],stage3_13[29],stage3_12[42]}
   );
   gpc615_5 gpc1711 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78]},
      {stage2_13[76]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[21],stage3_14[23],stage3_13[30],stage3_12[43]}
   );
   gpc615_5 gpc1712 (
      {stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_13[77]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[22],stage3_14[24],stage3_13[31],stage3_12[44]}
   );
   gpc615_5 gpc1713 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_13[78]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[23],stage3_14[25],stage3_13[32],stage3_12[45]}
   );
   gpc615_5 gpc1714 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93]},
      {stage2_13[79]},
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage3_16[12],stage3_15[24],stage3_14[26],stage3_13[33],stage3_12[46]}
   );
   gpc615_5 gpc1715 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[13],stage3_15[25],stage3_14[27]}
   );
   gpc615_5 gpc1716 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[14],stage3_15[26],stage3_14[28]}
   );
   gpc615_5 gpc1717 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[15],stage3_15[27],stage3_14[29]}
   );
   gpc615_5 gpc1718 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[16],stage3_15[28],stage3_14[30]}
   );
   gpc615_5 gpc1719 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], 1'b0},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[17],stage3_15[29],stage3_14[31]}
   );
   gpc615_5 gpc1720 (
      {stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9]},
      {stage2_16[30]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[5],stage3_17[5],stage3_16[18],stage3_15[30]}
   );
   gpc615_5 gpc1721 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[31]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[6],stage3_17[6],stage3_16[19],stage3_15[31]}
   );
   gpc615_5 gpc1722 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[32]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[7],stage3_17[7],stage3_16[20],stage3_15[32]}
   );
   gpc615_5 gpc1723 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[33]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[8],stage3_17[8],stage3_16[21],stage3_15[33]}
   );
   gpc615_5 gpc1724 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[34]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[9],stage3_17[9],stage3_16[22],stage3_15[34]}
   );
   gpc615_5 gpc1725 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[35]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[10],stage3_17[10],stage3_16[23],stage3_15[35]}
   );
   gpc615_5 gpc1726 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[36]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[11],stage3_17[11],stage3_16[24],stage3_15[36]}
   );
   gpc615_5 gpc1727 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[37]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[12],stage3_17[12],stage3_16[25],stage3_15[37]}
   );
   gpc615_5 gpc1728 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[38]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[13],stage3_17[13],stage3_16[26],stage3_15[38]}
   );
   gpc615_5 gpc1729 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[39]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[14],stage3_17[14],stage3_16[27],stage3_15[39]}
   );
   gpc615_5 gpc1730 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[40]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[15],stage3_17[15],stage3_16[28],stage3_15[40]}
   );
   gpc615_5 gpc1731 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[41]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[16],stage3_17[16],stage3_16[29],stage3_15[41]}
   );
   gpc615_5 gpc1732 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[42]},
      {stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77]},
      {stage3_19[12],stage3_18[17],stage3_17[17],stage3_16[30],stage3_15[42]}
   );
   gpc615_5 gpc1733 (
      {stage2_15[70], stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74]},
      {stage2_16[43]},
      {stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83]},
      {stage3_19[13],stage3_18[18],stage3_17[18],stage3_16[31],stage3_15[43]}
   );
   gpc606_5 gpc1734 (
      {stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47], stage2_16[48], stage2_16[49]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[19],stage3_17[19],stage3_16[32]}
   );
   gpc606_5 gpc1735 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[20],stage3_17[20],stage3_16[33]}
   );
   gpc606_5 gpc1736 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[21],stage3_17[21],stage3_16[34]}
   );
   gpc606_5 gpc1737 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[22],stage3_17[22],stage3_16[35]}
   );
   gpc606_5 gpc1738 (
      {stage2_17[84], stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], 1'b0},
      {stage3_21[0],stage3_20[4],stage3_19[18],stage3_18[23],stage3_17[23]}
   );
   gpc1_1 gpc1739 (
      {stage2_0[24]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1740 (
      {stage2_0[25]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1741 (
      {stage2_0[26]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1742 (
      {stage2_0[27]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1743 (
      {stage2_0[28]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1744 (
      {stage2_0[29]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1745 (
      {stage2_0[30]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1746 (
      {stage2_0[31]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1747 (
      {stage2_0[32]},
      {stage3_0[14]}
   );
   gpc1_1 gpc1748 (
      {stage2_0[33]},
      {stage3_0[15]}
   );
   gpc1_1 gpc1749 (
      {stage2_0[34]},
      {stage3_0[16]}
   );
   gpc1_1 gpc1750 (
      {stage2_0[35]},
      {stage3_0[17]}
   );
   gpc1_1 gpc1751 (
      {stage2_0[36]},
      {stage3_0[18]}
   );
   gpc1_1 gpc1752 (
      {stage2_0[37]},
      {stage3_0[19]}
   );
   gpc1_1 gpc1753 (
      {stage2_1[60]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1754 (
      {stage2_1[61]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1755 (
      {stage2_1[62]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1756 (
      {stage2_3[69]},
      {stage3_3[24]}
   );
   gpc1_1 gpc1757 (
      {stage2_3[70]},
      {stage3_3[25]}
   );
   gpc1_1 gpc1758 (
      {stage2_3[71]},
      {stage3_3[26]}
   );
   gpc1_1 gpc1759 (
      {stage2_3[72]},
      {stage3_3[27]}
   );
   gpc1_1 gpc1760 (
      {stage2_3[73]},
      {stage3_3[28]}
   );
   gpc1_1 gpc1761 (
      {stage2_3[74]},
      {stage3_3[29]}
   );
   gpc1_1 gpc1762 (
      {stage2_3[75]},
      {stage3_3[30]}
   );
   gpc1_1 gpc1763 (
      {stage2_3[76]},
      {stage3_3[31]}
   );
   gpc1_1 gpc1764 (
      {stage2_3[77]},
      {stage3_3[32]}
   );
   gpc1_1 gpc1765 (
      {stage2_3[78]},
      {stage3_3[33]}
   );
   gpc1_1 gpc1766 (
      {stage2_3[79]},
      {stage3_3[34]}
   );
   gpc1_1 gpc1767 (
      {stage2_3[80]},
      {stage3_3[35]}
   );
   gpc1_1 gpc1768 (
      {stage2_3[81]},
      {stage3_3[36]}
   );
   gpc1_1 gpc1769 (
      {stage2_3[82]},
      {stage3_3[37]}
   );
   gpc1_1 gpc1770 (
      {stage2_3[83]},
      {stage3_3[38]}
   );
   gpc1_1 gpc1771 (
      {stage2_3[84]},
      {stage3_3[39]}
   );
   gpc1_1 gpc1772 (
      {stage2_3[85]},
      {stage3_3[40]}
   );
   gpc1_1 gpc1773 (
      {stage2_4[101]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1774 (
      {stage2_4[102]},
      {stage3_4[34]}
   );
   gpc1_1 gpc1775 (
      {stage2_4[103]},
      {stage3_4[35]}
   );
   gpc1_1 gpc1776 (
      {stage2_4[104]},
      {stage3_4[36]}
   );
   gpc1_1 gpc1777 (
      {stage2_4[105]},
      {stage3_4[37]}
   );
   gpc1_1 gpc1778 (
      {stage2_4[106]},
      {stage3_4[38]}
   );
   gpc1_1 gpc1779 (
      {stage2_6[79]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1780 (
      {stage2_6[80]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1781 (
      {stage2_6[81]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1782 (
      {stage2_6[82]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1783 (
      {stage2_6[83]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1784 (
      {stage2_6[84]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1785 (
      {stage2_6[85]},
      {stage3_6[45]}
   );
   gpc1_1 gpc1786 (
      {stage2_6[86]},
      {stage3_6[46]}
   );
   gpc1_1 gpc1787 (
      {stage2_6[87]},
      {stage3_6[47]}
   );
   gpc1_1 gpc1788 (
      {stage2_6[88]},
      {stage3_6[48]}
   );
   gpc1_1 gpc1789 (
      {stage2_6[89]},
      {stage3_6[49]}
   );
   gpc1_1 gpc1790 (
      {stage2_8[100]},
      {stage3_8[42]}
   );
   gpc1_1 gpc1791 (
      {stage2_8[101]},
      {stage3_8[43]}
   );
   gpc1_1 gpc1792 (
      {stage2_8[102]},
      {stage3_8[44]}
   );
   gpc1_1 gpc1793 (
      {stage2_8[103]},
      {stage3_8[45]}
   );
   gpc1_1 gpc1794 (
      {stage2_8[104]},
      {stage3_8[46]}
   );
   gpc1_1 gpc1795 (
      {stage2_8[105]},
      {stage3_8[47]}
   );
   gpc1_1 gpc1796 (
      {stage2_9[80]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1797 (
      {stage2_10[77]},
      {stage3_10[31]}
   );
   gpc1_1 gpc1798 (
      {stage2_10[78]},
      {stage3_10[32]}
   );
   gpc1_1 gpc1799 (
      {stage2_10[79]},
      {stage3_10[33]}
   );
   gpc1_1 gpc1800 (
      {stage2_10[80]},
      {stage3_10[34]}
   );
   gpc1_1 gpc1801 (
      {stage2_10[81]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1802 (
      {stage2_10[82]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1803 (
      {stage2_10[83]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1804 (
      {stage2_10[84]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1805 (
      {stage2_10[85]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1806 (
      {stage2_10[86]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1807 (
      {stage2_10[87]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1808 (
      {stage2_10[88]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1809 (
      {stage2_10[89]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1810 (
      {stage2_13[80]},
      {stage3_13[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_13[81]},
      {stage3_13[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_13[82]},
      {stage3_13[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_13[83]},
      {stage3_13[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_13[84]},
      {stage3_13[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_13[85]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_16[68]},
      {stage3_16[36]}
   );
   gpc1_1 gpc1817 (
      {stage2_16[69]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1818 (
      {stage2_16[70]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1819 (
      {stage2_16[71]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1820 (
      {stage2_16[72]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1821 (
      {stage2_16[73]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1822 (
      {stage2_16[74]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1823 (
      {stage2_16[75]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1824 (
      {stage2_16[76]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1825 (
      {stage2_17[90]},
      {stage3_17[24]}
   );
   gpc1_1 gpc1826 (
      {stage2_17[91]},
      {stage3_17[25]}
   );
   gpc1_1 gpc1827 (
      {stage2_17[92]},
      {stage3_17[26]}
   );
   gpc1_1 gpc1828 (
      {stage2_17[93]},
      {stage3_17[27]}
   );
   gpc1_1 gpc1829 (
      {stage2_17[94]},
      {stage3_17[28]}
   );
   gpc1_1 gpc1830 (
      {stage2_17[95]},
      {stage3_17[29]}
   );
   gpc1_1 gpc1831 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1832 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc1406_5 gpc1833 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1834 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10], stage3_0[11]},
      {stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1343_5 gpc1835 (
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[10], stage3_2[11], stage3_2[12], stage3_2[13]},
      {stage3_3[1], stage3_3[2], stage3_3[3]},
      {stage3_4[0]},
      {stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1836 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9]},
      {stage4_5[1],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1837 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13]},
      {stage3_2[14]},
      {stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage4_5[2],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc615_5 gpc1838 (
      {stage3_3[16], stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20]},
      {stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[3],stage4_4[5],stage4_3[5]}
   );
   gpc615_5 gpc1839 (
      {stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25]},
      {stage3_4[2]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[4],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc1840 (
      {stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30]},
      {stage3_4[3]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[2],stage4_5[5],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc1841 (
      {stage3_3[31], stage3_3[32], stage3_3[33], stage3_3[34], stage3_3[35]},
      {stage3_4[4]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage4_7[3],stage4_6[3],stage4_5[6],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc1842 (
      {stage3_3[36], stage3_3[37], stage3_3[38], stage3_3[39], stage3_3[40]},
      {stage3_4[5]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage4_7[4],stage4_6[4],stage4_5[7],stage4_4[9],stage4_3[9]}
   );
   gpc1415_5 gpc1843 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[30]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[5],stage4_6[5],stage4_5[8],stage4_4[10]}
   );
   gpc606_5 gpc1844 (
      {stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[1],stage4_7[6],stage4_6[6],stage4_5[9],stage4_4[11]}
   );
   gpc606_5 gpc1845 (
      {stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22]},
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage4_8[2],stage4_7[7],stage4_6[7],stage4_5[10],stage4_4[12]}
   );
   gpc615_5 gpc1846 (
      {stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[31]},
      {stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21]},
      {stage4_8[3],stage4_7[8],stage4_6[8],stage4_5[11],stage4_4[13]}
   );
   gpc615_5 gpc1847 (
      {stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_5[32]},
      {stage3_6[22], stage3_6[23], stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27]},
      {stage4_8[4],stage4_7[9],stage4_6[9],stage4_5[12],stage4_4[14]}
   );
   gpc615_5 gpc1848 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37]},
      {stage3_5[33]},
      {stage3_6[28], stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage4_8[5],stage4_7[10],stage4_6[10],stage4_5[13],stage4_4[15]}
   );
   gpc606_5 gpc1849 (
      {stage3_5[34], stage3_5[35], stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39]},
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage4_9[0],stage4_8[6],stage4_7[11],stage4_6[11],stage4_5[14]}
   );
   gpc615_5 gpc1850 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[7],stage4_7[12],stage4_6[12]}
   );
   gpc615_5 gpc1851 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[8]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[8],stage4_7[13],stage4_6[13]}
   );
   gpc615_5 gpc1852 (
      {stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47], stage3_6[48]},
      {stage3_7[9]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[9],stage4_7[14],stage4_6[14]}
   );
   gpc615_5 gpc1853 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[18]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[4],stage4_8[10],stage4_7[15]}
   );
   gpc615_5 gpc1854 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[19]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[5],stage4_8[11],stage4_7[16]}
   );
   gpc615_5 gpc1855 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[20]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[6],stage4_8[12],stage4_7[17]}
   );
   gpc615_5 gpc1856 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[21]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[7],stage4_8[13],stage4_7[18]}
   );
   gpc615_5 gpc1857 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[22]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[8],stage4_8[14],stage4_7[19]}
   );
   gpc606_5 gpc1858 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[5],stage4_10[8],stage4_9[9],stage4_8[15]}
   );
   gpc606_5 gpc1859 (
      {stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[6],stage4_10[9],stage4_9[10],stage4_8[16]}
   );
   gpc606_5 gpc1860 (
      {stage3_8[35], stage3_8[36], stage3_8[37], stage3_8[38], stage3_8[39], stage3_8[40]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[7],stage4_10[10],stage4_9[11],stage4_8[17]}
   );
   gpc606_5 gpc1861 (
      {stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45], stage3_8[46]},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[8],stage4_10[11],stage4_9[12],stage4_8[18]}
   );
   gpc606_5 gpc1862 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[9],stage4_10[12],stage4_9[13]}
   );
   gpc606_5 gpc1863 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[10],stage4_10[13],stage4_9[14]}
   );
   gpc615_5 gpc1864 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[6],stage4_11[11],stage4_10[14]}
   );
   gpc615_5 gpc1865 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[7],stage4_11[12],stage4_10[15]}
   );
   gpc615_5 gpc1866 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[4],stage4_12[8],stage4_11[13],stage4_10[16]}
   );
   gpc615_5 gpc1867 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[15]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[5],stage4_12[9],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1868 (
      {stage3_11[16], stage3_11[17], stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[4],stage4_13[6],stage4_12[10],stage4_11[15]}
   );
   gpc606_5 gpc1869 (
      {stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[5],stage4_13[7],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc1870 (
      {stage3_11[28], stage3_11[29], stage3_11[30], stage3_11[31], stage3_11[32]},
      {stage3_12[24]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[6],stage4_13[8],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc1871 (
      {stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37]},
      {stage3_12[25]},
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage4_15[3],stage4_14[7],stage4_13[9],stage4_12[13],stage4_11[18]}
   );
   gpc117_4 gpc1872 (
      {stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32]},
      {stage3_13[24]},
      {stage3_14[0]},
      {stage4_15[4],stage4_14[8],stage4_13[10],stage4_12[14]}
   );
   gpc606_5 gpc1873 (
      {stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[5],stage4_14[9],stage4_13[11],stage4_12[15]}
   );
   gpc606_5 gpc1874 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[6],stage4_14[10],stage4_13[12]}
   );
   gpc606_5 gpc1875 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[7],stage4_14[11],stage4_13[13]}
   );
   gpc606_5 gpc1876 (
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[8],stage4_14[12]}
   );
   gpc615_5 gpc1877 (
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage3_15[12]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[9],stage4_14[13]}
   );
   gpc615_5 gpc1878 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22]},
      {stage3_15[13]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[10],stage4_14[14]}
   );
   gpc615_5 gpc1879 (
      {stage3_14[23], stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27]},
      {stage3_15[14]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[11],stage4_14[15]}
   );
   gpc606_5 gpc1880 (
      {stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[12]}
   );
   gpc615_5 gpc1881 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[24]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[13]}
   );
   gpc615_5 gpc1882 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[25]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[14]}
   );
   gpc606_5 gpc1883 (
      {stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29], stage3_16[30], stage3_16[31]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[7],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc1884 (
      {stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35], stage3_16[36], stage3_16[37]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[8],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc1885 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[9],stage4_17[11]}
   );
   gpc606_5 gpc1886 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[10],stage4_17[12]}
   );
   gpc1_1 gpc1887 (
      {stage3_0[12]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1888 (
      {stage3_0[13]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1889 (
      {stage3_0[14]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1890 (
      {stage3_0[15]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1891 (
      {stage3_0[16]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1892 (
      {stage3_0[17]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1893 (
      {stage3_0[18]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1894 (
      {stage3_0[19]},
      {stage4_0[9]}
   );
   gpc1_1 gpc1895 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1896 (
      {stage3_2[15]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1897 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1898 (
      {stage3_2[17]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1899 (
      {stage3_2[18]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1900 (
      {stage3_4[38]},
      {stage4_4[16]}
   );
   gpc1_1 gpc1901 (
      {stage3_6[49]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1902 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc1903 (
      {stage3_8[47]},
      {stage4_8[19]}
   );
   gpc1_1 gpc1904 (
      {stage3_9[42]},
      {stage4_9[15]}
   );
   gpc1_1 gpc1905 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc1906 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc1907 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc1908 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc1909 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc1910 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc1911 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc1912 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc1913 (
      {stage3_13[37]},
      {stage4_13[14]}
   );
   gpc1_1 gpc1914 (
      {stage3_13[38]},
      {stage4_13[15]}
   );
   gpc1_1 gpc1915 (
      {stage3_13[39]},
      {stage4_13[16]}
   );
   gpc1_1 gpc1916 (
      {stage3_14[28]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1917 (
      {stage3_14[29]},
      {stage4_14[17]}
   );
   gpc1_1 gpc1918 (
      {stage3_14[30]},
      {stage4_14[18]}
   );
   gpc1_1 gpc1919 (
      {stage3_14[31]},
      {stage4_14[19]}
   );
   gpc1_1 gpc1920 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc1921 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc1922 (
      {stage3_15[33]},
      {stage4_15[17]}
   );
   gpc1_1 gpc1923 (
      {stage3_15[34]},
      {stage4_15[18]}
   );
   gpc1_1 gpc1924 (
      {stage3_15[35]},
      {stage4_15[19]}
   );
   gpc1_1 gpc1925 (
      {stage3_15[36]},
      {stage4_15[20]}
   );
   gpc1_1 gpc1926 (
      {stage3_15[37]},
      {stage4_15[21]}
   );
   gpc1_1 gpc1927 (
      {stage3_15[38]},
      {stage4_15[22]}
   );
   gpc1_1 gpc1928 (
      {stage3_15[39]},
      {stage4_15[23]}
   );
   gpc1_1 gpc1929 (
      {stage3_15[40]},
      {stage4_15[24]}
   );
   gpc1_1 gpc1930 (
      {stage3_15[41]},
      {stage4_15[25]}
   );
   gpc1_1 gpc1931 (
      {stage3_15[42]},
      {stage4_15[26]}
   );
   gpc1_1 gpc1932 (
      {stage3_15[43]},
      {stage4_15[27]}
   );
   gpc1_1 gpc1933 (
      {stage3_16[38]},
      {stage4_16[12]}
   );
   gpc1_1 gpc1934 (
      {stage3_16[39]},
      {stage4_16[13]}
   );
   gpc1_1 gpc1935 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc1936 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc1937 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc1938 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc1939 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc1940 (
      {stage3_18[12]},
      {stage4_18[11]}
   );
   gpc1_1 gpc1941 (
      {stage3_18[13]},
      {stage4_18[12]}
   );
   gpc1_1 gpc1942 (
      {stage3_18[14]},
      {stage4_18[13]}
   );
   gpc1_1 gpc1943 (
      {stage3_18[15]},
      {stage4_18[14]}
   );
   gpc1_1 gpc1944 (
      {stage3_18[16]},
      {stage4_18[15]}
   );
   gpc1_1 gpc1945 (
      {stage3_18[17]},
      {stage4_18[16]}
   );
   gpc1_1 gpc1946 (
      {stage3_18[18]},
      {stage4_18[17]}
   );
   gpc1_1 gpc1947 (
      {stage3_18[19]},
      {stage4_18[18]}
   );
   gpc1_1 gpc1948 (
      {stage3_18[20]},
      {stage4_18[19]}
   );
   gpc1_1 gpc1949 (
      {stage3_18[21]},
      {stage4_18[20]}
   );
   gpc1_1 gpc1950 (
      {stage3_18[22]},
      {stage4_18[21]}
   );
   gpc1_1 gpc1951 (
      {stage3_18[23]},
      {stage4_18[22]}
   );
   gpc1_1 gpc1952 (
      {stage3_18[24]},
      {stage4_18[23]}
   );
   gpc1_1 gpc1953 (
      {stage3_18[25]},
      {stage4_18[24]}
   );
   gpc1_1 gpc1954 (
      {stage3_19[12]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1955 (
      {stage3_19[13]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1956 (
      {stage3_19[14]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1957 (
      {stage3_19[15]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1958 (
      {stage3_19[16]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1959 (
      {stage3_19[17]},
      {stage4_19[12]}
   );
   gpc1_1 gpc1960 (
      {stage3_19[18]},
      {stage4_19[13]}
   );
   gpc1_1 gpc1961 (
      {stage3_20[0]},
      {stage4_20[4]}
   );
   gpc1_1 gpc1962 (
      {stage3_20[1]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1963 (
      {stage3_20[2]},
      {stage4_20[6]}
   );
   gpc1_1 gpc1964 (
      {stage3_20[3]},
      {stage4_20[7]}
   );
   gpc1_1 gpc1965 (
      {stage3_20[4]},
      {stage4_20[8]}
   );
   gpc1_1 gpc1966 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc615_5 gpc1967 (
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4]},
      {stage4_4[0]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0]}
   );
   gpc2135_5 gpc1968 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[6], stage4_5[7], stage4_5[8]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1],stage5_4[1]}
   );
   gpc2135_5 gpc1969 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_6[1]},
      {stage4_7[2], stage4_7[3]},
      {stage5_8[1],stage5_7[2],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc2135_5 gpc1970 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[2]},
      {stage4_7[4], stage4_7[5]},
      {stage5_8[2],stage5_7[3],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc615_5 gpc1971 (
      {stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[4]}
   );
   gpc615_5 gpc1972 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage4_7[7]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[5]}
   );
   gpc2116_5 gpc1973 (
      {stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13]},
      {stage4_8[12]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[5],stage5_7[6]}
   );
   gpc606_5 gpc1974 (
      {stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[6],stage5_7[7]}
   );
   gpc623_5 gpc1975 (
      {stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4]}
   );
   gpc623_5 gpc1976 (
      {stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc1977 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6]}
   );
   gpc606_5 gpc1978 (
      {stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc7_3 gpc1979 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage5_13[4],stage5_12[4],stage5_11[6]}
   );
   gpc606_5 gpc1980 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[5],stage5_12[5]}
   );
   gpc606_5 gpc1981 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1982 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[7]}
   );
   gpc606_5 gpc1983 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[8]}
   );
   gpc615_5 gpc1984 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16]},
      {stage4_14[12]},
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[9]}
   );
   gpc7_3 gpc1985 (
      {stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19]},
      {stage5_16[5],stage5_15[5],stage5_14[7]}
   );
   gpc1163_5 gpc1986 (
      {stage4_15[18], stage4_15[19], stage4_15[20]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0]},
      {stage4_18[0]},
      {stage5_19[0],stage5_18[0],stage5_17[3],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc1987 (
      {stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25]},
      {stage4_16[6]},
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6]},
      {stage5_19[1],stage5_18[1],stage5_17[4],stage5_16[7],stage5_15[7]}
   );
   gpc606_5 gpc1988 (
      {stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[2],stage5_18[2],stage5_17[5],stage5_16[8]}
   );
   gpc606_5 gpc1989 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage5_20[1],stage5_19[3],stage5_18[3],stage5_17[6],stage5_16[9]}
   );
   gpc606_5 gpc1990 (
      {stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[4],stage5_18[4],stage5_17[7]}
   );
   gpc2135_5 gpc1991 (
      {stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[3],stage5_19[5],stage5_18[5]}
   );
   gpc117_4 gpc1992 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22], stage4_18[23], stage4_18[24]},
      {stage4_19[9]},
      {stage4_20[1]},
      {stage5_21[2],stage5_20[4],stage5_19[6],stage5_18[6]}
   );
   gpc1_1 gpc1993 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1994 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1995 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1996 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1997 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1998 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1999 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc2000 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc2001 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc2002 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc2003 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2004 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2005 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc2006 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc2007 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc2008 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc2009 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc2010 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2011 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2012 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2013 (
      {stage4_2[4]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2014 (
      {stage4_2[5]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2015 (
      {stage4_2[6]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2016 (
      {stage4_2[7]},
      {stage5_2[7]}
   );
   gpc1_1 gpc2017 (
      {stage4_2[8]},
      {stage5_2[8]}
   );
   gpc1_1 gpc2018 (
      {stage4_3[5]},
      {stage5_3[1]}
   );
   gpc1_1 gpc2019 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2020 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2021 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2022 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2023 (
      {stage4_4[16]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2024 (
      {stage4_6[13]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2025 (
      {stage4_6[14]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2026 (
      {stage4_6[15]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2027 (
      {stage4_7[20]},
      {stage5_7[8]}
   );
   gpc1_1 gpc2028 (
      {stage4_8[13]},
      {stage5_8[7]}
   );
   gpc1_1 gpc2029 (
      {stage4_8[14]},
      {stage5_8[8]}
   );
   gpc1_1 gpc2030 (
      {stage4_8[15]},
      {stage5_8[9]}
   );
   gpc1_1 gpc2031 (
      {stage4_8[16]},
      {stage5_8[10]}
   );
   gpc1_1 gpc2032 (
      {stage4_8[17]},
      {stage5_8[11]}
   );
   gpc1_1 gpc2033 (
      {stage4_8[18]},
      {stage5_8[12]}
   );
   gpc1_1 gpc2034 (
      {stage4_8[19]},
      {stage5_8[13]}
   );
   gpc1_1 gpc2035 (
      {stage4_9[13]},
      {stage5_9[6]}
   );
   gpc1_1 gpc2036 (
      {stage4_9[14]},
      {stage5_9[7]}
   );
   gpc1_1 gpc2037 (
      {stage4_9[15]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2038 (
      {stage4_15[26]},
      {stage5_15[8]}
   );
   gpc1_1 gpc2039 (
      {stage4_15[27]},
      {stage5_15[9]}
   );
   gpc1_1 gpc2040 (
      {stage4_19[10]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2041 (
      {stage4_19[11]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2042 (
      {stage4_19[12]},
      {stage5_19[9]}
   );
   gpc1_1 gpc2043 (
      {stage4_19[13]},
      {stage5_19[10]}
   );
   gpc1_1 gpc2044 (
      {stage4_20[2]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2045 (
      {stage4_20[3]},
      {stage5_20[6]}
   );
   gpc1_1 gpc2046 (
      {stage4_20[4]},
      {stage5_20[7]}
   );
   gpc1_1 gpc2047 (
      {stage4_20[5]},
      {stage5_20[8]}
   );
   gpc1_1 gpc2048 (
      {stage4_20[6]},
      {stage5_20[9]}
   );
   gpc1_1 gpc2049 (
      {stage4_20[7]},
      {stage5_20[10]}
   );
   gpc1_1 gpc2050 (
      {stage4_20[8]},
      {stage5_20[11]}
   );
   gpc1_1 gpc2051 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc2135_5 gpc2052 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0]},
      {stage5_3[0], stage5_3[1]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc135_4 gpc2053 (
      {stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[1],stage6_3[1],stage6_2[1]}
   );
   gpc615_5 gpc2054 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0]}
   );
   gpc623_5 gpc2055 (
      {stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[1], stage5_7[2]},
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc615_5 gpc2056 (
      {stage5_7[3], stage5_7[4], stage5_7[5], stage5_7[6], stage5_7[7]},
      {stage5_8[12]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc2057 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[3]}
   );
   gpc615_5 gpc2058 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[4]}
   );
   gpc135_4 gpc2059 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc2135_5 gpc2060 (
      {stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6], stage5_14[7]},
      {stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[3]}
   );
   gpc606_5 gpc2061 (
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage6_19[0],stage6_18[1],stage6_17[1],stage6_16[2],stage6_15[2]}
   );
   gpc7_3 gpc2062 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[2],stage6_17[2],stage6_16[3]}
   );
   gpc615_5 gpc2063 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3]}
   );
   gpc2135_5 gpc2064 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_21[0]},
      {stage5_22[0], 1'b0},
      {stage6_23[0],stage6_22[1],stage6_21[1],stage6_20[1],stage6_19[2]}
   );
   gpc615_5 gpc2065 (
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10]},
      {stage5_20[9]},
      {stage5_21[1], stage5_21[2], stage5_21[3], 1'b0, 1'b0, 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[2],stage6_20[2],stage6_19[3]}
   );
   gpc1_1 gpc2066 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2067 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2068 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2069 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2070 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2071 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2072 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc2073 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc2074 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2075 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2076 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2077 (
      {stage5_3[5]},
      {stage6_3[2]}
   );
   gpc1_1 gpc2078 (
      {stage5_4[1]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2079 (
      {stage5_4[2]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2080 (
      {stage5_4[3]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2081 (
      {stage5_4[4]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2082 (
      {stage5_5[0]},
      {stage6_5[1]}
   );
   gpc1_1 gpc2083 (
      {stage5_5[1]},
      {stage6_5[2]}
   );
   gpc1_1 gpc2084 (
      {stage5_5[2]},
      {stage6_5[3]}
   );
   gpc1_1 gpc2085 (
      {stage5_5[3]},
      {stage6_5[4]}
   );
   gpc1_1 gpc2086 (
      {stage5_6[8]},
      {stage6_6[2]}
   );
   gpc1_1 gpc2087 (
      {stage5_7[8]},
      {stage6_7[3]}
   );
   gpc1_1 gpc2088 (
      {stage5_8[13]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2089 (
      {stage5_9[6]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2090 (
      {stage5_9[7]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2091 (
      {stage5_9[8]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2092 (
      {stage5_13[6]},
      {stage6_13[3]}
   );
   gpc1_1 gpc2093 (
      {stage5_13[7]},
      {stage6_13[4]}
   );
   gpc1_1 gpc2094 (
      {stage5_13[8]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2095 (
      {stage5_13[9]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2096 (
      {stage5_16[8]},
      {stage6_16[4]}
   );
   gpc1_1 gpc2097 (
      {stage5_16[9]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2098 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2099 (
      {stage5_18[6]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2100 (
      {stage5_20[10]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2101 (
      {stage5_20[11]},
      {stage6_20[4]}
   );
   gpc2135_5 gpc2102 (
      {stage6_0[0], stage6_0[1], stage6_0[2], stage6_0[3], stage6_0[4]},
      {stage6_1[0], stage6_1[1], stage6_1[2]},
      {stage6_2[0]},
      {stage6_3[0], stage6_3[1]},
      {stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0],stage7_0[0]}
   );
   gpc615_5 gpc2103 (
      {stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4], 1'b0},
      {stage6_3[2]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage7_6[0],stage7_5[0],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc135_4 gpc2104 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[1],stage7_5[1]}
   );
   gpc1343_5 gpc2105 (
      {stage6_7[1], stage6_7[2], stage6_7[3]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc1343_5 gpc2106 (
      {stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1],stage7_9[1]}
   );
   gpc117_4 gpc2107 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_14[0]},
      {stage6_15[0]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc623_5 gpc2108 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc2109 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[0]},
      {stage6_20[0]},
      {stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1343_5 gpc2110 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc623_5 gpc2111 (
      {stage6_22[1], stage6_22[2], 1'b0},
      {stage6_23[0], stage6_23[1]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_24[0],stage7_23[1],stage7_22[1]}
   );
   gpc1_1 gpc2112 (
      {stage6_0[5]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2113 (
      {stage6_1[3]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2114 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor_CLA486_16 compressor_CLA486_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9f9601d1841e5d7f384f7945b135045b5dcd80d13371dde6177de3efabc9cb3f98e402a606dee3a81d53e3d418544e35cab150930c139a8edc6e4d131295f3cc7847d3e34f701b946128bf7467e003de065962c9242d68599bfed9771bb7289968455ef86cdd6a199ec429d784db49c89abd5028139c70d2090deb51f820f0e2b093c46580356eb8830969ca1b8414d839624fb8bb5fbdf24a859e0bf72c281bd407a20b79e0b141109671cd147ea57245d929b5dff2ec5efb65632aa4bf9a27c302afe1a19ba5ab730bba9ae01bdd602c372a1e5cecb01c53bdfb8081e8f9c83d8c586f6459649b5c934ca8144a714a64bd513d7930645a6128baa26403aa1b98bd22734e13217f2f985f236e63dfc5253fc0c5a7176a9c3fae40deffda982f1a7519f4ae88a7c31a6c786d8c8d0e63b54f46be680335c84f109aeac63e42727f7d6c5b51b35ac98ad4dfce94b31b5a567edd3c615da3fc86cae68046a0c73a25d580df4eca9155b04d3ad6d820a689d8ace7312595c3841fbf3c61e1d9814e43c17a500096796e67fedd42c2db4a574e714221caf61c243aa9d597b4d6e187b61589e08e7a09b586397e6e18ab9aa666fd6549e712f55d2f06f0a67e87de16b46fe5dffd24add52ce048ed0b66be629f1d44b6fd98a487e0672ccfe4b5d5201aab9883e3560cf5fecfded188d8059c92e3c348a8309da1e26b833b06d08846cc317fcdf50e924ef4f7d7105f22877c6cbd46a10577eac1677e4e298895c5e577b1d8fe2a4622f196855bd97523da8c57fe218c6674fd7e5a36224c5910619f7c3568ff0e14c9588c91a4f97a4d98c780ea1e315021cd44a0993ffc1fa0c3ae20d320a0dc864c5e7234c090c0dfdbc4dd041cc62c868d3c247741cc55f0d09fde33b40b99e199dddd7e23c09330a565b4a302222ae53952a33b2a7605a18808aad8c0dd51fa5f1f08a78bc7e1f18e1bf9c8e8ed2ea6a5f84dad8ab998051dde5f7d64d3149a1303a5075c2de370ab7087ffa8ecf3e8d865e53ccfb8a169808e474c3256fdc2f031ecf9aa8e03c8302d98ae22b25687fd76adf553b4a843e425f085249e98b226463fb93439b10cabca1b46d2a09a7afb034aed85f7e2b3d4eca0909e34a73a9c1c1b7cf32da8e5dfb85be2af48761399e4320a4a6178b201a94db2cf5adb110ec7f74a7f2d737ac312befa15b64e13f2b69d7fed02b1556918968203a3921eec4a42d1422c46c5690da904231ef5f75c5d4db05cfc78eb0613dd1ea950a54a5ce60ceba9422468ecb4ac73bc607560a1d6c34438874dd9b2a2a411e7aede13807c96f552d8299bb2915ab99748c921245ffad0feedef21bfed2f5aad33d20017ebb851f372;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd045f9396e1ad7b8ec9cba62116936cdd87a537069981c4d82377a7aeb90b44b9b3ef1595c01f37bc08c5e8c66b6a1a7f107c9d2082a098a112a72be0704bb84287d8825941a79a21d3be34dd3baa2a444952875ec07845b32e52974dd218c37397365632d1beae26e4b1d8296e26d1ab50be6139c0e16faa3d50f3140fae1db86c777622014a60cf4945f58c327aad9e8f2d419b6d2009b18eb94410c2faa0b611445bbd032939fb1cfc3caeb0fb6b1cc66e322904e2419cb99a44040625d4c2ba6c6f22e77a46465b5c2a0e8ae1f8c660ef3fe740b62130de516faa9087b26bbc77ded1541057b4d134b416f1de61f6b3ecfd96aee092da29db77476f1c6866e90e7e0bae7abe3f90e070865ff8404fa41cedc5b60082d524bbc03365e93f690f00542d1bd3930db1fea5f8dcf3c0764758bfb6f70f434ea343722200bb868008adf855a36f0b64492ca4ead6e2e645ccdcc44095fad8f8c374f8a0476499c0f5fdbc0fa7b4a911b06aae4c8d7b0ebf4e9237113d129d2ed9e222958fa8cce63a6bb8023921dddfb272674aacdc1e56de940c5ff926e47f894cd3843e3d81fdf7b3c92412950634e1f182503ec05242e636a3df50f06ad904ad8839067d5a3b3d87053d8d30817e2731d6f7268f1d69e07f864fd9e838e899ca0e76006fc76f0042bdccd7b84a4a1b117e793376459f420fe81f28943de50340caea67edec06b54ce773d1a8e42f9c4b189f0f4d27d9992c082360107faf62e19bd18831b785155b9a55c5ec74180c38e89c09ffb579c577c5f0b1f532bc06739c3aa7ea3ceaf6dfb00273caeaff3a5767f27ac9582c74a4a1ba6b74233cb4a7c00e9b7e77a8eb3952b1a4df681d62e7c5c6dda53e763659c803ca9b9a9ffafbe126b137943ebffe179da7f3c7d767ae049db42cc1ed4d1fd7cc0940a5ff386a4700d21597350ae90d81e451dccdcec4acafbfa061b386a39ac2c5e79b0f557962172a10cc374f4093db803a611f501f0b83a129a5ef9e8cd18adc2ce7446873a9b97a69531add49872bc6cd99f14dc127b865b84410040ef11aec81efccbd6028ebb2d24b75c4de0e441980eff8cf2db027de0e2d068738ddfa858c7ff54252599c21aa3a8333e2f69f8ca9d3bbaddd95a2710832c6746dc6fea133a3deec9edb4f027bfedc1dd542af6502da557d0892ab00ef5427d818f1e9971a4a53c892761707765dc6e7a659f60b83a5ef1e7330ec88cee4a091c5d2f3ce3abe104d9dde9fc2f4ab1cd42cc6efd38bbe0b1c331b2e4fa28d8b6760fc973f61c01fe0cc18f915d1f31185b1170e0645dc9e709135e97ffd4c153fb548555c2b8ee7f395dc187526cb5c8b9a67c2c6d6232f3caacb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb52fd36a45d8824e30b1c125c1ee33ca1726c5eb3ad52abdf4638705dd3d9c154c78919b128edccc20d7e5fcb6b2696d91f7a9ebe2b159ea4d53bf20549cb16960667e4a08e99e76a79c36f452f019116172eb94c4791d7ef8d727d17b8fd0512c69858b6a969bbe4cf8a09caa21d98bdba9ba93648dcc87f88b4161ab861d08ef0322f6e0e9d22899aee267addec58ebef7e0843710e0310745002f0dfd3ee9002d8f68d24a8a0c9b519109af74c3c8a80b35cf383d4ae979cc0f67b3b53f454c4ca4d77dfad48100d340f0630a4330ffc434e7e0a68e1989013eb80addfa788263f04b7f3fcaa4cc3eabba57d672d5b0340a3662253e959cabb7cf4f89e9dc12fa45d635376591f702df1cdc202c576f6ea00a785f53bed4ac511eac530d13a0367be947d52088dd9a1a160e831220834ecee8b02c7642f14ab264b6f2a2d962d82d5f5e36a3b9c592af4f4f1a682de623b248bc58c785399c12ee9d9179ea3074213b503becbe652c421b7a1f89450b58c256e695deb19d8fd20f29b10eace1ff66b80a210d2e90807804e95faf2c50d7c064851464d43b3d69eaa6d64f17810140a0cc1602d0fd2b7d625ae8345f540de380e4fc23069e7001f8e469471ef99b66a06b44ac00949b4400c2298e55328b61d5ae7bf8957cddfcb581242653344b19e98dc21c7c523fffa66d19ee71a9a867c1467a2bca8dbbd731cb53344f4e3d004c77a05f6de046a865d54bcad6c15d64f55037b4a52a7e771515f22eacf109e87103af96cdebd84a44944b0383272a7fe997e0f7674b66c5a1b70ccbb89537af9b7a1258b14dc39e766ba6ea709dcb87b996bbc4eddbf964bfc58f3ca15edbad89b712f679d61aaccc770a5a1d25a7d7b3e73a27e2b944ac411ddca5743ec6d8a883baa3252e7aec60678e4e3dec14b7c581c2c3ccb9af7e86742eeaea1f8283127c1f4ac2e48911d798cee8a017272e63c6cbbd3cf52cdb2774d2faa56145ec47a4d3404076bbadf904ada09a3e7131806e2041a2ae1d2be5dda21604945d4de6542108bb1c442a769161c9ba31f8cdd4a4e984a9cc95011a652c68d8825ede1a3cd3a31ade4f94bbd674822b1620d8375f883c7754299daa9870b434d085b22fe6a5b363ef4d7b6684166b43df77b88d405a31ecd19e1f2d9ec63c647f75d7d86c761225159488f1e065bbeafbcc690d61a2fabc54aabb0b999a4ec4aa90d9a07069604382fab1424084877d1b82af2bb070d83abc8f4c840b4f6d7771a8cca2d557ca152bd6d4292f7ffa1b77fbf177ebfc5f148d01fbed3748a101df2ceee6a5d297d6ec67b567db6e51ff25f3f8f75269f2e38d07e74b891bd9a4b5a6218bb1ef50405240767e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5f4dc038fc87d691eb8509744e8bd3c98cf367ac7296a665bf629593c784ed728b8fed187d23ceca49539cf193c79311fac57e3f32d14d9b06ff3749381ad39941beefd9c185b09e55e48dfa41138bfc5b32e4c1a709aefe19ab679ff3dd12d8bacd40cd7f186b2008abf9c0b39f2473c4f9a532f608b49f90728430844978e82e49086e4262d31d93ab269f5ac86798ee3bfdc707d087a91c7ab0a95e15b668b9355b49d844d872f8ddba385fff9fbdb12488c1c56a1d361dffd6779242247e8b3963a6085c55640e405c6515f32a019dcd63bfcf46565c9559439d196c16aa14bd7cf8b7dc371c17ddd841387ba451a287409bae9c0c52857a216285e9dc0d1b03626fd7a6b4c530ad98f614f9a4af30f17d0f86b66271e20a84f207b6750e4bd90986d4aadbc1ae77999fc0249206716edb54456dcf9313677a564244fe22fa83ea885665f941f7da6e35435a84b86d1f9c7ef15aa93d3f071d9eb5b41b29ee6688ca8b7269303ad485c4d268ca30b8fb54e135a933b8a0883b578a4d315e7470e3c2cd68a1a699768fdf9f498ed1f787a0a77ff994d3347955ac00b565757e4996e8930740036593b69c169161b5eb6002ecb5266599fbdfe6688097f339960859ea9841699110f9f1a7859023bebe3e6ab5cbfc3ee9237929a7a8d22bfc2cc68b12e8f41c0c78f4f099a2c9260f0cd692ec00803d44b59d959c82ab03d5a33a6240439b114e357be71e42228ae635c8042af0e03942755c1c27d564df990a945804428d14810acca69e04e8b73bbaea6d40b73a2b9784b9b6744bda23b1abf46e63881ba891aed7695ade64514dd77aac3972862fe068045e099f79c8a910332a57a6be4ccf434d19813c72e71974ac8f5dbcc05eb0aa4ec8f54d1e95f8636d1b876d625e4ca986eec43965c880eb005d4b1d9b2bd4c3ff9e2f0ce468732656eb0a3157cc511e85e7173bccb1ba0abbaddef0cf1033f670ae5def7bf5775858e870f0aaa7b1b60a907e849aafb9babaa9503ea04575d662c4ab482613f83525c43ba56b593c0a8f819ca5d000e018d40fefcc98aa5e0bd3128b8e355dff4b5145a7000c5de74bba63b8dab384f6e7ccc5506f621855bfc1921480cb16b83818cf4d2f6245ebc8ecf02dd3d1e2ff4b36815c799707964d6effed6cfbb1b22e069f6e9f866c3f99c6e5315b610f2d7de5c5cf2a12e1a7b7116a7e075b01a7b4fb99dd342b0ff81eaf297dd95891e4b5c66738b2aa8ce036d7f332b60dcd9016bba2dcb05bdcf8fc26326d77eb9779ce51d565b44938ce3682c95a32eb1c0f1f9accc0847d2d786dbfa574f1b03d23a5b6944b1c62249854448735240d6e407dcd6573b68e4dfb2f7c1099;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3ad85cd20e6f767d12b74fa213d9cb413e3416562a2d4a0fef3fe4ebe9ab0df7584d7d6b3fa0acfee5469ad08890c968a9bbf2c1fc704ab1c44d077158fc394e58470bea2b6c489881c3baca86082a8afd0e3ab30576c8565444a21701d991f313b8e1c0026ba4b68a5d2418b3a17d005dce682903384d4252915fe98170136597cbcefb7eb849d573f2a88aab7e018e4598509e4439864d7adfde5ea26312035865e39dfa6ce6b3aa879009736d58ff78944bc14c79161b87f6cb7a20b5551bbec7f4f8bb81f24e03008b8117921e4d4e098a5422c387f4cf63080a211bc6b3cf77f3a1f781d14add4b3bd5757212a85f621f1fad23bb4c4f09d661becaa31787c9b29c9e787a888e95577bb0fdd0496b824b3700ff56ab01f3dc34a18f6e7bb283e4f44999ac2230c0e8bbfaecfbfca7e2620c0031e0c92eae12ebdbdd0b7739956b53f4424b72e3e1877c83b8f68fc74c26c6b4eff79db0f84cc7af33c8918eb4ab8b31ef4e2ef85ad03156b41a45d7ea58f9b6dd7f3b73dbd224266c26ac789b9f3bbe7edbbdf36ed765146ff861869209654e3b2026c2073402ca68b463f9b747d2525ab356830d7b956879e9c39ad99eebb8be607a74c91a578cd22d89189e73ef37ffddb806e8d7e0c82e1a83552bf5910ebfd0923c5294b26dbb43f0892e2212c8a6dbbb242eae39aefda30f450f57ebb3494a2e00422de2857e589512c368ceb99a65f9d9dafbb6fd782d86a759c9d0ddbc809055f9cc71f919126f47bde166e2b9a59c793337f86395d859c3904c75203ff1d04dab985233cc585a1d01ae804e56dfc1f3a81fc84fcbe8914aaa882ae8a799958b60bdc48342d81ebb005e8424b0063a161ff5f75cdc89b72bd4370e2223d0ec6597ddfc2024b110dded71e9bdd1c0a3d42db01cf214284f99fce2e64d6c176c4f953023840e1d9bd61cd511219912e0c7efa879e1361e2f541b9a9865901f2f287456666fb421fd9c58b9e840bbe4d4a3db763e7641b378c242cefff73ea901cc9eb2e0187e518446a9ed65ae63048c2cb40a0f8b9decfc0aa577911e10d9dfbb6fee890688f30c4dd512c75866c080ebe4e2ba8c8e0d49429e108fd36a1ed9547e4972e99f25b2f55ea38d9e8f42412af3c65bc290c3d79f509e18e5d42fbe38ff2b2776fae20499f6cb5b9bcbc2ff1af7dfc9829af16589032092a0b58ae70d2c1015574926aef341707a3791dd9ac4c77f629bb1b794ca32366d0ddf09b96a8f2df2f9176c56e3a15eb0108b146e2a00a46703a2359e08b738006529198daf1d21d58d3fe6a6ebb7f075ab38a6e30a941987e97d6aeea31038cc990b308fa03ec2e684ee9c1a2ae2d6b986dc404c1415943d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9a9a95610fd1075bedaed217c64ea777b25ccc26f8bd1780ed0eb416a2d652ee8a7561de044917c41c2dfcf5dd774a6d55d34245a041d358ffa2c4f125e92d23ded63971ba30f9ea271f5465c26aaf0fb34249648938a69c7bfe853d920dff5242e84b0c8266a2334e0d46f1bb84fa8b86324913f8dbcaa67fe81003ddb7110c475aaf6738dc17d31449f3265f339dc480bcb2339834840bd02fca1ce81ef994041e4c9ad523fa4426a0dedb546eb67fd1db9694c57791c41ff5eb0c1d217c0aa992afb9fa2817d8fb954e36af272d767aa5be531749d9cae94001bfdcf6d295edab6239762edcc53622bbfa1b515d562fdbff09a8803005d26cd78fa7e8c1c67b446643bfeee83b7bb5b422ab57764745d679737417553ce1bcdc857c345c9b6bef64f56ef671253a062c1b6e9cfcff8b9617655a171c61a7c50f9d61b1a75c0a3bed5f3c82ccbf8fdca889f5c0cb8e80d67aae38d9bf1f22af8780863f5fc48239c55434faae334de8935f8b8c5a4bfbdfc3835839ffbe9b99a790061b27d0b6994d2573860077ca57ed0166007846a1907c748ab59c05148a7563038202b312c6d610a25cec27231a00490ffce440b99612f3d62e8adb8e3071a6235f283888646fa4ba5766b3618db16a70e1e31c6034247ab6e61501390a0c3a9877b72207226bc83da1ee32d737f2b583b4ee747c718dfae85d4aa5d7ec69cec8d3c72e26a56217daf08eafc7b537d5685b92474b25b31709adc2a47b91a4d2446278f7bcc1fd444b8dace9ecd0ef61f0708c0497b777037b357c7af696937d4205394e7edd9a2670d8006a8bebe00139272d9ea99a61ccc2c8d69518658bf93fa5fbf87c5442d8b51d2cd59b8dee55c6f72ec92f5438418ad29d02d255bd4e5b7034fea982fecb842ac08413d185fb69d49d2a54aeb610d9cbcfd4005bbdcf55d78203f2dc1525c4bbfc41fdafbd0b4da172579d6e6f03d5ccf52baa7d780c37f8f0c09ef3c7cca284f8a4d72ae7ab30f47a6b8bd363008a748fa939daed48421eab10c78cd585ac4b2728eb1aead1aaa815020a17b9bb7fa8df18aeb33a8a4e5c49986a8f48ef33d1c107e49012443c502a4f17632b474f85a7061fd04f56b16c60007078b3ecf8ca7f32464c404792d15abf8f8bfb4fa5edf42845aad1636725c07624f7ebebc952aa61d5abb683d0cb14a4a24380f0f5bc87a704528080d0d0c19187f999f915bd61f7ae7c5c1fb364649d12f9da2dfae53fe47b99eca932baec4d0cf7509a0648fa414acadb4180342412a8d9a82d6e1edebee4005aa263ce2d12fc78c4de6fd09db7612538be9a2404bd7eaf9a6ff9406859ee8d75607693d86cbee1b18f97d45c712b4e328e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3a0108c97ed68932d682e16209f46aac1a49a5ed3492f1b504958c357e7935356cc1ffd93e9094eaca09c27cef687c40334fa8efd9d1b1386759dfb4e5add315224f33ed910bbea7c059a3fbf7153081d6a51944c0d892ba8a882b7699594f0f9bfa646931efc8f129febe82e9d9b38a049293b837aee99f91a2f0fb5786dbd23c50110102028ec67b8f65469aad0201f539a96a6998dd9dcc3751731e155bf397463241ba0cd2835d6886447ddd00283829e05d5d6fec7a610a427c666e07411deb9b5f1eca83ed506adf742553b7714f935a21bbf24a7c8b52db3f7afbc1491a8440ac4780b0241713708d23af5630e97443c5f01c96f1098f427244de3ff92dde7fd6227423e4ae101deeb537a22d829cf628e9816235555c07a3732424e3a5d20ac80ba364a870620e10d1e633b176c47e124f39879156153b0c7ab7a19643dee93caa11098aff5b0da9a98fc60c4da3db46ba675caf879c087089f0fc376be401ef4d2bca682b3af97002d2b9d44d88b301865ea041b6eab6fd8e9a510a4fb616693c662184ed2d978290433f366ed59c1a125e5608a9f501724db5243b006d9dc9aa7d544c3f7f15a661c61cc86c814e585c774506da03107e1cbf2b2b1abef2bfe915f9816d4e2d04586609810aac8f5f98d21cc65bdb4f080cf96796b64f71407ae3914f0bd75392ca296034b1ea638f022c454c9e2d80a6cd64f746862eb6aed81a5fedd1746cebf948aa85d9194fb3c14d98b5280ae40f31f4e9373eaaed06e120e315a7a95f4c5be5e50dffd3d463c4ae43ccccf86d32e66bb5cd1230f43c680ed30c5715a2cbbcb5617d31e5838b4faf5bcffbe8d1977c8d88b1d14f0c2c7019bb8f41eabc4b8eb3a74a185c02e0d650b8036030795eb90d1df8908298b58829b89ca2dad80b0044cb1f1dfeb6a3fc6adfa174463be9f54deb368a240730a00faa05656c52b4218d0b564c209379c60eafcd9d3824e134393744394c98c55af0c4cb253f916ff6b8f1b01461ba295be1e56f80f1c8f53ec1a653486bf10ac686c690a04c16ab9b6f46b93ced9d472cf663def3d03d3a2e0d0949e453ee0eec1f53d1ea10dfe7093e7d51d5b2678de68140843ba83b9171bd072307ee7b79f421fc42bcfd9f40d141dc7b0f366a23a06f1f7e05406857c69b737557c07b96dc9575ab0c50da0980e7f2ee93ea59300ee13be52e510144f55b28ab775b7bd260237ce74e9b941e92842690e19a22c8193fa38a0478724b28ea3ad1330d6c8e3b9753ab4d9eeda6ce9f8bba95104bc77c2f9c990cda923d95199e2ea6fb3a6e8dcad2040495775b998835d6410a2feca39dab337efc01348dd7d771a91ec04bd5089ab7503af4fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd9ff734fda1f4cec73458af2fa3949f0c821ae84e30955909f0ca341427799603f25272f7fbbd7328e4f89ac7f2427bec6f6456aed4d7b81794200047db32fa4c5f79cb37f186629efb39c6bd90b2b5b1408bf6920d6d780e0b323afc6f92c837716fbb63dd08908a9db7536f2906d1de5ff488a0d7b4f767060db4e41f25cb28e348a8149c08c0e0bbd077d732e5616921f21d5558c09a2589515ccb65d5c836ad240f22aa0714ecd1b6bc7e25c08534a616086f9d671138ebbdc40182d3bce72d11fc5caef471d46e915612270ebbbb1c37f0ea542f822229746ee3fafac86c6efb4437a90b112deb27195b6bd244894a15c1a39777285efe4036b031f83614d01ca3e78167c103aa03f3e0869949ed8e6c2903052758eb9fd05df80b84cc8d4a19e895b32942ace012657c44eddee073feadfefff8e57dfd0f06629336f97ae38e39b89ce7e581e116ff8c40e5ca9a09e92659cbe1a29aaee870083662f836aa94a316cc70dd7fbd9719f6ed931876936ef0373dc9a99340d42c9b4ea8fab126f2c59b27f0dfdc181608f5aa4a96de990ca11b7f2837945c7680300374b72a5aeb08d197c2adbc27d6136579d1a7e754a5152e46a7c02f2887e074e724c9c7021c4bf175d8d3794c65fa75296cbb75f3bd26661e5766a23eb4e6e8841cdd64751d76da8fc873313e3dcf4748651a00139ba462f448c9486896258e6ab2bc00726bd00e11267e5b4db3ffec69ac8bb421453d6fa0188633ed13b19260b07b2469e70b2bf7e18219d54ef641a9c8326b58d0a016e3214f49ea3a0db4ba6273652da6408715902c6ece13cfb4e1c664ca097257fca2ad0bd7f41d32224db126f73c487e0d55e5140f10504de38810c05c37ff5797585be5b1d2db27b204263fc239f146d4e635a4344c44e9cafcda0dddd38566d647cbe9a7a25887812a66c47511c2c66371d201b20216683463617add455fee19e4666183e33e91019803d94a50cf94309bec3d11ffb1322a89124bd441f7d05219f9dd8671ae2160be983ce2752ccd2deed9fb124066a25e42efb0ddace1e0f6db764074660792ef9445675d15a8825edf7c321a8d3e9d9d0e0556dec1ba6bfafc70c1a0e9b645b8ba841b96aa9ccbd32cb6caa8dc95c05bef017a48c99ec569b8ac41906aece908f37ef1541c4b0864c2f15780a2d4ec01efb605c9991d30f7c0969b5293c508bfeee27a2080b60a9a2226e2d34f1de1cfe80752d1787e7d4d94ec0103679e318f7dffe143d3e79d8b881a4eb95f03665cd351b4ab0d5772de576a5b2807c080b13aa1123daa41e45abe312e1eeaad13bd5d30dfc9f46bcccec248a189b923667ad809b9c196a0bdd944f6194650c4232;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9b3180d7487e5dbdb5ba20a2728f89a3e4ec58b986833ff79fcc9518ad0fd739b1c20fe17401bdd82e5e34ba123cc54b2b7c0d24aee0a34ad9b548871546a5826e4d77585e182600191befa9b2991594192e5f8f31f55a036b6674809d48c7f9669545455474b3b8ecf01b2bf82034609a7d3aefee9c629eb233c58a03d531dd4834f0b7bcc9dc606cfea253647ec2afd04f1099c0bb2374f4a569725b4e454726304c5d6ced93835ac5c43687796fc7a72cceb4ee662cfda6410cfa640a3a70f9d8fe89fc2af6c72fb057036832f98b81de1752eedb3f93950d15334c04618f85bc34d7c79811e41848fc1f34e48a80a38bb760a800692e091a6dfb4cac5ff1736f28f19353ef2dcd87f6e2ccead21efa2dd43051b30a6546e4223977ebd3bb101e12c36e5cb0dc2e24f1b1c62aab34518c3466d721d7d6908f24dc89657eea6a809bf182a29e9dcffefa5d10e64f3a3ea0613dfad0eecacf44c9e95dc4703badb2927665b1e6e287b5896512cbab0c6cb60e9e3a5a074e9eabe2026c45f4c6bb021be6d7f100011149a80b4e0edd408268fca37ae8d2af4af24e19d4f29702f0a31d399f02d614cbd3fbe1ebdfecafa107f2d190bad94349cacac2cbf281c1dc54e7f62aca8b21cddd1a4b1fb165e9f4965e4545ea306ebfa33f86aa96d3a84012a9e3adcb754c6f6e9afbc502792594758ce8e80d95280503766b03ed840f4cc046ba552d9226310a27023f7c9d614b19a135f1b76cd726060e477db1afc1cdfbae0d70203e77ca1541c14639923ea3521a6cef1ad2d6238e2f1d3a0f6e2a330f0ee4c55dc1902461063a0623c98b5749c9c61f3bf25a9abce383ad72ddc18702f20baea3a34ca9de1ccc82b802a79dc99a9b5ec9277e4cff8927661d325d4cd8a876414b595838cbfaae7c2a5cfe5eef78a46d84ce524bccc1e3a6b4a2e6208e0b728b6b8b3d040d41464f99caba654a62699c2c2f2dd1f284a68f2b87145f9023880da72a60a1eee9fc0ec5c3a0882d3827a51cf6e3b63e4e0fc74547a455d45a3715f092d480adb1855b5d2723275749248e419e85a7da4c7006baff0d702561027491e4a92aea7bd0ef56805c7a449fed9ed018920453a46dd5dfa7f5c50da4233e02693c99f716af47afeff4a7ee6d564ff28bc104835581ad5b1c6310b2f822158e9718f5b732658c893de6216a89af4a773b7de9ed53c83362bbebc894ba20aa95c77941edae821f815902952141aebd9c8b8940725f74195a7da99a7c5cd573899feee27ddbf99d24763e203dcab279050b6355adc7f1be13cafc42b5bef1fe6aadc28f68f1a625970c560d8222a929ba300497d77e3651a775f3a0dbcef4d46633a8720e67ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb03e7960378009f3dbf96bddeeda157c3f89b5a2160228144ade6efd5dc0e3bf096b9c13cfd63f070a1deffbab7b31240346f10e5436e374e837fd26f59289623eb79628ec726186eb1c62aeeec87ab81649ed89f092d6f5d425b643387e2a6c3512688175f7902929c65a847d0746fa74b150ffc73fbb2c49405d69bba3873adff69ad908d95aadb0a1fe403fe684da160237a231941812f0f1df8f856d4c0522bf88fe212b3caa8cf15d8fecb0a455c4d16d191c3f78b74e9ecd81e230d862ce935a5f81f3348c0cdd24e0456cd0a50190bb578808ea9f39252f6f746d85d2a9f744fba5f4db1c5ba9777ccba28d90490c19b05b30a666e5f2306482b9eb7a6f05a893e476e260164cad1bf28c777eaf44d05a823b795ae4c250a821bc3342801980e49a8cabe910cc4e81061c6d6f8f716f14e4bcf1919a79d32b91af57b4dad2876bbe9aa21984f3c0d70950b30e4d0e0328d6dcd61f38f45bd538043e0bcb4b90ebc174181294c98e9511c093846ce334452cf8c2b76859afbf08be13da3910085350e9b81d7552ce640baa6f094a2a30843e239c9a5b692f25906dd6a2628ecfde06ecffa242f099f88935db3d9ec9caab82395310fc6fa90985b56b6d3a81c15f815bb90f7ab184100bbaf976f9506d02998fc527f55c382c942c6918d62ad0f90d36280b745cab2c0a98e54bf4e9d69445ef0bd4392bf25c78708353a2e4996f9ebaad3285b7d0b8b5a675bfcd8444c1d709a7604fddf026d54eb74acaf2a706ed593bb6e1a1096c276be6737e2f1c3721d55e835e783b5f2ce05dc8ac54c07d307d9a878abd9aff47c4960e10b6f061a506f57a0e14f8764540ced08297bf2e84887eba4eaa714c10d082a6006f6d0f84832183bd82b19f6748021b0f82405247ea3336000ce284111a2f5146896b9a349d063cb67d2ca09822fc8989c4ba083009524c40f2f023c20a5738d9b3e7cb2e01513000728c651ab79f00acb34a0fc9cfe3b4e884ea41df50f73276659fb165b30aadb8cd58201eea08e7e2ffc0101a03a9899d1da406ccb2312499344c4c757f4a41e06de03a7f8a0bc74a0f79aa952d29f961de50ac24d84cf33ec8450fcd9861418ee48d45b4f18faab3865e24c9ffc085bb028c03dcbc4fab6926eea28faad5905bddb9ecfcd149df3b5834661f9925b351dc143c3dd45f11ecc94e902eb3e5f0dd98a3e9b8edef775b075f164c5970ca90fdcf4e5f9c5c833decb32f710d26e668e6c7afa1f952341a418f20ebf3fd0864867fea9e222cb617dd8167e4b302701ac1b56b01c7b8b1e98cdcc62fd6f94a04fa9fc1185dd7713f5e16fa4f1080b98ff43e6f40388bf4d524c454ad5865ef2debb0cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5aef3bea56157e545e2f05d0da5c839e9fdc2d893f6ce7f452f633d143b81e7532750163c4c6daede1f89bd01b3969c2a171362677515fc49eb6c8e8955e3d90ca4405ac3115de3a6b0a3fcc86037f99c75b47352c22a601f3586d303683f869c8bcd404d9761cde488caab31255a025aa831794e99286d1f2d00dc5afe28f87b46784a3f35732def699ac193bfa2c520833228d58cffd4670b7e7c7a4e97b6ba5220cdbb394f60564f26483dbcf963a178d8e3c9b356fd0651c0958072ae65031581d5965cc9bf67e88b651d545b57185137e88c8f2779dc2c00a5272a0f9db3dd0887dec65c17c903345da4055831012ea4403d4cac7d61cdc1731906c977b3e94a2d20b957a0e69cf320aaa2c29d0799bdb3d65077563c8a54f1041872ed208cda523ed45ae4e086c70178ea5bb921c177780fd611f51b688036152458c91b05f6f88e665bd424a1fae2f7c50cdb3a7c9c234d5c644c7f7e17dc85481b6af20dbf483e54933cb951055057fc517ec48b4c8ee79fe61ecf71f17508f9a5d7fc2422e389d985e583e04b3c89a1ba9755e87941508950c81e1a817ad1f9b0fa6bc18d63ec3491bca228e7be939e132e161fa5c44b76745ea792c0a99d1c3f98fff9d1c3cf3edecba6c95ee701c605e7b1bafb2290cec26d8f30fbfc0e3ae029a28fc7661fdc2e047f7e63c59708be465b5f41e20390d2699ed6f29815dbc39d5f3bbf4ebad4e4966774424928ed4aec35846a9ce373b190408569b34dc25b6900b9da778bed464b70423b28ad36e6626d7cbe0708662b5b25a914194319545f7576ad9c049d750cc09cb4ae85d98f591c5e79f34980cce4604cc14270161b367fd327b076d57955edb29a46ca3fcf666ff9da9e35d8bbca54647ab20bc6ddb2ef87ee536a0efc9e2d7f593b30ebdad9b48123e47eb18b77248b0e8fb9971d2addd91b468d57115f21f6b51ff5fad051cfdbd35abdea1a2e1b638658cb4fd47bcf4b232254726d3d9230bdbd2178b4cca268eb8b82fe2d3afabcc2a1f3a2d89999b8e7749f3913f84f05771f0b4efdb8345e62c525d346ab56b34760581521ad0f303c2002c6c6d598c0058a3efe60c57ecbf2d8272e5cc79666afc5f40b936a13157789a81e55ef7a1c43f0418580f9f5c5adfae7937c030f46a0da94a6b9973ee8098609ec291c27268875b04af840d5b9be867090fbd86a2424f35ad8c92676bb93dfa6de0edfffccbc192143a46d31173c71256a33fa3c0ab8f0b828d42e7daed917ed8d2cdb095a9d52504bf109a3b567083bc58b78d95b0064c33848d3a46adceac2ad81563bd1e01d4e396c259b23b7346c21a7d17f2fb7b41c01657466cca912191e78e7d2e536c7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hbfdcdf88b1c1925aacfe021d67b9914aed2abd4c142bd9cdeeb6229d955e0ee93f254fa245d7c6edf9f161554cd64fa7dce38a9875fed156ab78a3b4fa796398b33a1e4a537933a5129d8e57c29bbef7da99591db63278d5c4c480a41feebdc18474d0332492cab20690aff88ad92963c438337a7e05e3bb29f111982288a06942a2689f43593353b4c99f49b0af164567fb33cd98c71c010fe1c793905c754f09cb73f51e7aa1af0dc34c83031cf2e41cad1dc85ea95717009bf095c8326c5b572f7862c0e0af8038d649bd2693f7da1b7bf8f7efb2802aebe53564784f6d3dde6c1acec18a8ba415a38beb1bf620415cbc289d0e81c43ebd80f247769a44379c43fc57a8478b4a254ae9285d495b3c472e1beb0e90a29ee6ec2c114f64f776e589257f48115a706b2af643e1786dfdeb83dde067527932dce7d1de8bd722303977e5febd7ea3f6a54b543185b05ac507ac40a34eab73e8073d44d91dfac1fd27fbb467300946be1f609106e059e6299eabda1c61b2a808a097a6563eb03469d1feec477c0e9ab9bbda0e203ba8eda45f48e2b50392f6b472a08255f9cbc08bdc3b8ed9abbf2dd92a88ad5b5665a5538cdb7fe4eb2cbb8b0d6d60d29cbf2eaacfccbeafd07287425ee441d5ad61ad96a17bc1fa23027c27f04e967899f335053eb8b4ad22b90d366c47d49f7314af72031836362cca7a999e455dba198b56c72d1d3573dff336cf25ee1d752af01412e5bfc0ad3d3136689cbc62fcf82ed65f30c970338d4a46083a2cc6252909ee1ce1553c548ba40ccd63345a11e7b68f5e5bb3d08645f529b778eb5eb49c5870c76621e89f6fff9a8d46b78cfc87e54c13e295ff96cf7e34b6b66fecf0f3bfba3b43b92d5d83be6cc4092dc7fdfd7719cde3ead4ae4ab1a3bf310d3e6f57fb279de6fd26623d7ee31457ab3554fdd60c5002e2f66553e38fffbac4a48b8991399ef5ee672c4153f062bbcce812121975e5460fe6d67271f77674004ca9eca77b500ec5eb770fdf41f00606fc754cbfda559f6d92e0a24d99a6ebb395cda342ce281f8e5be5ef7f5e099ec19c0c1da9382d430c8e8d4ca228eb09ebc092ae16f79d58fb3a1eecab32a85de727b5b5415d35db09fad15ea9ab64b7baab25657890f69756a7e827075830467295ad7307bb592f89e0eb18db670c7e7b4dc46768bc8c517935ca1b247f9adb5483b6f17856f968b9ab2220f2d1ad235c2a9df8bae0ef3e084320dc9cc454f005570bd674dc73d45a5145560c46b6ba57209ac4c297bee3abe699eb9688936faae02e15156c44f019ac75baadb4a0bdd5aa6f774541d427b2785dfdf7f5a9dfb7ed067519546c082ff434fec27b6006e2326a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8ba3ad2674dde391cb5f647b77a59184333fecf3ae52e446640f066681adbc4befd05f78756fe6646bdee9c92f698d48825230693f5eb45ff7d09ad77d83a26a329c1318d8ad046eec8c281c0fd1a2958b92c98dd84f049459bcd88ea7fea407a11f186ed24eaefe0c47441f11931d8842f54f839cbfa204c23c001c61edb41c29cfacba380c8b0655c339ac3a785944546462deae65550151e27b037306d0b1f25da334750e3aa6f76b1523878562dc8a5221d3fab8a01dfca2e6e19df1987b2447871c78722634e49ec2eb2488677b3c5a81db74b620351e657448dffb9a556cbb44917741898738349f368e4a6b203d38bcb33dbb3831b5aec75ba2edd5078f5cbee74170a3549b7fb29cfe5fc1d683d240ee97e58cbcccc39004b9a453f2ae79148e58647c794699982822246d117c3341cad3709e0b55eea832ad6ab7686cdf3656b7f63fac117f611c7b2016f1b0f9232f2373c6fdd59815d01f67c82fa26f0297bc0a05f9b11e76c69dfbda4d76507c5aa8cd157ab3d81a1a693572dabe98a7a0900c96ea204c89ead521086cffe458352b25db400776ec95925c4a49a6fda88197b0201eecb3deaf7450deff62bdc8aa8171c3f0c820aa06d85dd1783452ddf721eb508d98df38f425c0bb37b0e94695dc51c990712b384dd45389756bc9c16f7f57b6825bc55b3f2643b91db6d4e6ca69ce2ba346c9e6d205e88958afcadbcc35df4234c8730fa5b69a5829df38bb948dd97f150e589bffa5026bebd2c40d728271784556edf2159e00c1db521e950f787f9e64e97a874f18870e4a22973e855226db919049beb6d2b67965b088f2aa166b99d4feb714eb438d9680ddc02bdf593c4c98b98275a8e1a3d32116670b2c189196570ce93a444cbfb71590474d63ebdc01b511632ee2899bea6255bf1b534d5099bfbf97bcde1fc1fda03cfd5b89b9f11f8acfc4de32f5cd2c19e665128203de2c2a30cf5b8cbecc45d0a223eda9698b7adafe92d2042c124771c14464370a18f68d9acdf0f99a7907dd5a1eed06d2c47812e17c0f411a52218171b58b624d5ce126da1dc0f1597f7d11b389cc18f955de5b5243c6ba0bf9384ff566a09d99a319d3ff6e867a3896466bf7c13a9977eb28922336e3856f65a5d8471d067c4254fd70940288b6b20b9c28ba3bbb0ffbfda77ad45b54b11c6be750905768ce71beca4b43c0573f1d1cfa887ae221730a5f9f6a3fd14a997fb7068bcd90e329f626cd2c5d5b30453b660b537fd5832004ed5df4a0bb6156199c3dca1b24b36652b1f1642ff0ca4636c60a224be07f6a5549c16c408d4d2443c723e48746215bb0c1a6a244f51668c8dd882bcebcc0254554ff06f2663b7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf34509de39507e3024fd88117f91bf574a7872ec7dfb0a3030b8b7069d9bc45ffcb4390a66d56ce97de4b0c9eb895a172d0583fc36a41dec5381bd9a26d600d4bae5f81618b946a1417d6f19f7f3fcf828c299012408dffe09466b7ccea9305b145b123927d23f89f61b4cd877f2e12c7d9d050cfe9a906e0422af21fea110d5971ac19ac5b36933b399fa3bb7cefa286afbd854bfe2e69ee9982e121bfcea25224e2d3ef78060953a6f377286178311b6623ce5eb0bee84778be9678dca1d6cca6edd41441902074e9efd38a5f322883340a7b81ba3210c2d41bb2f541b8ec401f05c1d96c763048452f458611ddbd0956c33f87303183c190e4404792607d2f762caa351cf1f7454be649b4dbc6831deb57b85cbd404b18a383424135a5f71481f3ff28999e33d35ed7829abb3c7ebd2d419efe9f992a54202fb1d8955fa0c590b2fe5642efec5fc3382fe99894cad3acc79f1b555c8192b4b9112691b409c432976cf41cad5d880fa59e30dd34de63b6fd2131f076c01c239193e0f3f02fe2be57164c253b719f3e2302791291ee58160cd28f410e7ab8beaf5fb4d4e3430398245eb7193a210c5373c8660770a1d387b3adf69db3e476c47f3cd5d657da44ffa963b4aecd83ea955b2568b0e36eb0aee9289c0a11a58794a40176513e6911a46b7cf1f89e545567a8b710165f9efe83f16e75d0e2a4ddb993a371f7866a874ae092c8dffddc87de1cc2aa92ffc4b33d1ef2ea435a7fc16422a160edbb0d6fc1053cf87d0e653e5b4b7ee5c997b535bda3797084ad8b698d4122e49d100e9a0ebf1e63d7e93f1e732e797c4ebd6766e3fc7e55db3b77c1c58242d754f7e03c573f76f7c676622ea10cf439a7c35a867d6e5456eacb1fe008e76cdc5b1cfb9a3a617745b1f22fa9624c6f24294488f7edf7721953e4d64037db0f25b332f4206c3b98d0fe06c0e03ae093ad221681347cf477bcd3274d3fa460a8f232f88416e48001f4dcda25805f02623006d48f4cee75563256cac294ad8f42efe0f0ff5239245ecb184cb575cb12f2988f9f007c31865c7400c86091ceb65f3ff3f7b482eb9c1101fedb27e580ed61a4c5919bd8ea8d9177837d0e7943b595b1820aead10a532fc7c8c77f9e2bc353ebdc1e3978cbe9dd19cfcd02cbf1026a10305d35c73da579f7e4cfc1a6c28942c4f8b46bf678ac06f5623d42eafb1da4c9d26915491fc84d450d55cfcad550e9da527e6cca906848bddd43360a5171dc68dfe69b6adea6937699ac77cae859197c711e8dfaf063e7766716806eb49df733ebf1b6e1fd3ee20d5cdf8891d553ff40726043835c3b50469868d7fe90326bc25f2f0a154fae32ae9c82ac649e94e6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h96fcab16c412b3c886f9e7bc66f1b699fff185893e4ee174d54ba030d7ac24eaf1d626d7120bdc01856526658d79f9a9fd07c722e264662fa5809f56add6138cea3c235a39b3ced6c5e99dcc8a9ab606319bab96b6d9d51d18023130ed8977ea797ca0f37add9d0bae7367603de80487fb0cc39150030d1083c0e521d85595d6483c9303e18bd75ad1c699dba2c030d74167b3570cadad388488ad455e21e9b07b5b514da62758ab4cdf4d7cd2d46aa7de71490fb3f7fbae218f04f9622e02376ee3476db3cc7f77d4415a7f4377086b579d89dca6d17245be5fd327431ab179272df033fe012c16151503386018f66b409ef23c0da84197dd20142cc5fb9a5096272d175cb2561a533018b4054ce05c4246b2b917f2c6122fdda95aa8f3dbd0707c425ebf60af9879f8c6aa542cb7ea0ef6042f670cd280ef9a9c2a62e48f321e0f4c91c8ec6117fbce9ef9c469d702dcbf5a9637bd4bf71d5d4c6885f1b3ab03dabef6b52d837310c92d972888c4c7fbf74fa68ca6674048ed6a782b4603e6bdff5076ee9d8cf103cef7993be702501e68f3606975a0430de5cd71d360c0f0be2fe7c6f446afb04b2bc14fb177f9ab236fbb94dbc3ec4fb9bd13b82838772e145f1da10867b51eaf72535b69fc3995905d45ffef36be8ed458278773792c4461cc9290a6416b33ba0a6c061e016fdbf88d77c373c447b40fbea366d63b9eb49dfe2afcbd09d72275ffb14a0ae5c257d91e1311c906834aae066aad6ec8e0d46348025806d0aa6f79724449a5e3b7da2c8b9722152a1ba3662a5c71fa5033e935e551624e0ca9c9ce6f380f9ee0989d5cccb10542f017414515b12f1b4c8dbde664a7df74a77e6f42f2547ea65a9b90c05706cefefe78fae2677a1fc64877b8e9a54819f8e270b9a2adf149453af48c30f77d2d2e0e127208a808cee41e368b90c7ba0d977db85db4498ad10a38d200e67aba2ebdaddf2702a885a6ad818abe1be7d2704d4d6d09602c3731937ebb641771ade2741aca48b555caddef3c0f3c335ff7d71e83c008d8ecaf249118944072e5c406c071b9a275ac99d10f7ac8860333a5548ebc6547603b34bb5ef5c798e5d98e62f01805b39e10016ff434592fe6af51c16e920a89ff4e3252920365eb7ae4fcd05bfec54d0908a81259a4a31deb5bf66a377a8091ecdebef6d46c6e61a391f78caa46abd0b8acacba1519e6490e102be81d2f42f892fd00e61833ea7bda8e83a89154c70fa2a58b1a855e3d5b6a614d5061051568cfb2960b59aecc3b80ff511f89df1b2f3ef6325086b210a363339edb787a1a6747923e28ea8c7946c266a4bde6968c07620e9999c654be19b016514f01f5624398ae638f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'heffd62bdaedbeffd939c1b29bab5f70341413edeab44f2201bb78f3ca515f2de597d5da01f005656bfade6b95c47808124ea01620018bcd0591e5fa5a2ec25e6118c1f1119a5895ed17ae1a00f61ee759549546d4779b28899bce96132fc0ccb52471f89f06559bd7508ae49c6cbc5ba06035103ce68fc1ac44f73b0f69bfb034c1616fecd5d23aee539782e697edbfc48311776fff4b587727599162d12d4a868c0e15a34d833ee18a4e28acffdee98c8999901408f222115c191e6057db27bdd9d8ad06f12f724fbdc0359d92ccf2f094f51a10fc7080a0b0a552ab9a5c9478376d55f7b862ba7e705fa481e1d47ea271337785be0b469af0df549151260d9e7f61000c63578cd8c252f0a5401193a9e18fd8edd7b75fdd78ae71727a4a886b6af2e08b2ea35544f916e04206231c1a1654378e64233a938da6ca538fd89c230cc2378d8a7fe996e506779198500def8a7be3cab475f4360c0d6c76c22532d1aa8106927e7849cea2a3cc44bca2e62b809f75150e7a1aadd98e37bc3cd9388af7f8f5b236c522bba324bcc39d25d90b3fce669a3f81233d625a0177e785a627b48543ee588890be1d2491cd874142100bbac89380c841fea808ab250653004c8c2e79ee008befb933e9df78b2f157c74115938ddfc3c1f449591dc619e38fee4916036c33de4d51e9a792c3c1a81f7661165cb14db81a714ee7e03bd50fca009ef0b90b68a10ccadf91f4e3acdfeabb484d3736da198d7eb4299ed1c88f89c6391b75f50502b022f9e6ea0b6a11078c54eb3f6a6b5076349dad0dcd96f68fccd97723bf14be8244903d7130d36b842ecca6c785e0fbc0a49c9f0839093a1bc08c9d85787ec4e8f6fac4b934e26b29e79c99a5f42ed5a9feda9190ab225ceb47b893e2cde6766368bf3a70d4fb2fd870d3f010b6fa17ee7a2b1540216124b018e9f0cc2912d6cd5ee0432f0ab23aba0d5b81a2c180237a65e5561da5f0ad5d7a956d1196f7a12f3b096bdcf4e563cebbf6cae0a5cc078d3a939729b4b9d2363c82caac4cae3eea9a3cf75dc81406254bd2bf2e10f8b800893e4039b0b6f25aedda9e75add465db0c9493ae7e28c7f306d151d13127bebab2537d456839faec100ac62580df5f35071aa1e2242c671760b8c8b745a2036b97a46c0e002b297b9231a8240e2b5b78dca78c5a88166072c0d8ab836e77d3e87f5e113be7ff63a7aed10032f00a5372a44e3be4d607d01b92d86e2348d0707c32893bd94f147af899aa391c8455f4c3ba8bbfb10e3677633fde51be0e0c83f3cadd352a6dd52e3725573b2412fb58df524f4c6c01c88641acf4567d49f9f6c660f7c121e4ab6d97e8079d712c0c5e294118e073b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4e9cfbff2f922beaec6e81c90de1abe70e72235e2e011fda86792b83eb29764ca5c214d667c983eb4906fc2126c1ab702a732a7f5d24af698425b1a1442e45be4a0adfeb42a41748a1590c3e2e0d26accfe6679ddf1143aefbb2b4ffff6d36c97df63a3a7ebbf16936cb7b2440b94d0da28568196f923a7dd1260d6ec079458e6758724d8e48fafeccdec7089781a676b5ab5c4984e87dddcd9e79173fc1c3786dfe6b2d33b338b9559ddb6e10cf396c2ebafcbb11d48d69499ce7c026edd8dcd469f506790ba639df0379a4c0a78d4fed93a344621cfc62850cd72f606026074219fec6685a82f98539d1ab0d89a992e1ae245e7ac7fe553b3bb81f49a98d49e03fb1ba418fd428475549aa26d97298117af006f215260313f40a5ff037ff84f652dd005ecbfc27a057ff7d047d057f197d370fb47e715e77738fada25fb3155e6837095862e79aab5e8d8e914f8e3c89ffe5bea1381d4a493aa0893f9c400bb488834bf8bfe668657aee641a89707128949f9db41d63ff1123c6dd460234a52eea2049fd372384ff06c90d392a144141f26e7136aa1be49f4bb5583123c6b21484be8bcfee9e5451dff0c4fd4ba787df9e87a495bf56041e740e5f9ab36db04afe4d98f50c4a9a019e70f3c91a8254918566a2ec3dcb64b8e11b40c73d1df5d64ed7a8dbac364e876ee979cc1dbb2c8c8adab259ae63d2f85b89466ec884e3f0ec46c3e7ee8b3e83c8cb3ff4efa3fc33a1a39411ba3780b9afd78499a9d2a417350dc6f6cc617e2794ce8a3188fd5976eaf335bba6c78bff261bab6c7a9a9524e2daf6b8258c978f347d30059d2b3e873d9563ffa3dc5e23efd7d637d51c356b186676c1e384961c36c21369382b6275fdf18de293188f1f0dff4ecdf9ae7aa9e39ed2751268d24c24b5c4115c828bca89b443c636aab0fda2fbe42c5999fa83904ea6419e32c4855a13002c89b6d318432704a632ab902367416abf6db2c5ade80fb79c4d9f2a1fb55d3818ea47297cc1a8800f70cb3738144d7334c379c543fa32390154e8cd7f1084ddf057bf93171c4b328e08f5339a1dde8ea1689e099dcf20c77e4fc5040776c933d97f04d7eabd68a93b166b65ec77ef18655c43fc46a950f413f9cb149ef355cb2230a2d1680c8eaec314b96b545e1527b0fff098f2cc2ede4ee329ca407890fc5f3a069d1a57ea5aaaa55895c115aa34bbaf1af5072df2f2ab68df29a997095015e5566eedbaa199563083d189aa2f64c6750a2e941ccfa3862cc486b044a2b15e83dbcb24dbd1b44940a9af8a40570ca3ce3aa9c3793fcd2cd9c35673c02e4bda6aa58b06e2c42551fd62f35fd680b662a7dbd192b8175cf6ef26e464c48531;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1edec73da615b6a61cbc909c0edfa56426ba2686f7c1b981b6df96f8efcacb3b644c92b6c7c8517aa264dcae6d608e6e0f61d208d6c9075bbd516d74c194357c12d11dd088467ab5fbc33ecd8b7aeea4d066fd419c679d3b7f565be1296aab3ba0ec923417ad229c9e6c47f5b973927e0150923e8759e5bcb8c842c4b28357ede392f8e27e9179ff8263d06a60848b771e79de81b7a365b6f313b35e2e215bd95c7c1f3dfbcbad0c9c6f4b06bfeeecdfb25dcd4f43864a0cba8fe2d7c87df00a2f557ed9e9884876cced95a514ebaad827bff53c6f12412cbfff8eebc55a3d6294194a1b1380722ba31ec9ad25e5d79fc8c018de325ab309e21c3647071a842c91ce54a27818b232abbb83a719b444fb174a839d8ba0172365a236400356e95fc717025e6a9c08a367a10c1ba7c6486509c8ec415805abf0183ad3aee76d0e2c39f3ee19dc7bbd36a29bc37a74195db8c7e1a2f37f2f93357a3ff9ca210e97f90142a114391e9789c3e77cf5e112406b434cdd91c59fece5bcb4eec437efb0340b930f7b4f513cbd8dbb721e58013c9775851765847898ed05c16e84c3ea76958e59f21923b7c6b82594476777bf4fccccf2292dcb1780388bb1821cb179893612f20eba24d447e300d0e6518456527a4d70f2ff77d63239bc2efb8a2be56a54128c94450475babd3441a75d373ebca2d3cf30c25f5faa0b4e4d6364e46ac5b2131b4f0dd33faf2e55fc5add77f19cc8ed38428957de73f9406f455c6d81d8ea4729b7daaf31b90c5044b9c3df6c313e36a6559332e9ca6ebe25525cfcb9ad61b6b8f7a67ea53d9138a4720293dff0f7991917bc2de6181a7e7a006730442a357eea26cffed9f7618eaea771a201da2f05056fd993febeeebebe99c98540982265cfb5c42127a2db7c24f9823d74c8ecae5405bc8125829aa0f02f6eece35943c50dce3fbda3427178182dc5541f1966839932ca437c880439bb7a221129032b590376c8500059544a885f69b7230ad4393eab9db56ad30d3cbc9b4148ab0e6e2f70f76ad7d562dab40c2d22720474915843d04b228517b605cc84161b0c6cc598ab9f4de447855184b0c792ec1d2c5d8cce85f3259815ed13fd228c81e52c8ab00a8bac702d5fbedc3f75444b04bf04ac0b4386d902a6bfaa02fbe5374358b39ab7ba201ddc2dae074106eeb65f48a48cda3b0bb7d8ac386fed46760fb970add3fb634df40ae856397375b11a3c7da3939c51187a1c224471fe073bc08dad6cfbefe69554248250d54b29abadd4f5516cdd20d1fae1962d1de36e95bd85c15d966fd76d23614aef1791ff9c4f264d20ea7042739abcf31e5f52659548b96292f5d92980d4d23e064d5f45d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h90496cdb8b04bf86e1d7998b0b554bb065a7c0734564e44cd3fc90ff57334fa19b783fab305d90c8aa57ace3d0fa74c8021d5f3b3582cd973dfc9f50b4f4e9830e56b03e99fbef1a5ef268ffe662a4afa8a16316e6dad58883fa56cfc3068bd0ceaa112899ebb38ab13c3de064c6e3393b7283c2231d615de2184a1dd961322d9375990e74516a714009c583befc0a2d8fd4cf4a6df008d18b64a86f0da9e946b056f4668dceab59d930522efe0e0953a8eafeab129a91fde08500af71f32371153654906095f431a1548275fb90bf12b1e999db58cdc3825be4d555c8a082090787b42b3744fafac19178a74afc78486f0b4a949c61684bbc2d31e5dba434a00f75715c9bdce75c0d7d407439655dae0e32a8f4fbcd7aadbba404c92e2d9e31549852ebd075e1482037ec95452924f99f704ed31fc1d019ff259a35a0e386dd998664507b90472a4d65e8b527e93318ebd5e7d9b8a223cf331f9157c06d1983a3fdd6cd1a0444b3f6b077ed975b9c50a7ba7471f855faaeae557be2986a9a937b0fbf7dd8663018659de1f751b1d5a355fdc60158e8b3b8b7d2fb9cb98c953cba44ff434637355c251737ce3aaaf2cd32bb2f0169f32e5975763e66ea69456d3bc7911ba1a811744a0dcac9e6b60153a4dab1402623e622dcf58755c8f5a96621351b469af21ace24eaba3c778619cac6e5ba0678926a14702b91e378832ef286fdb676821c19d492ae474192d996a525b76dab5653c82a43aa5fc88613cfcc71fbf70fec2abc17dc4cef0a1f290ba951cec1ea3e7876ae8d0bb49d125070494d202e4ea79cad10907321066aa339b12016e939af4abcd984bee79350840c255a8a95d9f6c1c24c817fed73931ed4791cb7986c70da02965986fbe9766dd5792743f829c27a2b4bb68ab763ba14b14f0a0fa094480b0687016fab4f86b262d97fb8bf86002c4ff4e80caf1a10d2af2e0a61072070920a602d90b78c5dd12cfae14e140c2db135ecbc624ffa5df8170fc49096ac0e7b2e9265e225aa6c86d707e6b3ae08916a56d2e6ad5b3a3073f01c3b9b211b9259f4d4fe795620962abf38398a573b30c7eadeac2630bdce4a88fe95d7a5e3d2f0ea4a7be448d840019fbe171ada8d0d54dc1fbe4cd273b4a8bedcffb377aa724e09159fda56425d6ea1982e634a1937ea71888aec4d11f2f2699c14e01feef3f29e19adc9c5e4182c0d8b0fa489e74d43fa4f648148eecdb410c524957268c2c019f694941cd3c7680ef393a5c30fe0858c63a355a6405f0745415a091225d23cf77fd9c3f193f52a4dbd572f0862b37d6d4b2e641f5367e08141463b762af05e962d483f9c8dc3c2a8a2ee401b460f376bfe734e21b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hfa2cf1cbc02e3435ba75c47599497f9c9f24927630ab4a509dc4af5b481f72831bf2cfb03503451db776243609aa55af70bee74bb40fcf3a32248ed6ea76ffa63ab4c1d71672953070436e5fb029ce5ca2f3a894ced679c16ab6250beaa551f3aa9dec4088da2283cf84fa5507b12e3e89dd26f585c21b318b9c7689f7f100cc0a680a7a2d0d505121f4dc02af5f40caebb50f69a107c7bc2cb8ac2419c37c96a6d8f797930dee4a4a926ef5649fbac0e8010358a06415d856f8c2607240020c04fc0f17822873ac82bfa7eb5cba9f884110d405c5f3b519bfa386cc4d406f499e7050bdfa82131e16e7fc47b505fe90755e95ae364b7edca9530b12458d2bea06a8ce7709386264335e16287c6a8879b028d7254e2b8eb3213b981bf60d138a4d58c360f5ecacadde536b86295b772e688bc01f0dc97bab252a7b1f9c6fe98c26c8f397fdf9dfcd0a443b522d67ca28b308737f88cb60847df6b188740fd46f60675bea0a5bad001672c9a0777b08d724ea754c4894ba9f00f51c165befbc98eba006886a729e2e7ec189fb98548e20599812af08691733a21fb5112b38eb6432bd58647006fa11b6553fe366ce8a87608bdeeac6c410d6b981e819c0670abeb7276955acae156cf3257d51728a8953f2a43277c91b3091a6212da05356589286f1cacdba1753aa2f08be7f5e33aa16cc093bfb40ea604c3e2037f1a860c7f3e49a09c280e9d3acf91066ee82d70aa9beb79501305883bfc55f53d27a06a38e04d890da49c64caf0bfd311ee890ee63d44a8981910cff397fdb614e67c8127b20c9a3bd3a71907c20a8b0dbfbdcac4f11b666bbc8cc59215abd97cf45be595a1ec3245c0d290d6142f8280534e3d643176724e7bf1b14103da924403a6cc716126e465b7e5a008aeea377642d5ff1c9b0612d1a29545ca3e2ec149ad21d1f2adbc9ba009b7e067bce3debfbcd9fb3b6375a8205c0368f7f7f6180234a55c2d35efc29dd61849af933ee942fadc4e12f3493ccdd1d071bce2507395cfdf2ddf2cea218469c2949c42a92dcfe5625dd5579d4ab3eb3e2381f676963a082a353f7e4818c3cbbba319662f16ca613f882a79a489b71592e21ac1f69182a4b135d9f9ab0223c3b60496a4c1b76080a661ad299adf8849dac2666917774dc9bcad9609644cdae34abe471d78a285bc7062997735bddc5720d067c61bca450bde1cf6db81243baee6c76e95b78de1a0a951e042fbfb53fc119907a463d0e2e5c8e8e2e9a0d03515ea1b28f4de3a854548b3bea452456463fdacab73b9f89d018e0df75cf787e8985c7088d679d68820b20189fa0264d27c27fe87ed6556e1e73800a87d726dffa7e52b63c60593f68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5854ac0cd8c6880783a8bb18791324328acf207416c98b6fc8fb05a6a36c1b31a4acce4e45ee702e0acc76b662631b7617d44efa2962140a3bcffe1d7f0b00903744f29fe59df774063cabad25536671b4b84f17065d27d5f19492a1f73f17aa17a4e6706356ab430c2896087162c3bc96b248db8d4e3c807f139c6dbb007405c96dd0d1dd0d2b890a54ef9409898b7062224407bc026f8e4b4b4bb109b12f52f76afe3394290275296883fb34c5d23f21b2ac8f4155e452cb79c0f10e09270498c669bd836f71733f92da3e26fa3cf8ec6d7fdb1a73f19dccd352fb07315c6433571c99bed3066708357008d0af8e6cba628f5b9822a2bb86e4681f8874578a0186d2a48a6720add70a52b06fb8f29a895a063f1f665da64dc5c4742d0f54f65c258a47765a11bac46d7deae9796991fe19baa8408618c43eb0b221dc0429a90f6d49d2ffb4833b6a9bd61c03c359cebdded785fbe1d9b1534bcf237d26aa525e19b002003ca7e41897e838cd1aaae214a69cca291d7a26c038e36647e70abe131f3b737bdbdb974261e76ff8c9bcc333475cde5dcf3905ecc6198ae2887ed75824e5dea9b9c273571cb5dce2f0205070b292c5cc8fa8dec417853834b8bf610cb55e75ecea44e3931d74c61b431fd7bb1b9e65a9cc31f363fcc07be5fe18b9fd09928a188ff46bb845fb67a2b4c41f62afa8ee4379dd0f69c7b34323ef9941b82b33ba7f30b4f8e56c5f22aa78ab1ba0005eb81fc196468f1c6ab6dc69ae7a968f5e283663c3fc86732cf305a8471a5dcc63b5f2961b9370d5cf96f7eb0d0277d0ef6abaa7231b7f45120596e4d5e120e468b2942dfdd7d3224482978e880a241d28f982e0850625a713c16fcab7ef17e74c40265fe0df1f579da643b0259b4abfaf6e9886d7f6dc5cebfc76032a73ea6692c78048e3a57c6f8ab4e73f50c0c0c3a6ce3690d762b52d63c9042dfc710e730137dbba78c05261c89408fbbeeebd0aa93376f9dc215771b151eda2510b0a6bdbd6e197587bd31cf25a3fe3db72b84d8f7e78a6a59af59e2021a64fddf915e2624e0aa95e93151e3301bae5f00e760d61fb7995535298d116fc4b28ca8a4c01df41d2e86a9f5e670f85f5af49f8db48398372c7f72719a8d3242e4f5321e1cc902130e19372b4ce2e959ce13177e715fa3c28a725275e1e478e29bda6363fdbaf84108611f02476b2a8f4d7b5b73feb98d35061bb62767fa08a3a29aabd3c0096e1a29ead07bb47e0a043a44a67836a2a0141a1a2f4e292eaabdad446aa67ae7a59d59486e1e118d3a3564b13684ecbe9f1a7dc752beb03980a2923a58d471e5365f0d73fea021338edcb615b993ec1eab66272ffc38abda65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h82d7be3ea2df819aeb5b2682dd66218267f6a9c5c88f3d5cdad2b6b807e3c51fab489c6797009268760a145b75867cfc10d3148975b7a74050e087fadbadd81af431b0e3c458dbe4a1e7ce09912d2c69ed5568491fcc9e0cf2843a135887400d0ced0c6b977d6032c6190e3d18845012f16a473e2a2a0f81316630ce4dacb888f727404abde85a597d14e33e8b30ebf7ee63a64c1435a3975ddb46eb78f6b48359d16a622034afb0803f7ab8630947b725b16c5336b0b855d770dc36384644b1448430e9e035733c83d3c063832970c7e5f0b605650123358fc095fa9bc335b41a764b770431f50c93835f99da6f43f1a01513ecf75ac807697a21aa54ecb35dc76a8a24d08bc8b158bb041999fb1c85d2746245f03a7458c562fb2f75bc059130db0ec46ce12cd8e7ec905db53981435bfc0e2b21a07145c129a5cab586040d13b2675ead10a503526d3338cead7505cf252e21340250fa0e4efb4200ec10eeb754ce22449359a859e447b3c66810fc492e55e799458069422e55f43eb431b785047b3929ae2c2d6b5c8dbc421744f6dcd581d25e7dbd3a31b40e9820f2c04e0f7b341347644908cceb50efd63b15362662a745e4df7c45db6710f70b36de94214b4108ca5a73367597620108198fe2439068885fb8e73887864ea213975b7f298978bf7df270431fb126b55ecc02f2550430faabd04c32805596749e38099f57d3c3bca579b92e23734e918e91e0c892c437907e6f1ecb32933258f84eaf2edc5084f04239b19aa2131971dea4a3fb6a5204045dc248d82ba03331820d162d695fd393a699c65657776ee608d3f5c2fef8ecd7c3d5daabe46eb39e621a108dee82ddcf2d2f0db022e18e4b37ff12796763433cf5542cf6c420e27d24c68151eaf3613ab191ff0a342d6772eae539731168800587e48a77a0f96ab4b06bf89043645807f7855efa286ed4df7867e8b331635b7e276868b2a09afb12d38e65e02bd2ac25ad1ab9a32f6aa7a507b15c853f608f29df6e5b42f2a9efa723c82085cda32036fe5c0869afc6b74ccc9aefebc37c2785046f77dc064a58e9e93754d715a52cd9a5ffb71ad4d359f2983e3032f91132cd228274dd92b65c8adf679da1444c782f3b3e3ab1bdea2aa669718057cabe2609fa3991ea38e741a5534a863f8956bcfcf3dd9e8920971b75a8fc2598d1cb4ec97f539e48f5eb85fa295c3700d9b9ad8473ed0302e87539bdaf48db75d7950ef7c1a2a8b0669ce03b55a867574c02cae4e886829336ea6cbc69b7874f60234e2409816c726312f64419b60224940ee00d9f3162d1eaadf297e8f85136d7295f95ae68594d670e7652041ce32bec01f82e1797667e339a4734;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h93a0c3a04b293811a02d176b68276a3c35920980a8427db3a021082b66161f41534de57a175058af2cdfcb75501e87fd9770d5bf29e0cf0d3aed961cd651bfdd929a14826c8dade081391e859c99b0c63c07c5107def95a2db54e7670f0ab443d09de1bd49d47f8f6a87c2b7e7e52cae885b15b3ba40306c11143a573c895991ca030179e9e3f3f65ac2c21107066773e17527cbf8146061f91b5e354f031e73e85fc9ef6166bd3b7c78049793d7105de1f2b81d6df30f12ec9d79efc329aa7a2b6be70b78fe932c607725afa8608b2d912add2816ee1de3b5a3171589d3a5f5090eb4aa37b258841fb1b3d2e8eb30e733d691ac9e1eaa403052ca0a77836b74464f79319ced775a8ece05575c7bd251a31ef3f1de62e9631c5c31f9c421eccef49cf5a1263dd1fe7c4b32e9a587e90cab092cdfd8c8827e06023cfd3cf1c60c0400d94a76b9c08969f0308fa2f79bc300c7f056cbf40839453912861c795d193cff80d82c9910062884ba40f25db154153a15b1aa562f785f41cf234b5052cc1d8bad4e82911350245756635631c3089a02673313761aa4ed6dc3d56f5143ea58f5e5f3e06116a9b066b0585c4e6238e032f1e605e51a58f5ffcba1408fb4d3e89d78dbbce32bc0202dd16a7e1f14982a217a65c4a613c93875131f06db53be306b28dcb1e065e1371a3fb3150876204fff0359217a47c6232afd6ce01783c26da95f9b43899021c0162e32d9ad776c0a034b0f7283d96f6d8141946419bfa07a12a802365c9353a65dd2928901c75bda6f385132d197a8518575c7124b18c23c13d0bd308c39e646e3db45bb418148e8a5c23dbbde876d1320989d5511d7fd16aa393218ac8451dd77b901045d758803b5c26afd3334bbe0367e7ae15a5c1709339ebc2a514f1dfcc82bc6a0c589f5856c9ccf816dee892b65a2294953d5f4b9d54dae29c62164e53e479aece3a0b0df1b9573f90086a9866bd5175d9e1741be7da55a03ea94f2abf91f1645fa6eba242c4b3e776131934e8d53e59553521b1b82276c2a1baf55dc1139cad7f8a3df6d3fd13b1171d61c9b8898f74b9cd19073d13ef86d87e555c08be86e435a214ace0954abca64ee940e81a659ea9d828a469586835f09d9a80e4ef44ecf57480090121b6f2c1189719b5599b702c14a6f4768932cc556fd0da184615ebedfbd9965aea6bcee6df6b3c292fcc1b8bd42a6d9cb4ba86f87fb9f76cbbdf0948f224679702332b9092a224f119e74cacef29dcf77c52616f7683756a135b7db32f45ac5103b6de91c90adcb8b876d17ac5fa6a642803204f5b3833977957c72a58a9ee3e325285c955c9feafcad5165d46f6dfdb4ebec5c706f14a2ede6f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h13f4a04acf6122d953c12074c4dee734d94483b23f3bd7c55c406a29607099c4e5de11242c9cd353db6cb5cb3ab20766f8ccd02d88cd3e9cd417787d9875e4c48307de73404d7be2d33b142ab53065956a995ec148c7f819df4ede17079c7fa111d20983c7054fb4680d3f394fd6161fd628dd4f0c3337970036eb31d3b63dcae42aad185181aa4cb2c1b523d39e6a9f3f1742bad781727acb686551e236f356950aee0cd92a0616a81be662236a3ca5e189148dc28a02a7f2b0be4b5449d24f3d5141932393954fb4302614244803c829f9e76612ccc9490c09c58a4781c01700d091324e7b6b9590a3b405c38dc0817a0d810fc5eb90842ea3a5710924b9548ed189bb2da7e99e64756020746494dbc184544b7275fb63ea437fcbc911f7e8b704e565e94a5c7d81de7918684132ffa883a64b444343e58bee6d6d434f5ff1a52e19648b28d023b50ec614e5a514a7656aeb18733b1b9240dd69f96d742b1dbbb285b709d4a07834dede878bbd5f713e08d9ddc90ec83b21c92d424a7b03e2f72308c2d9aec9dc39371580478ed86f619813062c38b3f464c8ffba4a77c2ff209faf17e3a2ca025378a4721d7faadd7c04db1cd793ea9efc1d527535634e819390ae188a4309e90901cbcb6200d3b9f586c51fb934ecad9b79de3a5059697d3f2f227ba9ae89f2d701ef27b64e88b38d19681c5ef694298a18a5171e27cb26b2ccd19bc4bd4a149e423257f28c1f5286cd88bad451965189b62e72d9802d36234a884a6f455ba5b9b2d0f9a34e012df903955a600123eed5ce28ba8ec694ea51e9a7e0cd9819346d58b91127d12f04569ef9366bbce8eb1a9cddf6d3f61bdbec924f78ef1887561a089efac5381377fd170247728aa7c536cd5f77702e5d6ff8417e4f4842231c811bb5f9a0f46c0cf6be9fdce4eb4a1223fe5b652c6f56b22069fddfcd1d1f226b02635b32e2375781ddcb123a48392364373d3a32213b6d2d41eeac7c259c95b50c8c2829019306436480e257fd1592172d28e9ce57737f19f4369b608b97dac1154e86cf2532956b3419ba00b12a89e6fbf7b43ca2f5fd04365eb5a4dd5506770ddbb6fe4062503436baaab0449756558bbc6f5c170f267cb9f41b6523a75b0402ae86795c9aaf7f7b473b8a340c8c866ff1789056a9754bc49236a26d1d6d4eb2318a0574c52b9ed56e90168a7d6431e0e85de6deadad20abd912172bd0c2f82ddb1183a398eb176224616c69d45c7994d4c0af9aa77f7bdeebda8c2c51821650516e128d0afd56f24cdfb2573f6c82cc628dd0c1c9f0eac32cd94b2d310cae0ec91ea7d16ac6928d108e23b61bee4906175013211b1eb2b7543573058beaaed347df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc475186ed9294ca21641a18596a77059daed7766e15c4abe7a61d1b00d96be107038c7bf8140b6af75323e5e44d57e80eca4926b9b9f9dddea77a6590dfd8f6180e963b6a4bfb8d7581af8d925c1fc69946123bef36fcc1ddea937dd9f0749dddc534ed805484051f8c819c5b0deab604ebd885459a9c3605af8e8dcd7338d9b5bdc0acaefbf248ba08a19ab6ebbfa565b47b44c3848eb6c1650d225c3838f0be6384db731f80038c84999be367a1f1bec41c7107c0fd3f6591dafac73e90dad86efc90707d7690f59dd635dc8c986a8901b2e2f391c9721be75febb2b5d9607da2c4c630d273740641887c2b3f3c6f7a4546572c5c5bd23fd6af7a6d930c4bdd2f0caf2bba5757395aaee3e4f9a1da036005c884e5c9b8da0a07f64c9ee7c703f123cb5943ea30cfb3f57b566511608df2279317a8c4f89cbb41d7cc8ddc16f9fe0b067cfd5a562455777052a980bfc313e00712bd66150586d2a553620501a081dd4fb4bd86078631fcc3e772201120bb09c780cb867aac992727f2e4bfd2e31bca66dc826592d78b26b2451036f06fa446a1410e5c45f45eb8e6f5f79d991483a07e6c6e5d0875f999baace700d03ec5bfb8f01629a918774d4066d1c36be42eb84386f7da6a0f904512ea7d0425a37bd710a8c3c588e9ccb7de55f17fc2cb5b686e0a6c5b3453eadd10a76c3462a9dd0d6456b60312d60c86c324fb86b080daa9f223eeb168a35b621738db7973f08ba35fae2f05328c64323bc2c0a936a32f026c3aecc2f6ae799a9a8d748f63f69f7bb73a59a70c688e4adf7ea1a64fe87f6e1dae514137ffcb0afb4a04a559cf60dc2c5edfd2b8b79c7977fcc6ed5629253fbe2173d2edec000a548bfaf1474be839a40021ef77e1ff40b70169608cebae4186e7cefea2a1c5d260dbae847bd5942d94459a47877942a1126f2e062a071cb44f107705388a8cea7040cf4ca3f2b1eaa7b37e058d135f07f2937dead4f1f0b587cd544ea05022ab994ce29bdac398fb36e1ce24bfe42131a9ff949bd2d8f6eab173bbea200ad16c29749c058ce98791febf1e949d22f7ec46ecfe78c405ace449f8a43051975d11e4231fa9844fdd782e4a1ba6914b31c2d847791c2e0a78fb8dc05a0216dfcc89e7cc52e4b07499f905c87a900d3e073a33acba80dd80008da9726bf658847f2f8fee99768c1905fc65c0052f5904634a534435c5e350e2b2b15b4c9b5146972710d34fd58d34a124ae5e7428a2f18eab6a31dbc0e4509a3f659a7059fc8f453d0ffbf658bc88d103de0d261f8fef97ec4ecd62ac86189a414c4fe1a14d94ed3f06587a7d53582e80b08ec27ccfba0002756fb7038e686d93dcd8690c562fa95ab53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h166eec0e6c00cc07f2435a7f3202e59b7700ca2fc7a55670f8abd8b11a3cac30d90f5fde7de21547145b00befb781caf2adf82aa954c94912ddd572e22775542e2129f580b4de2890f50e2742fdf58d2287061427381ad0f6e56b6b30add35ccec1505289b06a0751df599bae031d3ef5a03ecd488e5f2a76d40b358606519ff1d1bbfa2e24c6269b68f3a422fe35dec243d0579cd0b76ba9079f046a0d4dbad4dc4d5e0f401b00664acb9fa199db14fea674079e31d354a3bd655962133c74a1a2e87585f47e55990b0eaaa613e2a09b2ab5b43ab637ac43a9770bc42138262e95fa7f549da8951144e40e61a9a86b9d6fc895e62d306ef379df5c52bf69692153a4df0c9b1e96b6f9a958d68ed0aa99cf6b7e1ac90967703ff864468ca7e1c404e927f6d9acbc8a3571be9259b8e3318945d07b8df7cf42cab0ad95bbd06dfeca0bf17381f833a4e8e9d2c31db2dc95988c8b64ee603b2eeb9ad95e7d162ac68e8682d0758dce17859f9e5ff288cd6ca993e6bf7d20dd0d2e9a4a50c079e15c8dabbdae852943d3737f7aa65e208e06a2ce31bb86fd468945e2703f68ed5a9893da5e73a2a4a04ba764102ee9c58be83b34862da599f0e24c825c7a0a34457f71ca31a1462c38ba86ca5d2223eae962214b911ddf0267b940f071735107ef9ac6966cb1889e9b20c2d265f533e55c34805f6842744f3cc73ce0e41d585e732216528d5d7dd12e19f297d496994ab787ccb362aa711cbb2e777886469071081f51cb026e7145ffb576ca2fb52665ef7a19256f05a7a99e9605259bfdd4cead214c1779a6715093a50823f6696d1f87c0dcecafb7c22e1e68e5bbde25b7586f3f4a82b874db57d917812bdc0565a5fb4fd6e71eb578bc7c208f5f5c28eb0e30dc3af5311eaddf2b0802b563b6172af18121d853c374c44d14f447762595d9aaa49b378feef61ecd74e896e9aa5704142873f0e96d5988ce99089b5acf9821af731b2f2d86ede191a111a0a9b5c9345475460aa587108b05b1683585b076aa138f44a65739204e8dea97997508424785236afebda8adfd9ce72513aafa6c1301f355aa666f254eae37a5ce61bac184a464080505625378ba51883ed4e3f2621518f1dd3611eddf1ee1c9ec94703a5390706bba0da9dd179c5871ab1f695229fce54075b58b16924e2274109fee9f1f4c670fbd492d7adaae6acf0a3311fe38175997451594f5a9a1c1ef9134481277c1f0bc701ca1b7a3cabc7bd600679ae7454551e857a8ba524de3f19d79f745675fddbb81c5f179ea06d48af22979f221dd831282f9d0dc4a13a898a6bf38a0bad6abdf06c909508ec3e6aa381dc788e1c30a0a6e281d616dca62b7fd207;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h53ee191432fa32e219040fa51d74397575182512fc5851c199a19bf9d17a11416167d85c908de94b53e8e6105c892ce188f38caa9ee98692d9bbcf6ac9ccef4d2287c97adf2daaf4db06f27fd05fbcac71a760f3c2ab10d4105421e1d9869517bf71ba691efc6f352a77083b0f1787d99a694b067f750c0fa8599a536bc51d62e5547e026de0fb157f4566087f0e0258d4ade222e2c39e30b170f9bc451c4846dc37fe63c195f08caa3da36ae6b5c560b76ddfcc377ae6059e1534ce3aa8489ad77f24820525a767042fc65c531d3f42b7674ea3312e6d896b208582309bd1a3e004d858663b37e0221886f13d45174b4de95c63738e1989e7d49050a8df863db6a249813c91d4d153d1c36b336467a8dc4235d5543bbbb3a9e0e796738a62daa198bfb387cc7598b38cb401df7d9765a9ce39029300976f6cd6423d0d2c3db01017f66925993e8a6324582e4ecb0ef29815aeac64d117ee56f8d749b802561974e80e01983c271836650b5662b376845f4975a065f1e18b27e4af3c9737bf8ceb51c09dcd4da3148fbad5b32e4ea8c9219ef3c917435a628621adfedb6d57507280855d4b69835c9e8a4e21032b52b09531bfafd49933df1774df4ea04f96d90ef3900e8af02b0f495d8eb18c4a44a5db506b0117dfa80681c1a47a684b5cb02d6df95739252aa280b6d7dddb35795cc29175162275926e2df2e540bcf1cfef66b5d703356469823bcc98f74e01caadcd767fc19a3a124972d3e008cb3e2f7d079caae73093f7510675cbf9f2981bd90296678ee41d6c4bf863206c9b695e206a2769653e06dc612773faf4f7f9e6f83d3b37e36ee5a492dca226c6867f4d3f61200ebdb1193f39784aa5315221bc7ee0191e19b760b4f785931ec6f1b51af58cef9114789886e384f8cbab072154bfacb5d928712f45d51ce222829547dc2e36e2ab8b1769d242029dd29ecfd7d1aed6357552c1a8bf5228b14d689fa3bf6d545ebdf1731e817617f688e52c0ac280b0da23068d4762622b9c0a2dbf568dabd647fccc0413d254a4a4abe83a99c5f5b2d81a0d08f5def87531f05fe3ecba23293471032490199e83a10a84c4a8d614ef5a44ffddd78fa007d3f46df5f57feb408a586526e9f55d6bada77a92cb8ae1567e988d26715444ee0cd13924ee2d08e0d42aa22727eba661d7d09a1d0859b814260977abdef97b186b07e575b5233afea158e740879e6a7600340899deae4849ff225045ca68c0bbbeaa6bb3ff20a4b9008ef1a7f5c66da81646acbfdf9778a44629bdb6d31acfb375d42c93f8201d253e7dd235fc5fdcac3cb34cffd3d171838d7c5e7e0778d4af9c814e070ee4f8911354e12361b72bd3463bd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5e50de6b0828466ddfc843b2d33ac8280d45e5233501eb6967b1c1ac619b7b9084a7391584effb631e5187c03d219fdb8f74791da240eec187df72d15c229f105aec984f1b41a8719eaac9f350a91c014d2dd32824ea205fa4d3c8cc61620fcd5296ba7b6c3785afff235a2495ddcf6913d75027f0b05294f043cde8528c87f8a885f5e5cab36200a72012180a50ffde979ac9556063a16b0c4b984ca5ce3957a07b1f940aaa1b37a737b607163fa3b5f49904513252bb19d72ec8b230da7c3236ca7226d5cdd3df9200596ef09085f7c65233e841762b1cdb39f6ae80a5acd27d1f8c2e985329b02709d8d113d9f7596fd900675516bd608e45f50301125e9c2bca7f5240ef499e3a0fa5a4edbc4cb8515494c361a483e565c4b49ec2ca590d2b31ffff2afddd078106617c36037a08a634d8c612c5fa526832fefc24c41e95c1ffa8486c7fa537d507c90d4821f0838816b9a536cb49a5f90048a5f5b9af2449f64b564ac267be038faf471d1e8ee6d9b66def180c5f2a9c8e5ac4f169a521389277a47e82e9244ffb7745f613ece7783e4f093791cac693a107676b4ee25f47fb2186d6a2ae3a0600c0908caa82781589c34ece168c0db0f113ef7abe4d1f4d8b73a7988d61c84a346e3fa333f5c86800f2c9e39f8e7c3f292d8adb44dcf30cd40c04cc7becb6097a1c2f9fd18d96fefb2ae69327308abdc1deaeed4f9f654296b12fc9cccbac271b818409d93d2fd78bf94e449d291f5562bb781707af5c5960fbf6b4cd5bcad12c260aa3489790476b7ff9b87862170a2426f8d1d1ecb110a9fd2c47bb14282d24fda0653bcf56667dd78c21fce5a3bc6687c1581bdf42dd085529892dd1d48a1fb9289cb682ead657f6c324d7f91d53eb947f57065ebaa3f5ad6d0c2a46854b5be8ae7be518bf4b6c39191d16fc1836c6eea97a79ef4b058f0300c5453d0a239555507619b23e4be3367ac6304d820db1d5a7eac5ffcc6b7bbfcca01fdc1cba68045bd54df140402baa92ea474d3babce3af495b363bd1a8aeb6f4652b722c61b068ea2c348b270d6f805f8fedaa7a103a62e6aaed20523c845c339dfe6b06bdb4db9f41985cf7f40dd30ee31043d51ba2671f7b7d64efe78509d3b7bfdf19ec11709ea548a762aa8d3a04b1df289cf151e4be49067270a9f23eb62c4e0d02de04bd669ce2881a824052e14339e43db4613621178fd3c028f2198db0feec59448f337aeea810565530390860006dc003df185138e95007d287c27654e781fb8eb5cf625d4472acb50149fb24c01f4e9453e13b78c88beab3657dd7b2a1a1e49d3a6b4e1b1fd750e794a6d174b5346df6618d8bcfdebfd19fd0bb3be37ec5e4083a29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha31ade9369e6b05807706ec9e4de085fb3481dcc47b45685fe502e94c35c567e8822eb21e77f8a65d7e1cb2bf19422cdfdd7d521bdb564e3b97f880e0387bf0c0a9732465eb3097ed98433d01ad3d80769054eaec9e579f831a2644903c22e470cf5289b3d3bdbb77bc406927547c520473c78b531f4eef9414b52db24b5a79920c95f66162f600b7fd413c3611c6fce8d07c8629029cb5096cbf83f898933c26123ada9c4f52f412cdd4edab155d9a8f32e1a4cedc31df19b2677da257b16e0db747d243713f28d0b884ba568fba6e1ffab42adceedf8079b2822149fe3a08f941c456e3865df56b27aff0c1e63727069da75a10f56e761ab5f93b3a2cb90cb418c5cb72e8599b1d63de6c2bab31a867eee2944afd49953cdebbe3a26f9bda2187d998d6800704db619caf014a0d278762e3d1c4a92fd1d9fab30aad7f4cdf48d0fe37cc73d3e777885d30bc9fda4e0de495f7b03fd427061f81c3ae4339a2f83250405f5e15724e9443586bb3817fcec3a2f00abc5767766b5988c2a4460f768438e764c90bdbb048e4e23bad866faf1bb5345885b9904b97c6eee989c040cdd238e47ae7d5c908b506e91ca84e65556fccffcc1e1f0197b0dfe9f221b7e77e1bbf79e14d395a260e9f271f5309a9e308d51e1da6bdef2f81dd53b4c3d02deeee7db052f386d3be0c320866f8ff138a61a0c9d1425535b1a264daa02e469f01cde27c7024269d40c073095e0acaf28d943d060ed3470fcedc3a8b916e64e1f94eae8a2e93f17896ef767b6113da702b5361dfb2d0947dadd4b558c476603a42cbe63e95ea935d407b887ca0289e4415fa433fbd5a9e5ffce818756985c401373e51e8263d0c6d69779300c6c3e688868c8224f92eccf62550a1d88c49309a679d0f06075ceceb17e0ef0806e43eb03a3326e783436b82b8d4a8b1b636a0a341c0da801c0b8ea05f43774fa5bdd65e170faa290343e8ca0d5ab27ce448001f5a4e990e839342b0c713d7fc75bef48db0ee1a558365dc188b6eb858a029119a061eed5a1bbfabffd7eb8e544e24fe7fcfaf639019080d70a6952b8f4b4d016c584cd1ef5ad7e6de9bae076d10f9834517195e2921de5a93ed8511167464bad3b0a0443fa1a5f3eb75d2a9501c568d35ff3005ef6e8d204be2dab75fede52baac17af96fd2824d6ec96b04ca3ea7cc74fbda6aa1a78347e3a197a2407da66407bdb59f0e2ff5299f1d50438a401f8861c8054d6b6ee366dcc66f011eb70f0224ada3ae3064bc387ffded4d937fd45df1e20deb571ef0c1a072fb00195700cd42bc60c808b33eb8bde342223f1e18eac612159cda2d3bb8dd6ac0fa533bb20529f4b4e3f004eab23085d9b83cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcd79ed1494c62f92d21e09a8fba6f261c95337ca15f930042e9e4ff0264cab0c12382bfc55d203bfd30abbbd15de11ed78e75adf262d132dd6368c48c5923c9911265ff0544ab6b3d2708ebeb5ea7c327e84b440bfaf73f4fc349c0af80a168d86d64766116f779534189b2cad64fce262aae4fc9038b807a29fb5beb11107de86efb14efa83fce68d791b070e4f914e09e1abd0bbc781d9fa73397ebb3b34390e78994ddbe31b795a560b077bba817ac9ccea8f683583cb0d852a0c3e90fb626c73d54d7d2776b7d08aee9b86d9764eaa6cf66e844674f6c2e1b42b19e323d4ecb5ac0bce61df0837c77b24a8f49089ee93922cbceab24db2e09499747492e747b1e1371cd14f8340e6fc1adbcb03bd7e0153a8cb1a22fcacafd0d6df8c0727de456ff4db1e00b99cba70a829910315e9d02ab8101064c7a3e6df16473a8b66c2361f7ea5ae7f5b6d55548653953451fc82707698dde151165f1ad629f80071adf239cfff29badbf6e76eda5e7cd1fd5d801b1983c87e6edf517c91c458773a5550e0b5cbeebff2c62c4a76b6df949ec55d8ebba36ebf913443ffaf77ca3dcfae7769a40c13cc2705be363d770a9c0a8c799f3697a789e0a74bbf204a5650689487026448a87de24853741f71955be29a9ab042f114b785b4b47174702b950e7015030e48c5024476c6ea03543458835675282f3668333a9dc2584b35baf4a1a90a11c0ac7c312c9f22ca6652d0602b169078741cf6d05cd087343f38cea154b15762d9fdb55f9266a1cc252e7a233a1e77310e0df72fa669cb8d68b1c8dc4fa532743c32ee8ab0491bc0c2bdd8d6bf4010c4c7538472cd8de871b8b49aac65e4d562152b58e7480292d182dddb269250d226464edebff7aa4e6b6e83ebd78fcaac3099103f822e58c04ea0715af3c7ba703d54c2c901d813c62dfc957c814469e85777e629bfdd91c807128c54ae88ecafad7e5a3fcd200e952e5f4a2422e4aeb3d7f45cab42888b8896a66022a578921c1ee30d7b0ca2e42ac7f5ad79fe3f8e8374607cf80650b2d781e6d257e21105321848ddbb6e80abbf8741646d985f455a17a439621694bf39faea0c3c8b03d2d8c7bca60665a37dbf7aa03853c67c19a3f6a3403d14de365bbc0d8ddde52f8d084a3197af016a7858903d0e69e8252ba02f1d6d71f0826cfe62a5c4bfe04cb48c1d8dd336ffeb08b5665ca5eb2c793aaae381e6dc5f6dcc229791d64bf281d9ddd128c7eaed4e8833339ba6021c1beb319fc36e442158014d68cb8a7665cd14aad80c1072de50f980b964dd634769ee08ee6af83cf81459043031af1e30cb056e1273fb133d04d2236a007dfbb12906bb0d817aff4a708a181dc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd5eea55a9276afaa78d2b930592d03db55995ed29ce1482d563284b20d4db4f12cd1d724ec19064823cb4d0d7311c92a680e5ebbc02a4c33ff7f8b13d4350955f92928181a85eaba20548feab5d1ef794768a63196d2cc65c5623794c10ebbc080647e8f5118a9ba9b4d42ac011c35308262decc3791dcbb3bf1c21ced8aa4794808e090cfd74efb83307642f69a1fa3bc459a8f8df400cfee3c9a8d5b059f050662877d27c9219ca15a3f32133ad54cc3853f61390bc47858e9ad5e80bbc55d4c348a07c35c2545e816865d61c0e3f4009dd88296109eb17f8fefdfc82c909f0a7f0552225d46691a989cba8a29b21b805125eb1ec5995312a8b1e37e41efa081d0fb7318e30b0517cd2c00defe73d31dc4d7b8e77fa8d639c277e0bd921d9b2b79c5cbeee17047a5708f64e496b441731af651e66033e5f5533365bb6770dcdc2bb17f4e06a0f74a0c36e586d73eb2eb800d93283f44e3a5ad720fe875b9ca71e38245c1a9c6054898e9d9c6f1e54fa740a9c704a06a46baf96ffba6088094ca318465629db2f39698f9e6a65bedfc74f394c10e5ef8f4540d3921fe0cc2da6db15bc7740435c0008ffa0ab4fc014b9ffbf266e037af579716d3408d79ef98fa20ed598d265eee922cd236f593db5071d64b0133e6bfc1f8051c160ae51bafde3a30e7962b8799b3aa278e08bdd215f9ddec4098d21aad65000ea07aa5c6c3d0e9955ee87caeed1c688d52cf08499939935378cc0c8cfde21d457bab9397053ab9829b5a42b4efcd3e73783f4c8c2c5a71a148d69b23f728403339366f793be904b80a1163a28bae8947f5a0dc6a1f9eb366aa5681eac0618b5d3d444f3ff2ece6e6a9d32968c53d6b29ece461759566a7061b8af36d93e4d49a0a1344c6a8077a3a4cef24a9dad800ed9c276539fb8ad46507a48920dce1dfc73ca219770d4e03503725cf3078717eae9ba1967cf1629f3c7678333f1498b8476643ee1ca9137a613e0ba9d32e0a8cf4510597cf55479cf431aa8f476b66c22cbcbabfa99923109377cb126a42d5615dda7295e465961b211646529f574a9f22d47b32486ad6001e2b55ad4507f1b31c005fe265d74254c1fdf9287201f19c93b5faef926fa73479fc3d57531201e6439d9c22f7c28526db7e176d1a251f2bd9e265fd0618371ab9a40545d8f6c6a1b06d4a243efcb6b5493d92ba6ae31d79913b0b8ba506288b4079042879696eedc71a1be0524d186c677b9253d61fd91bff0cb0d9b2b1383a17919b84dd7500f607d7155011199d8d2aa81b7aeb2e469ff4bb81b4308e2d653abe7eec5194359ad415f7f3d434ccac65955406de266750a0c2091a3a528dbbe8fd35bb8230c27fb687;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3fd61bdb755032562c73ac3ff2d72da848d85c25e2461b9a00047bc709ca791db7c92acc1e986cca91d2b8ee6417addab5f1c73df3c63de679ce8bcc6100373189eba7e026eab20194fb6455ce4ccdb3758d8681d2a76b7f5b5b7f02fd4403973d54a9cf15159cf84d029c9d67d03e9877f7a440cd4cb3fdc156fe986bef0a33afee064a9ce8b58b963c7932f8241b5ae69b65b2fd9a5d2cc23e7f4752685d0bbe0e04e391085fea19899b40a1bcb9880cf8a5914e3627c92ce3f0801eeee031cb2aa8921eae996ef32bb5d49636abbc5d67c03ff5d28ff6eafef1d67885f71e30b937057167ebb909dbd2b3d86a15c8fc9800acdbb93195d12e0d81a99cf7e6b4db60036b17c63f3589bbf330ba7ce5e97c965dd4448d8d3b9e0484aa7aee06300a316df1e0b3e6dcca2b3dd00565e2a9fab5f2c2793252aed8de1c56c8d6224b043539dea3bf02926b51c45b02736a03320783863445959d319b5c2a8f42fa3069883965229f858e4f732e72be7c027c2f3375a232fe49be5d114760c0c80660d3e6fd532812c160c506fd9cca3d9bdbbc18bdcd9323d74da7499c61550644fcab47f24ee30b0a45a2ff1515e551e7cb38abc01a60d6b8b8a23b74a636288115e34f8fdc061a133f975d59ecf6d86d067eab071e891f1a7ebe72ed94e375024605eb6c1a72291a730889fb79bf5e05cd36282291d626aadc8f61c316551973d2a0e7d039ae6ef56c26fa3bd390e7669599af5d179fdae4fb57dbe4635b1745ebe3ed3acb907e142f8ec2013b254b41e06926ac162cf90d2389b9179695c55594e559052fb25642dffe85289001eda55e953f55d9ef165a9681510d0e642335bb388fdfbaec756c9db809bf21b980be177de6b74fb1df73d1b3ccc9ec4ea3eab0364457f5c2dc4cb3765a1f866e1dea0efdb41621073ec64387cda1a04f844095c2d5525d9cf002b2d312b12e2e0de8bab9b02c9e264a7c08b63c63da61eec10e2c41f47b71d2dd54880de49c62d58d18d237c65ca8f54cce5014579bad613f98586d6382997c9e69972b24b510e4cb74f2f03c8c376771eaf64c6611bab7a1729a336dbcd716301490d9dab300f187058f55672012b5bb69dda60aeaf21721ef0bf0849f3a143f9c1f0be1039f6b798d1ed03d4cf4ee4793b32d7fc920e87d9987155345586d4d1c74d18013f977d9b10de1d9ee1e288244307d8efa21d0c50586c52f95efbc539fc97417f59c622a187dd3d10e61270e6808fbd8be8a5554cfc31217c7671917ad92a7d721024f97eb33fe9490a7eff57912d7cbc7acb68e2b6b873b1f4a1635df67ed2b375e98b9d8f5f9fd61309636a6141eb15f1801da0c4ee307d923d10e129f29f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h85c787437787b03d22bfced1c796ac3adbf9c8af4e1cd188ff9ad31eb69e91d55c9101625d207433bab9b68e90cbadc5138b2be357d4cced0133420c89c90f5b69b8c6b29bde06005ecbac22a979d709019704a39d2d7df45193a9c5a61c7ea81073bab62f09d71b62391c46502413a2fa436daa4f5c48b165c655d891c2e8204f4624260e8d345fdfa57ca26d1c0c5d56953aaf451066a0ab018d370e0173a7b899450cf8d33b14f61349b2ef4163339f4067b0c0fcc6f5ed25745015eed9896be3556f56377dba884ec45b326ac87db46d271a5110cdd1e855a0d0dc133fadd96c0a141e1b977d94639bc1e37090c67c034785fa1a63457a905a80a7d7dbff94048abacfc94334aa7aaecb32dda9bad6a2a985ae7b4d6f00933970163e83f64bb0e3210133f494e014e78cc90a809a2fa366b3af5c571808bca66e5306e8159a5eb7c5d2faff30f606e5ce612d2eae12f5062123b731b249b82220a2fe83f0f9f11e445c6c406ae121a145379eea7349751977aff2e7289b0c56e4a84099c2d177adcec54adf66eeb22a55b9996369f47e70048bdac4ef63c0b65200c415162eaa93d347bd5785a58a7e1f691e1dbd88f76fd1c5607d76a561028fc002c91b41f5fbcaad381d5dc8c033b8a83131df3534a4b54ce2d762614b128f992856c90b0b5aed3497aee8367007723e8c0ab800660be279e018df484410fc3e52d1be79f7df37ef88a769a0f92584909f44fdc42c0213ecb44e37021a3bc0b555cfe84fa7f1e10283906782404730cf65add9298461465de98495d9eecba3a0e1a1561d1efeaae4df55005228094db050dd27c60157e026be0cef103056b8afe44933b491ffbfba131e86bb7c5efbb4d16064b70b337a1b86c11b14f697f2acb305bce7e11083e827766e0f8d6e97788c59ead7955d438b940dfaed3954d9677df0359d7ccbfb2ceaa05d074b78bd0f4bd2ae2a3aa30f0e6939f84dc8e17a78332e9071376acb5e5bd2a1b6cd644baca6d06a8b421a1e04f1e1162e08c53a72844bb4c63857269f0f7223cc2c3959277349c8cb816f88e48e8c925ec87e7ce8f90fc3154ee600e72fc984e6c56bc642d22989f9828d97480314e5d18ac1bab0d4fe805c1e73239d8509df8c0dc6451ae2e61b35e400b444e23f0c43c141ef461fcc3571f0804f206cbe6e278de0de4c4b8434bb20f9637427e198b0a540ffb23845a7e6831f071372415683cd8c2f980570e5a0f74109181ac8d45c03482012b07b212f542ffab466bdd898989ae815bcb27022c4b29dc91f51601768365f4ef1f6c5ea0b3052f8053e949128a76eabe6dfa5ab2b547b7ab79798f70b6fad3c1ebbf90f4870c999023960943e2fbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdc4715cdd9eba49bb76764b4115f2a0f7ffb976161759d900619a7d928abf4155ec6f745b89fb023a8e5c4a49ff5b3f93efb6d56df8b3aac850348f9dfb6fc66eb46f54ad7291304fc82baa43789a2f6f8c7370c8096e648ca12fe1ed21b1a42e14855df3949540663dd6908447d78d2ef85b42c7d68a0fc7f3d1bf773187279b0b614176a3a0b7c974eac7effca32a027e375daa48f6a0d3e2b414babfcd77bf31c903ec6ffb54e39da4c8daab37345311ed33daf5fd2cae7f3b5ef13dc2077b346699c15d64d7b41df123a21dde2f57fcd5f478abddf67b1c5077ab1cb1227cb285c53d92d66372400da0a423373cea27db4bc987c1bd8842fc95c72e99c00e5c127d01cc55577ace375dd256feda8c1ccc4c0a270e3efee0b567737f0b8248e700dac613fed33ca97081d42eb54a94418d12e25c7855241ba84f239d8744f46ba4bd68926cba7794af28e62ea5219375d884a1c3bb9201142d7d917249f38bf0b7ef3c23cfd01ac59d7e37350236aaefb8ff0f0abca62e2fc94f236f80098ddbdbc2252609ac563d72a946fc6a759dbba64d090e373f59cd5fcb1b0a31d2d95b65070fbc4aa34cfcef12bf150fca9a40c85de0b77e69584d8ae872db82203eb82990507fbc3c6a9af3ae15c5a047cff1f54f7cee0f252b2e729375bd0a93d1e470a2e395ea351eaa0c9eb3bb2c0a27da36cd2a301e511b256e64afc089ff569051313002adf6109b5b254c44e0c6d749889af1f2968970bc7c659696184bf0904417bb31bb5e9a2cfe9e8a79be2c2a1ee7d57a3f6aa11d181be92944ed4dccf14263fe9f903b8699eac0dfed378b913d2b31c76e38ff22e20ffa986e28d38d0bd4f8e071bf7fa54e89d14eabb32f7cfed735ebe416bb98d393149c4f84d3ba0de4a2c270cabe5bb0b33926292316cdc5c46560f3de1bbb34062aa492be9e65c6fad59b2af6e2c0e342647ef2429653560582b2b5b18cbf4aed21e156152a80264e3d93320a9b713d6de9eb32a7deacdee331cfc899aafba26da3be17620a67a2b93e7adcedb4378f9ce8fa98dd0fcefde2721d3d726887023e0d7fcdb5077c45c78562c799738904ebe8d165a1c38f3b52aa62119a5f305b3faba91b7979acf674353ae38147ed456cd88afb9fc2f66d6c3242e3f161bc2d0f4e3e432e2beae91e068f08d9ba9d2b700988281f4b6b40bf0191f9ca61093d8ea42b21f1835de73db1b4eb4b67f7692caa3c2b7c494eada7f4d99c2dd43d3690b3e4b1b1877db1e088ac6d28a75db71117b58b529873102165689a1d74b46ccbcb79d48dc02fe77968057d16f5a8274ecc2bb54b3906b2d3f7f609f397276cca10042df70acf9a40ec6d1031c9adf544d46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb12167e242d7d9f4eb98a808cc84115316b846ec6769a878a7b4ab9073c7a2ad4c82e8395cc29de34f3783ae4f107951496398ff0a8f6791ba4a79507967ed638b8519c995598b898a4112a7e07785dea5dbd9c63d4d8f2fe43f42db1630c8847c9b8c979b107fac2807e27213b5145f11964220ccab4395408233a6ea7cba1a4ea5b61d322c1b214e9bbd9f7cf9806b3f8d9787d3a23dd696a95f1f7862d2adb781e88adadd60ebd17167cad19eab1baa2b52a6a85cc649c87b78ec25dd60eb4cc843e4d1c68aa85bffd45b7e24e754194e3003a4c62e59b0db19bb677f76b5e715826c8624c2d468956146b6207aab3deb66df7789c538d12cbf252dc6366263bfbbb4feb9255982f6ce04673ae3ed342ac26aae799d718e7c6eb0d64f9a796e70d2035dc5addf8a9551971151af4a64deaa809c716ed525e5a674b688116c344ad853f781417ad20af950cc48a917bdd4e5ed8aaea0067ceda7423983f3a1474c3bbac1359028addd6c909ca28aef1de495e4486f6d595e8c49e26fc44fe530192847bd0a377a8eb7299a57045ceabfc66a6bcaa4f599209f972234eb7aaf1ed96580f3501d970ada634019bfed5579ddb0faf9a81b124d87bf8253c6698af518f0326cb193dc4cb4d3bccb66a408db26fc87561cfc7f9b4546f3bfc212179c58a92a3412a999743e80ef4dff5fa1fc731ae9ec3c5d03f6f97b3f7c412558bd1310adb0cb70407d811083f6080e8ca59ea4712106e80450b240c1eec17f443b94d6d80635605aa0b71250245cc07cd0af609bebf21b9f70ebd12ae716b8d962f6c7da02028456ee9ea8e6b2df355ecd2211ede808bcabd2104db8e8e91df4ff27f1dde092791d637915ff77225320622d4e2fe398fba9c7558021d97db41285b531c2258ef43ce41129a1a077583a5f18e66886d7dd39f8a55054ad35368e2f1819d3c907ae64f4c5859f93b62912ceb3d665a91fcd0a4e78caf207f09ef672ce2f109743f6f30299d70fc5c0013b30ab2d27600faa623bd9d39f03be3d1848988a21a284ae4532cc03d80680907ca5b638765097071614ecd95e2c64df52cdd713a115f9e36f5975b94240c296ebf9a12e14e92b17a5fd42863a1395d865c12b454aa4d133d2a281e820b305ac4bc0ecd69dbd8a92f9c695e462fc2caf13f48a72de07d2b2b7daa907cb8413715f2b5a1fe2425db56c490698892f43f371359fa3bd3890442cf02bbac12ebbb05ec3349cdda42201b9599f14b8b7a7f67696ca92d557e6ffa7db13f2e7c8d2af2d3609a9de54e62280b10f9a5c0e51390d6b901d993cd6f53e425957338ce3244fbbab070d202fa0423d37266d578b5d83e6fe7f792044533f8cc85711;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h589d2caa8b1e914f4d65e19565e302b13c4bfdb51dae3a7c20511b800a3cf7f7356610a28de9880fb05d8b4d58f9eab7b28a868a9e1ea3ebf580465f7ffe5b665b18d54251577da80c6b8172e8e767307ab2af618c77528c2ffc89c877daa0fa2893bfe466b2ffed09a255c0cb8a89fbeae9a8ac2d0ea30658cd1bcfd5b4c9db277fe1f3d62078ef63c5635a17e96418933897d40c529c46e9f11534db9418c8e29ddfbc3c73d8e0066f44696a81aa9923c792cda669ebfb2cd035593e35ecfbdc0d2e641a8a550cdfabac622c2ee419e7f1c60773d12fb2b8fc51c8ef38e9bc930cb58c3a373e8a79e8c11dd7cdf2dc9675b0a3e164b4fa36a095576e064cd18d4709b74ff88509f151d924f2919b76f35f0c39cb24f17f22f4e138268e7201d52d3b7a2a65b1d10d854e6690abd18cc4b80e24ea982eb34f5bd7f95540a57f04e9ac60582a516dab93cd5040ab0cccbf20f43163967ed856b29f4cc6aafec8f984cd6a2a6fbaa2bd0d29695fbe0f47e16179b8b6df9bbaaf35a32fb1f7d6ff130adc250d6d9a0ad785517e0321c7552d3bd83ea6b816bc039e58022b23fbe2cb2caff608faba476adc0819a3fdd4e95cde0a4572f526e20382a61a2bf2324dc80d879f708df674770481f35b417b5ccdcc4588a1569d6bb0c775725effdb8e421fdb4df332a951f7533a2d9f736ba6616459598f4d0120abf8d9eea2b496b60225f26c95d76b76b55f24866d5f4252d0046d23fa170c2ca1d8516aa2aa731f8afec30f8bf3e7c60aac49d1987b15e964f046ae38f65e3f96ae28b6cccf06eae98accb5a33ca9fe7059322092539f22e999acd5706a6be88feeafc739416c9ad90d402c26457359ea1b9bfa59fcc7b57ab338e0b0a8598decf1b7e3edb2d4c3448350090f1baf57262da57036daf067dbf3d9d0b330596f67ad3701815e2076af722fecdb54277e9af57d4ad75d5ca9c72ddae4824967841723e469b1a78e2b5eb3c7a43e45e1fd66b87b76f90c0172433ae66c02315dc879c7d67653cb5f974ad49e28981b8612fce1535f71e2fbc1d602229f41b9a8a732aaeae86f226ed323a04ba51aeaa3aaf40f290c0db51db989c7ce17ee1c9d34ce645e7046671df9afcf83d41e54e304f4d14da1950bdc63f225cad89b464a50232cf6c8ff2f0aa17965a83143764d89f6f480bfd5009daeb7217d2200b5ac9f860a94b18049d549dfc01e64dddcaa37f78c64891c115b9e88147bb3c6c8a63c0731e7fc4309ee9683124cf7b5c4d9fd0cff9055797c6496c3654572775fc0db478b14fa675a72c0566738c897712718066288fdd5b848b0809fa0670504a3982c78e0b3de96002d3a103486a0f287c38df2fed9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcd9c765911a7a506e0a7e396ea2089351ff120ca93fa7e09b4d6352876968ba2c7c2c0345d8534eac27d55d488f8bb52be0b8fdb329756b57a7902f7c7e25c4e716c8c9d85c530caf23b19833811fe564d98c96f368fb07f4a963c8846d0ffe6d6a3cc64120e1eaece63e6a8e13dc0a8673a64c4a31450de08aa8d06a57ba7b2ab493cc6521d6ba6a1b2c958c911b6e732187d9f546cb0a6d9770bf8b1e7cc920841f31f2a69d463e4b6eb2b1effd26c90ecfc6cb1a249d6210ab534f798fde85fe9823e57d60aae1e2d45cf45f5940ca231732d0ba3d913b2473299f6ecb5cb9bbde22154afe564975e93f5c529634b18f4015e169dd9ccc63f9b75d608197713a1b12b391c0bfd0e6aa430aff3f21ef21f5e95ea82967f5d5aacd6d0742eb1a9f8ae916f3ff53b3af7adb79bcf6f23c467d1ec8bc3d476997f590d49bce6399a939ad09eb9365a7f3842e25b957b06d513c065b1764178a8b966fbcfb96ed101509f04758d58cccc6614f87f2cf5eee513da09fec79e48d6ecf2c4d658c16fb2828a0fe2d95d03e7e642361589f47140a7cd3706b0625f4b23666a927c94df6068874209dcea7069a8ab6ffbdb5e5fc7a01259f7dfe7a493c3a01ce8adc179b93cc7caba8eece1d19dedf71d4a1138e0958eb10330e731b0ffff3360a3096e970a772df832e6734b7b99600af40511eddb978ea73a6413deed4e7bb429ac8dc5114009b794b4be6a48486b703f30fba90dc7882d16c8ff0a979eee8a7f26b448b86b7a7575ad726659b2abee051ebf1745791d33e481eca33703b0d2f3557cf6e2c732837310af4e4e47b1a43e10ff5c23719903aef1c64ef37495697e04a1fd4ab48fc6f2561992da3b803a1a8686be753965f2935566c4f26efde7f5b4a9dc92374f8a79df90155561409e3faaf36f4ce41b5a67d9254cfded4e4cbcc6125500b5470b16979965dd42585d119e37cac51cb2a3225a10fc63aa0308bfe5c255445070947eb8abbc3f7f0bd1ad4b78696c6f4ea4d6ac5a47ba662b831637115f3e6dda347fedff89899ba79b2afa7aedd024686c52a61d5868b849e22ded99894d6e85c88b37b65b87ce767e0e30605f67b127fcbf6650910da886790f71d524df0f95b662dc9237359c0263a1c11907fc66e2aad6d9493df12c15c858ff380a09e2cc75632631fed11532eb5d7a6b86f838bed6236bad46004761953f2be2cf20249695ee79d215191797774f266544df31e05f445f5fdccc8e033712e63c8376999e1f072bc4419f326b6e0ffb4e8d4aaf880109a61b99a42138f1376587c8982d750abee4c71597c8999effac8b1d4d56e37b535caa53047c8f416b96da4f2379686791e456d229c095;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf68e67ad7543b8922fbf5890928f6530b2f7a67046dfc650fe6f661e6ebd2ed4b81b4c198e9bcd2e84c0e38ae38ee5df1fbf2539f065473b80d45fa237215e8486dfd46dd0dad4cfe9e9e3aaec62cbab8f039012eeb2e05d2f353cfc527e6af415c31d54d3391bd87ae3e4e55c48baf1bff626a54841f8d507913b1c4df2dff8c5a5b844035bf55364ea14140402e95c71f9f2067d31d61cc9834f55aa12ad2d2c276a0dd9a901e3fcab25e0729f916fea2a9b7c7fb0f3e255db30ce041343a79e743fa2a7cd745fc779b239bdc8f37e0d2d9425720f4f60a56984892ab432932dfd33cb39b5673cc42512429994eebcf3f6a3905ec37270716836b74f92437f5a5d5b7a8c1d0f81837a988837663ed50247deee99181efe21b5c68cb7c578d5528565b2d358be9eaebb6fb3edab47d8c774100bf6641ea0686eabadf6d034a314a18db584fc212e332f9781e9d71b476f2814df6dcf5a30f0c6ad3fc8facf5dc4bc791aa2659bf4cea0565937c5161263d051f18916ba170fbc731593c8a0e144288485fe52e6657c0665750c9483c1cdb1bd205a1f81701e994d19eef94dc864d3beecf06b84856d311723633aa7fa2cd34732fdb912d5a0b20308616c893d876545a329adabec1da9f7f42d2d46174807812a627b6c2f55a84dd8f72d47a6f2f0b2fb4fa568066a2b162445b40ea22ed0f8827bd21fa1cc2e23e2381684efcefec2de591785a0d0b86592b28344e3cf83c66066dafcc9b05cecd903fa4d46f8f30f3e50cf2a28037125f7c82991f729c6a28652f6d74cb9b590d9de6394a24e7839b4b7f87ee83651a3cdf52b08aa5d00a6db181061a69294727ffd900aecbd4ba957330254b71f7f589288300e589f8d587dd0bd9d3732917282b4022d2d842599918cf7a67c0b12552db3a14b06d083fb25b5d76c048fcaf9e1ffc468d22973002e765f1bf96d268a9821204b0271ffcee72cb1b4ea050323c43f901d7ab751f6eedf005aa167f46a37ff9a4456d483f854d3a42feec4176db237df73bd1127b247138880ad96d68177f599b6a21b77a7f3e478d2ad40acfbb6645c3ec70a780858fe9717d968c4c4030c3f64df22f90605c09a28509e6da05d1d5b05a57b9d8d73dbef13485a3dbe0b252631a789bce0f82308b4ec6fe78677f31bb218a5344d30b49b5e039703f5e9c3253c8d3239336b05a86e3c4db4e5f20c47c65e65ed41152edb5fa83191d023ef4f84c103a0f7f186b670ce6e813d69c4b3158d3ab574ce7a79dd75f60cbaea6761e9035c970e04897c80f7610b344629b85fbc64c994faab3d85c9deb1ea29a1ca8a8d55bf736b97ad43a8b9e6049dfd167d6bd4c8f918813d9b47fbd8b66e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcc5eed1562b3b9a9b883a8f857a96acc068883c5862db7ebae7baa721f1dcffbf683de30dda13ce28061de19174c1712f147fb0cc104afac5626fda9a4e0c5f0ba4a753c0fba5bc226756c3cdd6addf9d3451e27421bb49b0c422af004fde96b1ec587e3854a52d5b7e3fa7ec1745897e7d9186cca5157fdabd8daba20294289155533b7f581b40707a4b2051901808a74b1e4e13c66995e4eed9c624d0b2c95164768e58ceca75098e69c5434c1cbb17a0c2678f8cbe8aff546cb62567e416f796f27e42af0fe7dca2bc63f864849e3e098d1dd5b60de09a92024856d714bb07b26c8f1be6956c8b652da8a632962de611400a0e6f928282a403187bf392a258875186fde5aa9714debca2f804bb934b1184350ebe3f6e048c110b5681ff88e0195e757bd9e8f40deb0353d2c5a3ef627badfd9bc965fa78398b036f3abe73e9db9877d1d1a2da9d8bb7e04e17f32a06bafe9567afc9bf64d8f65c76f43b0860c44112a4d5b2bef7065359e453b59fddb2f8c5dfa3e48d729a526f60db200eb8019c798c7a6b16c5fcbd0bbd1865dd6774741a746dc9b549ab6044bf97cdaea652ec2b7ede93792e9d11282a3282f08f3b270ff53423302a82464fad425abd3101dabc21ca00f4f75d08fa0316002ad732ec7e6fed24a34c2c5d578f95412d7e7b9616dd40deb2055ec7ac24b0d7e5244db14c827bfdef7149d0a7d45d20c70b2bf770a970094a112b60cf8c09be1d740c0ca53f232c90e99b9e3ac7dd22e2ab5d64079caa92cc1b23a24d4c293957336ffde2333b4e6b8e9a46f87c6ad56f7bbcf044375e8c00ac8f778e5cf0d0e2c54331ddae524dc859d4c417a8b97798612729d7c46d2f37c9981cf6be6169a96a70358e298a2f1faa124ee318efe08ef2a9e1b93d470dfdccf345eafd8bb85747c5eb73bd9415a915cf63ce3c67e300912888fe2dbe2bef50832dd5e545c4080045e3e66ab4c9f7fabf932c4190db11bcc855c3d25fb8165a636a6f77578d5488a9df35efa2dc731408cc28f13ec360c310e75d9700ac2b179d557aea685cdb364eba6b6bf3ca8a4527aecc8677642dcce31c01418b252275d537ba1edb61acfa76590f537e10d6737065be8b879934c17d7e0d85d96ca9d324b1507c10e006e9d0374d763d94379f8c6bf398f115cb333cc03a3650ad7ab2b85e48263d61e024e14db842323257e4370dc85cc2800d211522faa8e4f5e64b7e6c7338b3fb9fe2406ffcadeb427b4852cdb8c471123a16eb96897cb7224e7bd23697bc19a71f11a95aae831a5e43529498f2191992abf9209fb59000b691f59d02c121ec1ac7462df0ea8475f5694a0cd0cd707f5f11996c8a6520ed9658e5b5930ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h886e32fd0431420d9e6e5697e930e21f60dd44aad5b6e61df831d5f47dfe985defdcdd0b3469ea19ebe046798da9437a470ba10d6d0f210b9daaf726a6cfd78dbc0c33308a8040d2d6ea56d4f47565ff2a06da117f429bb7c82d33ac7fa1164b41a7e69766f319e8a2e442a90b0a1fbafe9b0770d8774bccd3e2c3436deab54f1294434bc46a56088ddc6a16f57411a1a8c06dec177214eeb501e14c4e843cdf8bc84f1859fddb4f52bf3cdab1cb7835e64930605377d74e871f61621d76ee3cecbe2b32964c2cde72e6d00ecc2138b38f0ad72babcf09ce9e8c66f390825e898c164f23d30cca6b2486c67ce42a563617deea33a98105c54c40b5746b6d55920d8409082e60756b5266ec0f87be58423601bd65dfeb090e535a5a6500213937a8a10039a48d6cf8216f2221407d9d142bf3215712c1c4e56eb6c8f38bda7869a4c49baf66cb00d3659903a7c60a6c7f58ab9453b476fed7cdebe6d5b057ecb2834163963323a6a5f1479b9560a6a1abbca5bb97c21789a2b630a55bea8d7a07806e2c176d7cb43679542bbe31f2702e52f69943b0b3cebcea4dd06afaee5dff35a1bcd150351457f8581fe02f858e862ab7b0e0631c46e3ed5b05f68eb4e4c990e058f6959d85d7ea7bc31a00b549e803f2228c1272003193f5873bad81664d561da0764b5f9b83cff8dcfb9b4db0eced5534f486c4892bca3c8b5e1d31538da61d2d13db411c1b4fe25c1df87ac18fee29e7b8a44f3cab2ca4bc9e80b61631abf84cdd973aa752645e627190c344588916ea7c8ab40e2370ce86c90f74e97b96f7396a3d44f3dc6b4ba3ddc3ccbb794c5c5af3d84c1a26b372df1787bc4be2ca040b0462a2029789758cc0e00939c729388803465ac5befe205fe2bf24b928162578f45189ed88eb4aabefe2b974e4cda9e20204d4371182681d371d0af1330d612451c7072ece0c203c26c3e07f79a0c4cf44870c636023e1dacd462e13862981dee72f92d55842e3e1b83ed77e044421352c590061ddf9de2c8f1654723605c09b058c33344ed7d0b58e2c342f8aece2c5da80a7c36ac0a58935d260d57e6e0a969163a76f0f7047a1345ce822e18db965003ba10717247ab4ef27332dc3cf21cd43337fd385813766d030bebaf08be8c5d7e32fa44a907958df6a580553f2904bc798f83cf1df368ae95e85f6908bcf976949b70c25febf8b46a949af7f8bca3bda94e462f485808ab5bb989683b9898892cb65ac4d13273f254cdd80c13fb3fd303936ea09356457f97dd597f5f3490855f160faa1067c1c283359d760784441afb3c487639fd226e8789f1e75d9a7bd7b782a50338ce3070d2d79a9ef5ce19c9b31a60a8a6461fc72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd35ebbe913371bed6fd02f380fd2e72d7a767283d9c35a9870fa7334ad501e75f014d59b906eaac46e5b85f896cd519724442f900cae7017de2d085f5d5c2a988c2b2b51ffae5519411cd45997385699aa4c28033c27443711f40408a19b5a328db9584f1f2bf19b9a2d49421cfddddec4a67c480b6a22c9410a8d28fcc061a79a9585902d1d69f76d9df1fa73e3e782e6c4abc4fecc4d6c3056ea3861ce8d9cc8d428bf185cf32f2eeda02e0a99f5b19d7ffd6a2fe764e6912a1544042233018717b2159643da19fa3c5301ee31890c0925aeb83838a911366191f86e18333106dc93620b2f656c2a01b4db478f092b2a43ba4d503e59ead8479113ed8cd329c1a18203adc5390f0cc8cffebbdabf28a8b181296ac03bf44cd46a8d1185ca183f364fff91b77f5613e4caa3981d510ba289a7cf1fced51fcdf723b803e8db5f83573bba9cdc105ebe3fd9ab5ca5faa072d03cbecdcfcc7d8293e7e8de65e825d909ff73a30cca1ae8d9c602417300fa2ba05c3ef44902f0886c4a12580e7b39aceff4aa6f9cd8a2813ba0302393b36b2d724317c959f24d0d7e07489ef0ba86aca4caa6268ee5eea9b1e7102135f22b9435e265da78cda1e168e5f60f72a92ec09553db35c4acc725427509c7f0bde193d464f0fdacf214aa192d53dbc8d60286ff8e92e7a71ebef72bfe6f73669476576003923bee25a84cc5bd4a7bc60f8879d3a48143aa119643ba9259b17f6c6286fc8950696339c8d2b19d4bfac5173426ce95328885639d4d7750fd21b25b0672b4fa5a268fa5f3177f103643605cb6327e7ef2c4c14d4b5a8b468a459acd2f9387c412c19507ed3a4161ddcbfb3476b4512d41b90f9d948255994e151929f922507e84d84e2f3573438f375d4e7ab335c93ae53e72ee3f8feaaf5fdd674d39685500e9e37316242426cd157f31074113a003a6dc32cef237a3fa9c1f95047ac2f5eb4d7f441c2566b49b364de53fb0c8e221cac961e867e2c62357b19ce8115c2eaa4534176374e975a0e37b1c266229979ee4f4ce89a8ac33f98b696f8c5455bac2051cfbc1cb27f592a021f1a3957d7e85edf4c35d296cd4f76d151ab35dba99df3c145704ecb70bca436d8fdc9809a0081bb6804f1e63b0208262f2de001a0c62077b34a32932f5aefc04e02bc028cb47865f762975c8831877507a548185d4befdd6a163383bf86c3c6f72da9fb240aeb7253ef50dbc2a9739a3cc809e83fa6dcc4f7aa718222ca9f96284180a7bc71b0e7ca46c9c1d39474170dbd6ff50ca168bc7f6fdafb1dbf5ef6b77d5a87e6efdf7425af6c1758ff522dc179ab46af2ed5bbcfab8159a4a4dbfd4e33fbec004174fe82e486f10782f52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6975a3d608ac65acf1cd47b254b394ac51426db12b682ca4a0b3bd1e54198af6ef62ce9c0a2146ec3c4667c7084d04281e516f7aad53f01b13b1b2ec7a80deaf091efb485889a54b5c839b182e263c9a94944cb64d749356acff064449e2911996fb1a4e92988d97b751f32a18dca414bd7f315c2121ba83665306d359e4c4fff2843ca1f84de4d53e3e09058dd5ba3059c234bde41c48cd09dbb7bd66df878f3b62cf43614f0b3b14413ae6f9ef95ebedf8ff75723fd129772d0086e428b8fbac008319baa14b56fdbf4f34ab3646fb759eb0e02858d8fdf17c1b466e8b14aa34db44adba741d562ac50e5fff39e9edd49d9da38a2a90beb0a7f3afffcad2efed4a2c79398bcf54116fcbcbcec85add05722c6b40203efab6610aa739a2c9ffbb6d780467ea9bf502b1da72916766b093bd1d2722719e6217193f457f537d5cf9c01da7abac16bfe8b838dab3e91887c650422b8680b7968294fd6191c0941f484528c45d866b026424697ee8721592755994f27a209784687d66262b8ba5e6d2131e01cd08cda1d30684d5cd7442aceb8a6c1c1a120552f5738f3d2ac39d6825e9e5be9efd1f9a7c7b6639e6a245170a71275217bc7219215cdd7959ccc22543581be1f2cd190ae3ea813bcde969ef0d44bbea4cc5246fb626ca828d9ee93546b7ddb38e063dcbdda92b27b753ad9a9d9e56b01b4c55c4acae41615dbb0477a017ee27199dce1435630e818fb058f0e6601e31cf4f408840fb1e38112cf14d497397f75f1b252ad3a26b2570e3ab65d8d96859e79081e75bcefce6e1eb3a82a5ea9be6ecfadc6ddf060327057199c8341a3451803a82c53e4bd8fd444c72e701977d8a4342d56c3fcfd78010b65e148a32ce661dbf4ef0bc4871771f5843ed8fb5098913496eaff19072962f25f0ab0c2dfda909bddb1f4199c8c2fc6b124c584f73a010aaea6a794cf8d08ff2aeea9f03ff67fe3ed4f897552e00ca182aa84ef00210c8d67cddf2b9cd4f7aedb503032bbe0db1192df2d25b95b141e24f8e8e18a23a01f99f8fb5d51f00b64d42607273dadc40da3cd2f057d91e0ac606ca851e06bfe25524d02413c2014126b961a98a57fb51bfed1bcb0c787c80f31d23557a0d433af2913dc97a4a6a545acf1bae6a6adba5aeb086ae045e43b457e2cf4a891ea08170a9c91563854422f243731e87957e0882af2653351c32537c2f8db4afe5eafa9ce1ceb38ad855ef2f5146dff4139453a53fe3ebb6aaf6317f5183a1c31f639c759d6a9b195fa67c3c7306db491f55eb35599bc1a07838f84336c4976f6d1ec9c5b0224b998aeb0489cbd1919f607526ff36dd7298ba89243e3f85e14c0fa573dc847a393cddef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h58263eaa0e67bb17ebfe158e67a77fd41b9dcb5614ed2e50de5ab5bc42c16450ef15b6c76cbcb9eabc98e3eb3b26a52ed053fb85471b0fc49c36bfcdad957a9ba7e3ebd2522679555dcddaf6a535ddbcc8266617e369cd9fa35002bff2cb521b66b389a0ae5de550043170f816ade8fe9946d8940073300ea0deede0849cb1f3a5c865d7581d46213604d953059e8734d742fecccf4740a68861930af02d5befd6c22d20da66400cb5fba8b3913fc65e1de4bf1e19d5d114029d786bdf62f94ce1a07e5c718002fe7f379515d235d975cfd1e4f11e225b5f3fa3bdf6188da70ba7240c76d9d17cb234e7b5fbd67f4b21ad8a7e9cafdcd0a5e9bb2386a57e54dcf2609587027ca4feba12d4c464d6718d7d251d899485cf483b59ec0e0283cb5b8d47e147e70f7f4057ecb8bf7d70f4a395696b514e2118978bce30e9dbf706163b0f8334b13ade9c515c2dee2ab76f143e3adef28396d258627ed9482720241cb0fd663c44c0bb6f8b06d90e96dee746292a156a8f617142291136b068ad28d063817e01ac2566f88531f25e9e580df6072d8df22ff9b7d4c9bfa707c40ec60a7350b4dfeab22b953280b34394e61553c0f58d05c2320723a7e9c87084756b804d95c11a74f6fc75b45b6f54f80b2cef22961adf5e5e8069b641ab0d6c2977d2337f59710d5d77cac1a76432fea8c9aa50dde009ae40aed1c02881462ef8e4ebe0b453f09e429f69b8eef3c71a79a56694a5b84ee843aa70ffc3c2dfc290259067b2061fa1f42602560b4649187fa3faaec05b3f4145bfb1ceb24f2d1c8bc3052e870bc7fa0375bd532d8a87fd629d960e1e1316e314f7d0248bd80c87a9ee7f449a3f7aa468af0db9245181b48f59f2621b96dbe773d4f20408a866207890df3fa02ccf2bb36c059a8c886a53d1917a3cee63a3680b35f1a85a60c28968a1d9aeff75b65ae0560a54f7d73239c56f4af3d3621af4f8f2df23b5b04771fe39b7c665055ab9d47df63825af38c0a6590ecfefd35f9fed43574619db73614b75148d9e5f596201f6e0760e62391ee7b49ee228f30c61eee79e68c6413562b77c3e6c8cb2b6f1b0898352c91606e2d17f90a02d36a308834bb5757cf5472fe50788f3727097f35d45f1c7c87b9382e98e82933da19633855d64a9847e7a10b04b7721b2907f5b1ca5b01e2c4f3fafac0cd84c9505c21ac70dd6df32745d3618b519c451e9f36bd89ccb3c92d912583003478d8e4dae59c05730410fe68bfdcdc83738ec5d80dc149944a07126a64a9d082745b9c2f63fe36c65ebfdf8ed8bfb819a343cb8d9b686012208387309924567f133b3096407a4398c28615e677eb5c00748c7ae56099b2603453d38b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h305946ccd345b2f8d2499013ab148f6b8359c0c3f0da7ecb306b538856d43dbeea5b6b7fa3e2fecfa264f0397762bc2db692244e5cbe20ac596223fc5af88d69633e016ef8d9913190f32499650f86bde138524e4103099ef814be824eaa49046931c2e2ba0256bd2a78dff7d737e829580ff2b14ac077558821e4c0c465f448097b3711ad34e7f62d1ecbfd6a94d8cb85bf9ee7f4fb0c2cfa42665ac9c6849d0ef9df466cf7fdf5ae7644846dcfe2a5fe6186eef8fd23ac60c9b4756358401ac79a0233d48780c2edbdc8bd12048dcbb30496501aee207a01e0495c2cf939100aac3dadace5a8a1cdb26e0a853e7a70555a4d97fa44c3ce2d032ff90443d9778eff7dd257a6cc7112b3bbfb577e9c41292be7cd17c768428d4c9f8676bcd6ffe589d7a3d99e910c79f896ffcfb81450f040b9d941ec6b3b870db6864674a927fe2ce7896a10e0ea6c0af1d403fbc01ca5c09ae0d60a741ff4baa8768fd63bd3a450044d52374c4ea7ccad59e5497de2afca8007f536911ca6103fb33d67187c56f0aa9b6d71e64d1e36016b2d702d8a333f69cc49dd622a70204760413e39ad89a0590b1e3c0c29850a506cae7edc328233100173016ff444b72258fda440a3efb47341e0c6182cb2a35684cc82c8b3e29753244799f2b4b9f45b8876aa8b623e25b936effe1e8f63d393962b5936d011b0c6f6b5eed5bb1da9de4271f66baa41ca105c74c1b798836534596b80f07cd39ec2d2b4d1f657e1762ffa034f4c2d418fcfcf2acb874feb37e684ce91b5d592881ebc6a530468c5b75963728ad58f84d48822d26c84f5ce25c8bafe29df12d14d8f3fa8b58da8c953f8a7e722ec3765424d7de7ce6e271643c5355c4cd34817ec59ef158b08c168872d91f8b186298c85f9a010511c1d228ee0a1c405a609d27ec8f52e037ad534d8766ff8e782e08b728611e5e1b642cebc995a20f56655d22dbad966c475c645756cdc7e896e0cd30a34973376058a73501b4ada3779d1e9aae520cf8777722f8d8c3a45b928a61fde172e4e0f1c517e257bbe3a6626fbaad78e3cae12cdc05c5f987dfb14a7fbca8958031a4bff052c2040f936f95176aaed26fb638767363ec31ab14de25de606e18e202eef31bcc63a88ba5b08c517200037e12a82560cd612bfc5c9dee243edd20f400d58320e18d3212c0b8c0c54472529e84887cdd5071f8258e3aa558c5adf91958ded19e410b10e2a19a9fd0a3ef3e7154a0a06cbc1fc9ac7178367744c237ce7a5ce8a024d7e7ca05e2b773cfa78b32a9ce2e325f5125ba277a0cfcec63615c977b2fb118a6f1f681ef30c6af5dfb54b68b0b4d28aee67f6105b516ad98b092da0e288c94a4f6679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf1c80cb9059b3f101eb272163cd5acaf400f0eb53c3bc494dcee3db428d555d0773fcc915b094f9a16a9dcd43de054201717f6f03a9e6858cda0717aad61b74c293ec1644dc0a910369bc4a183537f14345b92dddd31aaa14a61cf95bfcfb9c4501ad03c33185a292b4d751f4f9f76e07877c1de8f03be60c6f3468ff4ffcfdfb187cc433da49b9f4b501adfd0b2b6601f7d7b52db432ef2c4ab14ee64d86d6679a879c64e0f4ec3f3bc3a746cf84474162d23d8de7664c6c242867fb76ae3b3a5499bf64c4695a08820ec0aa88366333d785efcad2261f479d45ee700f528b884600f2276befc8099b19294b868128fff0f19b541160ed37f96dd40d724c7215c48a298d824d2dc4aac48b2122d6a83eba1a175fd564d5a7e474258a4683a8d0f822ca4621a843d8d991576b533d74eb810928f05c6a972ad1bf7aa8f5803cb1a9d9bfd688c66cb932e54e6977eafeed351283abfea17311a6a725b8a7d908e9f8c660be313c404cb88557852286266661d8ae0180636b3a646ca2fc39e22932db1453ccf425a239080e9bff5c99dbca92a7d0a0a1dc6ce94cd5c04b5ed60a146f796f2b1276577f884c80a5c9a7ea5778738b0ffda1f81db657570ddff5f792047c4522dabc0c1b3580d009b012b301764bd82d6118f7339ad902963bde742fbf57493203897a2b24eac7da1a716f879e8844fec0c9dfef8a7b0f4ad5852067552ce9a85c7f5ba00a7413c90cc9cb291d94462d038b2a8b4ec169113fe73c93d1f8b26dae4d82fb7fdaf3299566fb18f03bb3c5d737acf2686f32e0b9986a586e4a5d881399f1689e5d7fdc96e0e5ace1e46b149fe3f77b557cb448112847a261ce8792f019729edcdd8877d7dbb8f999b09347c2a5ec3c143bb99e8e1838382b37e0a1e849814b043442670ebae5844a63633ae69d2d1a84928f3d144c3c5e3a7dce4ce07f2dc1c37dcb80ac5bea58791f97ee58163dd657c00ba470d2f4b606d5f6f6f2553c5088e51eaef854e29978fabeb73bca316d260bdb8717f8e52b711b284636a3a459f7fc57d358fa0acbfc5363c9e0d74be809d8b224736174142fedf2b99a0018cb152a58b4cab91e84f27ade75d82e11ab1f8d2ee6ad9e78bbfb5c6cea720289e3883d84a5b58b2d8167396647443ad55be1b02330cff06d0a7055859f703b31b6e38ffcabe80113e8c924edeffdccaad9aba618e1d27f70b6f5e78c440634a6619207be8fabaf29ab1846b706d5d1815c201497096a523cf7a70cc15391e1b372b10f65cac7097a64db426540ae9aeb7a2729ec8120cb923d833cc8639a5c4c6373e9213c753a5029e67dfac75d8bb21aec39444bb93843b4649ef42da65ed2cd9eaee7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb09029531bc3da5e3c99d65dacf59dda3f7337e3dbab60954918a86f2bc62f2cf6c6bc92fc4b97f4f4a20192e45fbbbc833381a31adaf9223b9b32b57e4967195a84a83bbd66e03b9f6bbebef3cfd5ba0d59519e09eff20c9876070bea4fc82d4839fc8b980ade2b2a5c04c2c6d4c496dc478fe5353425b49ff5194104c3f963894437ea90c45c1a2a0059adc0f49e6d008f5f849bcda8ee98407381160a97381fb3712b3611e74d74b586b34dc336af6d1e1620d85cefcab5153185927bebb5300a07f293deaaa5a02436b445868688a3b463d5fdbe1c5d2b701b08385e6bc4551b276d6a82592a4e1c006ff5a783c2f071f3468dd5815a5e7fa88c068f1553ccc7828b8b6c70029e4852d37de102c1abe3209589d887d5e2e2f1c4ae88451f3fe19e97c600c74f6182d88e4558fe4ef629a25e5ed2a6f31c28a445ab8d7205e8e2f951c0fbddbe968c922d360c52b961297ca28e240fa5e6628005b80de0097b6dfdd9394d7453800c4d42ae4adaa87df13a8a868f2da1a95c6e01083b37d79d8c2fcce284f7f26c7985134f826542e6c7f5c182724ac0bb26641ddcaa4564448ffb23b93ea3b4f6758ba39459e03e7b31997774a0c80709a5bcde26686a1f19a615c80980cc37d508e5a807636ce21a5f6631b199be657e0455b00d4c2dd6b77a7e90636044198607d0a6f15a3bc7fe565f8c5a8081d3aa38644aa78fdc2a7cabe6a04d4e9f0c28736879afe9893b6699eb42c78fee06b7209d9f19222104dd4334612c00b3f3ea0e469f351e5dfebcd9c4557047e8fef2d81a55c5c949b63f8b0c3acc8da3cc049b5f976711aef5e308d9768c1cff68b6b9b4459c96f1eeffd21464ed88145f3601f7b027d7268b1a2125835c19390b490c802dbfd91c5b0ebbf702ebed197a443635a2744c285987c8359e275ff8aa272ffd437243d4e718eeb7476c09d456d01af32d29d0c8413ada9c9ffc9623291e35a4b6e9cd9d3a1fb45657b7a480e0614b93cc375eeba6c542571b89e1e3afcc5da6c7f30bde055932dec59e169cc9164d9de93fe52620aec261823b7dc91d4cb0614acff776aa1725aa15d0f24708118a5e864298296a0d76c7f7335aa3cf7772a27b1ed04b0651b40f6a83074d1f031ec886b51991330ebd2b063f613b0d35f3b5409d7196a98f944256e336b0aedec05bcbc5f02768508c63763ca350c114473e4c22c6ecd3b58c4ca1dac5fb1b68a0736d907ff8141eda896a3bca9a8ac3b23ca8deb59216efbae575bf53d053ab610f6aa26d0300db1a1e51631a98dbda864146c9aa6a56a8a4866e8856e0ba334f1e478f76da10346f222cb112c6b708de5e21674163a07c34ecc5edf45b3023ed8e01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h62ebaba19f0af8a142993016231530fe8c489013f415aacb7e59b4771ae35af9379b5a1da9b3c9d213a09afcacbb363901be8b1d9a074967fcbc7befec25ffbb9569a9317f4cc292eadee564f97a6bdf175f5558ece715660e0e255885330ec135f0b8bcb6742a6dbb9951d3e554bc74f05daa448bacd489571bb37e9900566a2bee6cbac9618acd9e57a8500970eeeb6a8a28e18ed7b9b0078784c140e3649cd0f379c6a98def1504148963c2a347592da9e1e4eebd9116837bded241e7225568c50a2407795e8c92039d6d7c7f95e3d76fc9e5744e9f121e59981c7235fdde9fbf425af4d49c71f26f69e902d38a050fd10283b9f120c5a1619638cc78a1dff1a7b5d591bab3cfea0be1fbe59dd46f49dc03508719df02912eee1bf14d23546c5770b810223fa63552483aab395a04769099c0d2d6b1922ad853fda7b2fd6f9be4daa8d6acd158a182ca067ff23c6de99c998dbeb2b7403ea9ae6124cc00b72e93ffaa6b5637f7b3038cb73c0495a363a9506684701d5d7f0a8c8ae32b00e69c9149120e311d20e5eded25f28cb1c35978b68f1a2a6671e4b573ea6c03d52e899cf98bf5d0c0576268c200e9023a820c7535c5d6b10560f366447a67bb1081f59d7c97548120e839dbbd2f50231e5599ffc75519633458dd1da7926fa6722968e0e76d6b44430b66f1e8302094cc075184e5885870e3621a0641960eadc1e7c1db258fe2682347975f62d60604be096e59d911a014788800a7d2715b23b39b3921db5e16d6d532add9c05180abe7217d060ac737c8e988c66fa8a7a447f00e32cf567216706b27ce1ad9aa031271dcebdd60efa3e759ccfc27f13be379997cb863e3ef4552eed3d1b2dabc9f7f491bee69d27d2ee2a639bf3589b4ee4743aedcd1c31f89d76c3f9606845cc9da93f8a19456e9f27a5d75bbfaa14baa93a84cfeff0af33420fd50f1b9b923ca6b2051ce9fa870f3209a09d60735d33fe4b7550373a7631f460269dbd92e13e3524c46cb3d4706db20d6df3716d06b76ff0f516c08ce2256f8d5ecf43ce89b0af83c31e5106e9bdb0a076f1312a3dc2f5167a2c84372400154e1b79b8a7bd6154004d6718d8bfe5b490d4a375bfa60bbea87618558af4e4ba74ed77e6a422c2cf9c3374c5bc75ff917228ec2393c17c4565361c3383c7b0b74953c7e90641ccfefb7515aed4d2f6dcaa5bff4b9eac70fb896319822afcf935bca3f79560a475583c21c64a1dd27105edb57247daaf74ad61dba5839b20b977f67dccb5eb2fdfc562f5c72a2ecf24b33b5fe88751f4904df3a8d6d037df06b1e432f78e4ebb6c2b840fdb1f9b5b00f85c3109748a307830440ba84dd39caa7c13bb4b92a3db0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb9ab1d9c758817cf979d5734dbca40aefb7cb4dd3cc38c9699132c6e30c3721f6945510fbcdfb046ddce3aac0b9e841a0a1fd37daba4b1753b3a9d7f0e2cbf6e00565b86882b359087d184493c380bef4139e24ad29fa3aad002158894bede79d4b16cb285d0709089fac509af52ae579c4aa56967c454fc290de05b99346d80e27cf09f172c59578ee8991849a413a66dbf02b4598a27b9abb0defc13ff4a3007e58d9066d13d60c0940111557c1f6c7d5fd50ed334a17b8b9eb4e79a213ed8625c881e7972c950df5e56ad4c1f4c7fb1a40072383d15d5ec21326cf18e99f008d5a1fa287ee50b51fe70da477a8dcad7dc2fe079dabe2db53161709509cd5de176d5e1a24c54c5611d847a892ecfc667c47077b38c9980514ccc315a0f58176417a8a5710105ec8bbdff5a23de8231ceb9625cae05b155318d202760429bd7a07c0526369e11337105d0fc2f50954f12d7f231b4b99b2ef9cf43c247e319c3a25ba98c27cbdc9b305889bb0c9eb8105769b41d786d5ebd9871133c226233e069673a8d8fcdb8417ec9469f7f9851cacbd23cc3f3e3b000dd721340fc19b54690728ca08c160ba69da50b2daca174a24fb00fe3e0baad4efde554ca25201914971da8a62c69c7f7f4e2a2d98c71f3c59edd5c6598123bfa332f41d56d0135f11eedb039c32daab4ae62f80452e4ebaaea9df16fa90011cda1735da05bc8eb1223270b0f837afe0bf88d4914005fe9c15e39fb08e606b6368b962252c707babb893f4d852a0148f49957d95fab440c04cd63360a96bf2cd7e3686f165563a3c36b5d88bd1356ae2a9a0bb9ceb9245fe30ceb47d3853b6c56c51e4a23691dcf92c105ea37c9f495cb152188a277a66130ad23667ea5b3ccb8eaf84495e9921190a3c073265a130c14444677f4e59cd782cb43d6ca75a35ced9ece9a98dd7cca58f46287b0c0297346f52ee8072de08dbaca7ac8676915c9e745e5dbd20d6dac6e06d41bc72791a008b9bd78e2169f5ade831418093d41e237ad2edd7433321c71d5679f7982229e0814a654f969b7485694da02b35228c039404cb0a6bf8eebaedc7a33a35c37d20c4059190bf8c3d9bc3958878c964cdde76d2b353dc1216fe2625ddd468ee093a23f982e241fdace3de6b213199649142ccd5d6ac3c79260bad6ecb82aa04e13e3e0eddef4c33469eb0c4f05b16e0f3e79cc9214ea2dee7a5180ca28e1a798945fe29749601f7766b64cd56ebfea0ded62b18f48f4bbe84708f4e0a5b4a36b99cbcdacb17850bb657eabb5cd982c4cec300fcd9be8214fa64df952e5ca8f761f09f3509c03641d0a726031a7d865c9c51af2f2cc10e93c89244eb240a32257ccd351ade9f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5dbab084a4a7c351253c1e026b87f058b3b0e53bdda69d5a055a1dc252b31aae129232dfd9d45371e51dba2ffb89d1873a5f9688efe72c857913bd48b8e0358e2df85c5599128ef257e7de5e7d6cfb841484b3ef084084d8c0aeb7e7d3c0d5a781f853e676830c7ca85337080391a5ddd972c3a207d075987c52ebb6a0a1fda758c8f46814671e6acd8d9f02105dd8daffa41fef58af193379b811913a3c9e1c8cd2992fb64db7caf8d90981e6c929b8768f63e7a3e527c35280f4fbcf245bcd705cafa5c4bd709a01e9676f35d7e9c91061d6e8ce589414c40130c4440482fd0418776e7b7f35a307aaf98d48e1db5c69c25fe35b00b6d70901c2974d1d1732b343c409dc495eda86463a341b89cf3323f53abab37c219bd42024ea113f1f947f10b7ae44093626cc189953ed44300ea91905cb360bb71d36bab68059b8440b893b9baa23acda43e37c34628a6aa685ded568e9d56d575f0aaed92b716dca1ae39ef7746b1af45d45a1ec35b8647d553528a40aa55f25310933e60b51c492ffdcccedc4823979f55b4485aa32bb2233353a3f2564b0c75fe52e885c351f01ebbf62f21ec9adde3e9e9e1d1ab67f6877fda7b71c88eecad8ea4dcebe41eea117755c35c946e9793ca7d1ab91e77cb2f6d43c7511489484448113b72cc5bceb7c6cab9e81584fd28dfeea77e073f1a8252fa36e3b97004472049a34cd06016179a4ab5fc667c1b6c1f831df90f52490c230a2349a7be2be6d6e2ffa7f3d74d69a05f9034da0a2404c50629b68b1ddd665c462cfdcd56b6f53d7e6ef8f424970568cd21b023f671829712e002a00494dfec0a55927f28d3828fff46ebc3a000284503e8e0775d92542776386bf5a4ceaa034648d4d19df2d02bc1f30a761f71fc156550f93839097b369905e50c05215e1cc13a68b9befff64771b247e2f2f02324859984c044ab115528d98696e19ea35adeb43b9617e271c19f2622eef977b0e0431492d41cc5d2d0ffdb990f447187c597d07cbbfebd7b508c0413e3993ea7988541f1575d37da4cc3caf022befc3359add5f379cfb45a8bcb0d171d387758c59fb96de7f4b26c60aeb1dc6f7d02fb1614b36418fbaab06dfb59b45e079b2e34a5a55a73bb6d8f2acad2ec3477e540e71698babd8701a1db9aedab2aa6eadd6d7d6aba8a0bf63b784b51b4c5a54934d2f8d5e67697b5999ecbe08c2d2ed6dac062bdd5fb48a56a17ae447c459581424d4015ba5c0e1eef5d5eab6afd57367b7abdab95ea009da7efd73c423d1c16bc400984c2e5e40d80ca458a0aa24ec9a698b9320079780e573254ede19ae00d50a780814623e3164e3af51c4d82d93c880782a201e1e05fb964df3a3a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6d14fcc9e9239ef888ba501e0b9c3cb8676a1a7d8ebfb2fb8e07f3adad342982a1f3c799e85dc1681f0a3f337603ea41fada89624be48872e34234ab1f2246e931415a9b8c3be366830a9769f52f94f480bb0258c9d37649e8c6bef7b7c42dff28b568d8e34c3d028ee2c09e9f6aac150fba50e4896cd466ca4ec283262c5260375a25fc38ee11e0d654c399baa9b4d671eb9e502adb6f70148d8ca0ad298ad287e14c794755c666847dcffd9686dd939d82bf13fe1c1ae6e62747cb73fc9f852d936897c59faf479af3825b14e6dd1571979ace2f76c2e755e3ca449e38c251e4a3dbba353dedd1f275ac27d84c32e2f8e25d84743fb5ea51319e6515cde8dfba8f7e2662cd1023e61d59dd57fea2d69861bba109ce4dddf7c03cc360969ac5633b4714def7f6b26008223764c3a92ef3be95ae39dbb1824a1a7ef070a1237824d4a6b8bae4911b5547529bda54b9c34da76214a50bd82ea5bb7270cc712a4c644aba521f111a0d08f487d464128e7e51d6226877f38c3368639d0ac2f4c141e301590fcf5cb0e2ff6f289b3894270cca140d99c4495d9c308ad1d539b059a01513d346ec8f290f3f80fb36f63dda39bc01c12fe17187ced89c6396ba3a00cac2b5fa0a3e123b9fe8de40b5a70d91cd8709c594826dc760baa087256749042500d8e49623d0700f16d2d323eba4c06bbaec11cea7390d822bc3373557c1d20a0cf033045b29d12fec63790f00a8815c4a2f7124a9d1ae3f8ef039d865c87a3914193224adb54cd25da80c63b5ad4e41bdb86aab7f0e067c770683cdaffece4f23a0cd18af868d02ecae47604b8ce56054720a47fc5b8f0917779c2cc6c203d8c574b5b1f38776be7d2b5681fa7143a2a18f805ff45e2787c3d6eefd3a97a2247dfb67ea7e962d7e34e354321ae7cef77411116fb61c6b3334dcbf38b25d378d2df648036761bf21c7663e468b0501ffd4e7fde78b7e93e5a8befc91e1bb83a3a3c68cf9972af0ffc376943cc53b05a8e7961b40b6e22e473f2fd8d3ca95c6ab14ecbf7715dcf144f5693edec07cf6ab59bead516313479f2390d4cca63c09a5d4435e0c3541d161d26f064165a8a3ed3d1b7760a927219015fd7e25955bc66751ad680266bad57fe782325fcc3e29edf6e52b49ffa094085e97dbeeabe8bddee53ff59bcc507ce988792996324abaf2dc7d3bfa32cb0ba699baaf94691aaf264f06cfb0db522da71ce8099fdccec28e4fe2f1c740e764402aeb141abcb0b6f7095cfa2fd2a85452ebc12e923b107e04510ddff274aca6e134e651767aa8439e81bf336eed3577df54a7f8825db47a31ae9023dff4dbfa625c23b7ceb0906efa60c758827bd60ede30955655;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf12f0c3ee49a61abe6a6d6f298a2bcf27d27e098d44089474d9cfd168dd6396804372ead3ccdee94802d48cf9b70ddf3870700654ef3d8f41f77d232e2fd063b588ecc0c7e36604c4ec0261ab4673e13904b9ddd58ea95fe0e50af73a2b21f50397ae24fdc925442b77f2d827bdf091c08186f346b1a2615f5c40ef5e471c5bb8d8c6fb74d0b9424d2ef8d10b11e6d092a77173b01bc86b83329f2df1874713b8af79a0679a7f0cceafd4c4120f0daa417d865cf80319eccacedc5a891e861245bd74f19c97a44f4d4a3ae9bf179a514aa0af0d03e30842f3c4bfe1f5afad553c4fc9c186b849f30837f2ee6fd8f033fb77fed8f4e66ed6aa553704192efa4ad8dc77835ae3a07a53636082b8e02a8da347276d11bb0c2b624c323034fa0a2f8f5b6ea542c6046ad80cc0161b03d19c59b7a14c3b0925113c0ecbdb415cfcfece06bc9b44c9a6dc06fe5bb210ef7e7509b81593903cdf61137a5bc614b27d2196d40fd4c51466a5f1bce23c282c14fb3c19b97eb9f777dd15a6b7ee944be81cee724cef97bf528c17778c6f5958f8cc58316f056c23689898c581e0d1a28eb120aae5640294f66508c74e51f155e995a6f7226cd5ca2274d5582a01f0378bd9544b2c189ed43ad0d38593b0b0420881a6f5d839911bf615b9f40c7f222244312d7d6c70b18e982bceb2f6aef3c79ab27232471a90d7be74715e9c243e0529f9f1e7254e84a814795636a49846f3b366d600a9a7e1d75f474e3cbd1c123da8768f5c20f1a1957fecd91b6994918ddfa236022163b6aac3ac6ab1f02b516b2e9d557a59597ca82e27c7418c806c9cc21b00c856787961608ecce8e37214135f81ed58f7688a3dd661a182799d8beb7caae01c1ec61f4aacefc380e1411f140670b4d2c2a3034f7b5c798dd16b770c65145989db7527fa958b681c6c0288b44e9c0c41ccb70f3d99dd2376d613378768a64ee0dfd4e5d0dfbbb5a0c01f7febdd04417d34d162dd00dab951f5a51ab2ab2550e5cc43e92083e39202540430a0250135842f06fc7dca41757570e7516606d36ef1932b6dc35cc90a10d2803b0ff64a9743fcbb782762b127c8214e94f9044223cc95003b0e55e1d0e8d3ea29a7d1164fa022a31c6de3353d417de4699e03ade1939754641735c2135e0cab86059f084d79b2145e43525fff36c990f2e89e5af2f4f19de13d503cf930e6f19a8b17996a4d48c998525d5bd4d2f81ad76788ab6dcdaaebafa1f6f2e71e109182ace1632613dccca1228dd7a2555ca6211ce0925f032c9581bf311dc8d35a22f2fb70db5df6510a5193cb0332cda61903332a20e2163f864702a8336ad75e602419f3b7c6d65f05f74514a7e320f6ae7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h7b2971755402f10c777ab21b7b5d69aa2766f85fa8a5a467a5c48ff2b5251e54ffced4781a037c57c499b00d1fc6004d401e145325bc657c3d3d89a3ee600fd9db5758c549de9c4736a8c7499c7f0ff9f9d5d44cb372a9bff838dc5101500b47b49847a9d7399bb8143dc01e72ec21f9fd37752a4b111c917d38980945054cbe27ed14713547025362de1f6fb695befaaad192fff6d2a657755024ae524d027f0b56f9dc5c1c47eb78e0be7d1dadc423014b1855d651c5c114a04ead9b9857519895a684a1599120d4c17499439b45cba558966dfbb5fc0926fad910c4a8e39a925a4f65dc7f4b19ea7615c665412848d8ed263534d97af6cf86239a0c454874cf22bdb4b4ef2c03fc070781146051c6fd7e94acf3a1ca78c779a7196a0354da1bb94e263a0fe3a16625e345821dfed948511f41f6c6cea56b20007fb5fac6360cee14914d92f0341f03ca6b0af7f6cc5f99c7deb9fd7a4bc1fbbdc0cc9d928d1f272e213637f2b9daf65808825c53a3efce566c44319483928c6d18f0eb493b8a07d4c5e5e2a0297c515016f7c37c71f522511d03f44927f843ced5ba0d2a838182890709e0ca0f9dc9b60b701122b67deeb1aa75163229b9ef4ba667577c9f695a77984ad8f3a05349445f6fdc06ce5a00cda34ecfef0b6f4909c0cf3673bd2a6b24183d6520c594f8f7772f95ba8a208bd4fb157602eeffa49e6c1840737c61b493e780ec10348e58bf9a6062241efdc1ce9652e443ed5109b5842e4df9067388ac6aa0c2225f367233af4ea2d51ddfafc11353a12162ad570e3c5270f26d234e14c8848e3252c1b29c04a2e89ccbc91f8170756767a0fee4886b053f5664d4ccbb4f71704cabac2b61323bd906e7f0c3f6b1b945cc562e59d04bf22ee258fcdd73689b6cb5e31eac6d417189fd0c350ff444e76b58706846346f9c9c1cf614c024207abd9023b08a7d585349ca031c776102013db5123e9f41cc0c956a7f52a9d9c63ae2bf034e02dd980c4a8cd605fa5cec343f2416160bc357e535ecc08ba36b5fd11345452ee08ca0f2fa2c23b13b58d516d29c028541cf75407821000ccb4f9901c42e7c2ab33a8249d7c06b2b1c47d7473a843714d5065125495b613f1098ca0c58536f3a83bb7634c6f3932b3ba28624c5b954cd907c814cec6537dbcd564ddce730da1776f51f39ed8b9d39a4f31042c5b8cf5114a5baf0d61ae8181e8eb142dd311cbc12769280ca4cf9d9b9e80fa3451b6271628e177775feb596a1185bdc63df62da186ef6b484b59841b4209d58c0b4f021babdc8613712c1d96a93cd6e1441395cfb79d32039a9f93db4a80592c22dbcd1f21940b707a5fd9200060991accc73a440ead9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h29500f0af1f6d6f6a2a8eaa3fe140f092a99cab721f252d3b17d4334312dbbf3f39dcedd89ead325d1cf53840798bafbd0990d5c5b40859c4b25972c380ba6a5049683845e9e31b5a1271922f31e252e13da08af71ddb66b5deb411215bbf5d3a5fdc7c3100cf6ffe12752a5bc30e8d7e7b7a81e30669a2e1ccdffcbd3568e8beeab11174c278b368354e5a3fa06c260a51a87b61132d2e0941cfb53569b0c9b82f32391cfaa1b633ea43f66a629de12891ff71393163c14f4aa4c88b190bcd3969d7619abbc78deb3b54a28fb9047876c0ab87dd7509c7010c96a52d53b9dd6f1e090ae05978a061b378cdde369c8bb52b6d4cd879ca2d5cdb0b4330bb7a0dfd4968291a3c8251f2c213574cb3b2348f809dc46def027ec8488fcf312f86025438b11aa589d7fe5a128c05dd6816ed70cb26624df5afea29bac27f1b0d76dc2403c4172104509312db6985b0fea4cf08916667f14550ecbb1eb52a982cb0cf9bd84290bf1489e932d359cdfec5b56d4ba7dc758c6a28523b2a925a672d5b135e8a5cece73a35baa5525fb33705ab8a6d2e6b95639a66363ddb311bb3eb6b96f7c17c473349cd861dbfaa5471c81246ba696d5cb93b7e5c98949fe49091ca7113824e959cb5f1f7055566e87f8971cfae7fda83bab23ba8574395ce03ac157d8cbdba215f293c941bb4b799625bc2686d5a2d34df40541618ed4d139f1ebda5f2440f61303cb210cf6f61e74b3d483a36c606669ef08d4a3a8b191147227efe8a81e6074dc7e5855963bc595c7dc14f085059e5eabbb2f665045b2b10038faa80ccdac5cd29911aa7fbdacdb6e55e695f0e50ed16f2f25d97e4fb7b8e630de5a6d0d4f7c15c5511e117805964fbd19cef4a7aca04b8875942ce94d37c9e6fe146678bf02a6fb8e0fdfd023a9879b09a360f456c2fcb2f18add03f980931239328ad3878c6ba0821125edbd2300ebf5deaced63f40acb262ca8d5b0d481c454e0722fae9cb1b92bde87aa88e7a5ddd70d65d1cf759ba12972ab628d2e44b7ab4662d7f02410b2e362651b048c68667136e0e72628323ec63d88cda63b06a363df5dbf723dbd170eb660d3dd2f088fa0014cc0fbc5c06e4c478e425651b4899ac84f33d47f992a09aa6d5246311f6b642ca068fb2b004518f8f1a54e9b28e4e90cb43895183d527273270fee0db28772c916bad2c725b0ff586d2829279fb2d6a7965ba691cb5431bf29906520d65dd82709e7f7ea1ed36bd4d8d52f0a4e49c10aa6272f88ec03185c066ad226abcf322694411d98ff6957d3e32f08a9f711058332e6b356c4948410c34523b1672b34b23b7c898d0b15fc9d7ec9780551f270bc0e72909e77bb6d8cc2753d98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9ff2418eb6cfdf96bdb93dcfb3a7868dc2bd2694f5e888ab657a414051bbb109cf4fa96c808aee05a376dd3938363fa54170c20445c1e3a54b25b075e4f47c99ab4322e59cb17bf424b8cbe1c85cc72393d7be24e3a96c5fffc47b73513b1cc0cb8338752cfdd0c3942b2a313aef3190afd3d167e04a594123b5501d72637db6fcd3f585ecd39e25a960862af9055420b9feaef8bc0377a9ec8ebfaf42951a7220c0fa19ff74ce913e4f43bc6f9a8a31d3669628652ac096b3874724f26a8c76e926b0dff38b46b4d461f1ad9726de67eebfe9f5f731743b75d1589ea5bec88b4de3d5135eafa63a97a69d9d528a7b995f4368294267d71d888f46544db41c39a5c848d59f037ec905db1cab809daa0a1522a2554960033343d7794493237bc53b173cf3188305747b4cf365c8cbefde73faf9250d2ed612e1d80ed6d4baa817ba656f74f62a003ba759dbe717d7cb4ba8e01c201ef07b23112affea28f44e3d9b24563cba2311471a39457940702af721095e7b81bcc2eac8590f9ce5bad78ea586e98eec33be3ba6c707e671cafe5761dbc34bbf8e6fce93a542082504200bc91a830e29e6258026dc625cbf851e860c3640b54e6a6d9f3e07af43fc24ceed7fb074a01d8e77f2d3907726343924ab0409355464c656f2f1b962822b5d77892a19f8b572ab2edd7124a5102da7779f59179ff45dc2fff1755997ea815f3244f8231a2e7ed498bf72d4f346b1b9d69d30db68fb4399be717b588f8cda2421d4ca9de83722f8bdbac4a7fd3cef3d79e23ea6106d1b2657d38ac01d8d83a6d3ceceaf2263dbad453396d913bb0563eefa6a3401228ae8d93466265989ec2efabcad4fde558a3eec30c869522d76d8fa536dc2d9f176c85e9c4629ef54e9518263966678a4be4605efc8bc01bb48775a7864a8cdec0f88dcf149f2fae47f26178e455bb851918327201f3f6e258b91f03b18e4758cc0e360f85a08c91559b5e8a42b9f4e6f699e4222fd68d4777b11b1ccd6e3eaf0a75b98782acc95c5149fe674d743e44ab7c72ceda2060e8abc8e6b281a17a5b868ef66958c1dcb81455123c565156311a8e2f80092ed18a064de9a992cf8426c36e2077a6f6369bd7554ff9568d37c83ae71f8c84694775857b1e37408b4f2f3b6ba9d51d2cfca7cc4524fb0ca3d8f53489c08c0aae17d83fc6ee54fadd89f7a9c8303b97d61fef8c7af726b22ebaac39e3a98bd402ebab1313793008067c34b57e17561f7938add038f676ffed49d90415ff26a8c2768d06dde29bc7c06f4ddf05c49935fc1bc101a0a63fa9a1d29197d8070f3b68173970410cf684d00a659653b3f2c2ecdae815c607bc03d835cc148ebfe463cb66315;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1c075128a9372fdee7d0492c3d70fc726c55a4b8a78f6a61589be00fd9c61b718d8bf32a8e7c46bf5e034837a4f62e22989b713565b7bd050647d796bb6702f8c680bfcde29a003c33acd8070000dafc24b7227ec343a2eba4e2dfa54d29145f16322bd7d1ad3cb35a3844006059d226d15a1831c89c9b559547ab116516dd6ebe574bed67f52b8d99b259a1cd444fdd9b2830f684cb35f865a4752fbd299734f4d45cd35120a831ce690b8d16e1f046e6cee1366bcc4f8c2adb2e07f050f820e1084cc0d6de842424d69bcd68e3917d19052bfbf79d80cc7a560ccc2815a8b34a29884d9f2719f6f0c57ce14cd508bb08454ed44159344d8db8ad51767f63362dfae887223baa05dae99d540886843c7d50bd77541eb38205acd6425b78bdd070027d1138fe2ca4bc2dd86cb0e79bd1cd6fdf8a726bc0ee513123d77deb687b7bb98e1e28ad7992f4d3703697d2e38ce7ee3d0493c547ba96d5b3a82399a55864bd06451ef612dbbd8d401baa1296f9adc992251baf682aae19105da0046b9765c87ef86ff05ec84fde47b380063873c22e9e9087d7d4fa6bc42fbd84c068a840cb07cac14237ca2b4e6bee76692faa7ab6d8623ffc9a1d8f9614b2e833c6adcec7ffc38110aff907eea49457dd0873a37c7dbe8b1ec122c1293313615957425476f0f5ac660cd13822d793b6466bd0cdd866f624502e0bbb04785fcfbb2a5488703f3ea813314f72483369e7f1017c55f463224892215346ab5ce99d0421ebff0e75bb87ba9b4e3b04be03229442e07b04ad07bdd4681055cdbaa75710e619c9a1755ba752adc52b217c8e56ff62bb074f12f150593a21b26210d6c8fc8a4410d3178e886cc2d88c17832efeac1b2996c71c39299b915de6520d8bc50e2f7b9a5c7cb14adb786f2e87db95749340b130ad0f0b3b4545d2fa5aa4c31729d6229602cb8c508a1e93b7b8cfee7be8b2e9866d3374f5baefd0f27843b96a1e0ab7c7781bfd04e6dccf6fa092a0b8f680bcf7cac460f073276b03848c418999034f8050ac4f4293403a4b70be38812e282bcf0793925e3b57e5a1857cbce2bcbfb5563a8a5c6ab871736879087c67edeceeb75cf79eae2448ae833291f1112c4dc76f7e6edc627b3786055c56cb1dd8376705c7073bda9790759bbb70350fff5efab54ed8c64361fbec8c60405350ea6dd4760768fdc2ee6c7bc002e35834d028128659a018a772f7abbd96a0deea9d6526c8ab6bd94b4ad092348591762aeea6cc53a16286964e4b6f8a4266d3362106a4a8288e2713f99a4330a843385aeb62fdfde02b6ea3da7b9fc0db5e8f57f0cac40ec29277131ddd88b0f681335838b2fc93efbb5a980b0bdbe906b2fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h423526617372713cc4152db4079ac752e943687df52c9bc2fa1c0f85430425d22acfac144a6082e8bfbc59b077c24717a2dc4e27de4c14dc6d8fc5eebc08f30012031d45d2fb59c72846de44670ff2098f2c79a552e00dc4c421d0f22ff29ee465545e05de8dd7706c13e81c9467f6ef4b1defb3ae866dceb6e7d7eb486b04ce080f7c410e56709ca4d0678a3c6a4e081dad2a7462f2c487975df31c8339ca3db4c9e82881387cb4867b027bb6b9bace1d098d197762857440da369795ecf639375b471bdb440aa2afc40649aeab26e024300ffffd80c8a58ff7cb17bbe5d19d1f7af91f3d8fecb7d302fd9fd62316c9e48af9e69c83d88879af827d9eec667264b68010ac81b9ce40f149cccf836b58cd2f6ddb789d966f25edfac0c829b92447065257b4bd8af35608a81016e255034e3529bcff0860311884be75f04ecce78e34ad99b15c53151359514696bd79130a85bbe0e125d7866afc13e38a3cfff59347d8e416cfd20068c66423068655ac2327f9b7a8b0c81c4cdef0229a9069bc5a37578968084b05fd7836dcd9590b0fcb66470539cb61f706edaba51bc315665eb10fc496773fba4d92a386158556d059fe1c518293b38dcd0f4c452e77958eec97a097f8c185d55703c8364da5b209f9cb2e1473b029e5b52eb76dfb815333d4668d62e4df85af9087db85443611157133bd1166ea8cd5e749425b3b5056766040e0a88dd8b208997af5a9338adf5103430e5bb94489a5662bc03158ba6dbb52cd6a34df39b69fee5c898dfa6e8d5e39e2412dc77d2e41bfbac45f4e780dde7c94313350bdd05de462f727913992ca502ed762fb7276f3b4419129db0be20aef762ef130dbd663350db5a19221382b885e6db72b663e609461abb19e2d9400fe6b75bdcef765b6bb8fe9a69685d5666fe53dcf7d8120dccfe835d621bde1612eb8c8ccd036a4e406352f84505c3255e9def89a2eac4eefde7ded4d6b8778cd500d437927c7135f9728f6a282addb4a8b4318f62501828dc3f5cefbd8b79bdbc0a05237de7161e8571d904854b56b6f44eb4d76a8a184f635d4ba690b6fb0d4685ae7483f208e09a7c1a63ef627e89a6fe140ab108c6fa822c1fa600c60481846ffc82bb1a65f4b471a04a3103a76342a7008ee766d689108ae449db73bf49ccb23b5b966623ef995218040d46053faf4351b23b46372c7104cd1dfca2e25a0f8cd51153c5f672df682a7b76a1b8c02cd52f6af374a8fecb3506c2612c263a54197db2d9585d1a71fe0344e010c2eaeed09336114976cb29fbb6e39111960d8021c325a642b45eb802daaaae20de2b6d83571e01e36d364db39d9d7cf7468e9530ef7bdd1a2bd4d260d3c14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf6674e3882897685eab1ad676d2f91d8ec1dfd7a59ad2b374117071bdd0aaf2bd07a639ee8a0c637045f32e7858e291e59eddd245aa2450b627afc6370883c718b6fc609eda8e8dbda8beeaab2711db19d23067473056761411f1793d4e03bf5de9ad4e061b29a587fb32eb03f4a9c9756a3718c9b8289e0d933050b718a6fcca203b03fff2e8541d78784c9e9a29f3db91a620c78e401a9d36fbc31ecc159d05f7986de212da783d8a610c84d7621a8c096b4d3f5a10d1c57ff76a2e137ac4f9f281c832cc6d2d714652e96bcecdbbe4ae09ad387453d6eeeb8aa29cfaa5a0f9203c97e2402f7736accf3ae569872bb2e62033231120e32a5a63cdf1069c22c3e599912ed242bc552f7fb42df4f54a5be531e968084603eb9c8eb964dd64432220eed6c40d704377100470ef47ab5247222aff7ad1c0c3d9fc91373a01a89bc045ace8544cb29484a4007ccd163b3fc24686b6bba1b5566ad17076477d815a6353638d1bb8fcfc256a26d439fe1888b916e6d3fa98fbe4d76fb80530f110dd0ddf24c6b5a1e42518f310d7a6d8af5ee9b7359fc1dba7245d1c846dacf642d828ae344723c3274a9d4f3f56a331cef01f1d0b103d9152cefc9cace1f60bac9911e9fa417767f408593247a0fdd2d35cb010043b8540ed0acdd12c005e01f8436f136793c33dd336db246eef4f6071d882573317fb638b4ec1da0bf00270bbd4d0f3a29819e6df76e88a289e2c0f461f48e4596b74a9bfbfa2e1adf011b90903072a30f14c7a75d1e0395de4b35f835ce44e0387e7dfa77d3dcf564ea230833c06033d01f53329fc0024954368a63b228d6428190c488dd08482d6ae8ae657eff3cea6d600396b561e26462f00a14feb1d88d318018d8f94a7c8cb0015ef789cfc4d86a16743bc040766b25d76b4ce7bc359f870846881ec17afddada8eca12846a6b070c00ac16a0e4fdc46ed23ca6d458d820086935eb550d144fbddf08eea9b4ec5729faf3c0d00d634d8bb7a1e23e1a738750dd072d3d21bcdc1616cc3d5154346dfa159a0b55dd4a6ba910d16052550eb69d6a8f5b20e2d1a0ceb72182c1a86f40b5ad4227bbcfcc9834da84beec662d49a0c3efb4f5307bea78b01dbfefec42b71336ea88b344c361cda53398c977b48a4e75e00c7492468cac7f715cde7d035dd829b8e5e13aab36ee5603dbc41fff62633a53eae03f697a48127e908df5ac0b98d704162b190bcb611d93fe1ae4b54408f29c11f33777e48d3792f83fd757340fdfa4d6278ac80da6940aa83f5c0fad51b2fece24196a3161a15cfa48ade9eb0c70fc51932d6ce491dee74c9782abc6a5814a75ea4247b24fe59cddf3945a62edab9ea1883b722128;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h34c9b810f2adaee67e7b11571f0d08975f1042f9893c229e5936557874ada45f404d1996842affeba2e5ed3444065ea6c227bdef1be75696f80de9a81d2670a00cc5f5690bcae78c2fd450f1a66d5aa18bc2fbbb260f5567782de002cd25eb036a541bf9d0133a1e0d1b749cd8a64272c99dd3b94dc593fc1a5da7ea6a10212625ba4973244bd4f1593395c9d4835a6cb780ca250bca8eb19f422fd20af009c83bb2b8374ec007cb0935f1e78b17222d2299eb1a8ec9d305cb9edc0836bac06aed06e394e38161d9a49cf0de0a4030bfab3df57257f4e6917ae3e3c74f3f50e2358797468da39947c6bd8ec79d8262af391667b0a0b7a0fb2c029b38d29b9a938615d007b44f4ad9cdc59b86e3e6b5cd6d25da517d0b5fd96abc295c97956ff0155e01d2a1b9af21e5a3aceb8d7c58c6eac0565c1e3995b393d4dcacd5813b3069316a666e64730e3cd5a724e841bd24004c5c6e5fb1cd9af253e55d780cc71e6a321b0105e0847ab3c32658108d2b365f40449541f40fd3733f1ff7c774213e1b64e5e51779c66383f37bffe4cb3437b4426aee224b90553d9806b2f8a581c476757557aa4c3330b4ede1c8fac1995075ddd60531721325cef0619b9037b58c0247ebdbc6d3dc3594ae65f54243383b7deba776000e8707cd03e9b267a95c106fca63e64ef56f774c49a28394312f994aaa9a7558abe52bf2a61ecea08a5270aab5ab6cae1a695f0422b9cfe65fcc16653b284dcccf532621e67dba0ff82931970570e8f6df827c8f6ac130e44f2c5668f3a5a940535342ec59f2050d5500d2e01d4687c3a31cb9d1f05e6c54bc4c0fe4987c19474eed86a435a22da8ee923ea3a53942d55f4be95e042c0926c39c4ff772bf3f029be66883ce811e400a36a9905d7ebed5c7073f038e3dba63fe7137fda3864a508aa9c884c47fc46f63f75391e3481060fbcd46fa663dd0a6c71907ae916084c77bce8856053b788f3cf5d3229e25d2a0000af1c1b5bf217802f0d03c9be64e4d8d188d2c8cc484ed15a81af221ae4a584ae9ac342ee8ba31012e1c8441688b478706ee555711d152a7be50a7c25aee7769ad3e13593bdf923484105c3a638739f88dce112a984c72fbf63201725bc04f38171b6068644086bf61305929e32edc82c7bb43fdebaf36307b9d837b4a2740860942c048a7bef2b80986545508dd2ff4ac2a84b2c26f8f59986eedbae8d799c8d8d64644a6e9dc42fccf62278a5598294b10fbf0f027e548ba184e336a0507b511858da6e4548dbc3b8e43b03c22434c7fbb4cd894a63d39879884d5a647636064ebfe716a397a7b083b0ab01b8f51c72f45484fc222683db86271c780a3bde0204d27af5917;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf2ad85e47895281399dc3188b4a92d3432762be03a03c5206d75ea64e43e478f13bc9c8c01f3cd0cb656a4df968e22282c3a3225de2fd55c0465283e34fad1a0d0fa24ad4923af5f398ee742d29cdb46b4e4b0ecec28aa2f3fc210d074c8e466990922bb2fbab26d6cfbd435832a12aaf1e829ea23daa663c870dd03fa1bb32581cf0be0db26f9b0fd3c78cf3d1a8273f411546b506904e067acec04c0586097621c9d5e0851e6c24f2e919254843659183c6523791d4956412d86f29acbaaf28df58e8089eeb5b210a49c966c7644aa4e70cce235ddbdbe75155a6acedd2702f2a549a2f543f55b2d01dab46ad2c3df6d066e996981dc31aedac4afc0196cbfcc1214d7420c07d41553cdb069b8a8b857e9c1e4bb653517e58227f6abfb7ee678b6b388612bffe4dbaba4a2b4134e20e18439cad7bcb779e8d201fa836aacaf541a3369604b2c96ebf526259e55793debfb09e180e47b08dac056a3392cf671c1aa69554dbc76c1e078cf1a735975156a2eac28ba801a99865a63c298ef33909f70be4c3b075cd2f01324ee2fc2d19f620c7cbce6f91cfcb0a2f506f8dd9f20fe8629725bef641654ff35917d147e9aa697ca27180467236bfc7693bb6f6870dcd2a5baec03160daaf441100e4fabab865a9848b3ac9894765d22fd2aecba2485318836e866de072210d2eb5f2ffba55b7b663c7212b55b455d9fbfa0dd6323aae0a3302fe75911cc52edce5b558faed29f316c32358e3be22456ae17a61ff14f2bb13c26e95dc4da223cffd7c652e7a9915c370e129738bbbbd5591e2486e9d255ba20e67cbe823b3ffb09a18f9a58ec3dd0aff9f364f5f7028d1bb44a6d305838af2b6d56b852cad92228ba482827773a4ec2901efac675b7d54fda626d311f04a74e319b845fc9e6308e23cfeaf066df91ab131d708e71a8461a07a5ee1d76d7060f1b940c1b1bda8c2e2d94c4a4146088d83662d229fdf02502967ade28d3054199b368dbec5a18d0a589cb965afdca6376e22bc01132f6299d254282efdb63f93b49ef23fb616e69aff3e819a0b38ad745c42e96ff8b2e002f4d12c1f923064dcbe941a3931b1b2e97414a1d4970be08e076c475f8d4ac36c6124f09599a8ed0f19a21acb88695ef21ce2724a81e82647b90fd01b69cd74df9c89909ae2ace71af4feb430ba9bb5c4269307fb7f3e3e274219614ecb2ebf2bad98aa9620a1296c54017b3b071edda23cdf02d0826f36582965548d9ac376543f163ea3fcaa38491b395479406c8a1e2e323efb8debd7c50b5cd243fa4ebf8d7ba8a29c3b41a2119936c8139d322db2368a275ba31fbe007c6367549243dc02b6b67c027ce8cc98c51edf8f6ca53ba37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9b6474bba087b93f75c37015a2cc3d6891df0fe00b52d9255b8941ad6c914eca98d499b36c5895dc663cb6d52feef6517d006b9f706766ba6e7d2b90cdf4de35711c5f9e6a77853be4d8a42ee65368fb941e7253a9461fd90bdbd7e0e316660c0f29f9886ad07b0ec10b5ad67e9b2a04d415d6c5bd59466b1d055664f8c013990c3ed0881c090b47217e61a4c8a2afa9eddf7df413f1cdc3b40e2b139ca5817b99efcd9fea4685da2c132ead7772d20ab2af06ba98d3b6700e2dbc89a2066b9740c7023c296eddac70ba3a6649054b319a14583d3614b7cfe0122073040f0cfc4ef35a8a424573118ee6c506f087152eb73bd4850a4e9e5eb8b46ee52511ecf7d05a1352ac43d86a78b802fa188a62aadd7ac235b362220e908b7c27cb1054a43ead335376d6e5fc49d729f59d932bbb471956548393986a4cad02f7e87ac663e02fffd8ffb347d4826f31f90c0ce2a198ec93afc2e1aed1202c3fd8af299ad0fd1e4bcceb174c987b6bbd42e8dd6c37bbe03d282991e7806658eb242b1f7ef04e9cf9b268ecadc3589affb91339a50139d53a280989da29d013ce3eae7ccae18f3ce58be0316479babb68e6c95a7dd6898c7ed63abb910d6ad518d8c708c9be2aa784766f381a0acd2f666e875c585a11b7147363d6d6f06314b752f9edb455b12767d1974b3907f76d69f216488ebd240baa793b5190e6c2b2703bb7b95df74e81ffc8ec4848760b7b8d1c2e143435859734df7515f5a3896675f513e72dba198fe247a902dd29e6e7a88391d31f46c9e98089e20b8e8847553e024158bc3efbfeeee0a129945429c5b47701439cc875451d4657f8fdc5cdab0322d1d05c0bedc32177498a7d5dee1958ec26367d61bfa847142ae3e1eaedbdd632dca49fbbbbc3ff265c815c7105b300087fbeaf1d98c557b04094449e47feecb99148b7bfba9e5ae905b3e3f36d90cdf9dcea2699aa945c3bf5607e255d1a9c47518354f5d26e97a46a5ad4c000465f399e458772d1cfba8feb34417e4ddaf3679fad56e8e9cfd7e494b719e7ea3349f8bf870ce435b4b5de4d94a9f34d1cc9f46c38ac89835667f90f4ec07d153f74e4c0ef69ca03244025a70d37272817aecf2489cfcd961aef6a94f7685e01bbe68b308618a37fab788ff9d289fc25dc3c76926d93a9914ec3738b91e64c59113edc27fcaac5372692c4067bc44502d666079d85a93c175a4467f7e3834367ffb95ee4cee88bd7e17c4c4d4908ee645e8c81db4665f47c28395f63bd7c8488e56d239014ec97cb9558d7739f7f3a71af3a958efcda2c3158ea8d5fd0bad714da7fdca3494bae5d9c20705778201b0257ad9b3d790f6355a2ce21f29e360ac9d40930;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5402061bd97cce5e64549f4ee29846bd3e57a19bd3f87e2f05cfbcd6e47ab2060fae87fde1ecf96862764bc18a6d0b3f7a23870d9da31db1bd2987b5686f5da552c0b4d89e57692b20d93207a0a1526b1d951b1b660a8427237befa721c34348dbb4c01e6cd54810df90c4b3f76b99ffa11eba4a9e5b0772fa72b351a1453eb000dc95fdf82e8a6a3af89c1a53b3d94ef2652c7a46fa2d2e1b9b0651bcf0fb436d2a1de0e96cb652d8fd897bc596e48a18e174e0ac4f5ebbaae56a88b5fb3c08866adbe407f382fd6aefc95abbc1a0de3fe1fcc57e6b2e7f4b06ec8211d2525b29d4f32f585d78f93344fff63fe6f70fe47dbbdbe7e8db43af40944fcfc0072a56d35775d00deffdd81cbdaf48f702157d7d1f25b68756c326e2e6e2352895eaf8b3823ff11de359895a641f6a5d2f4f20cd4f256fe02f2c013585c486066f29e4438bbcd80c267b20c633603def794f89eab06b7175f7675202ca4165cada97451bfb70199f91e9ec886dd020fca8fc282972b634cca48c39991a98e580a0e6024b182685ae1886a1c7b003bbbdce3809d3dd1c3b0faf1a8c4e2bf3b1f0f4cd72b42c9315a3817e5c903e4f058068d294580e3edd28bd28ec9f02d3e2989dfe56bf7b796a8caf3ede8e03856c232b73808a72a28c03a1e8b60480e87880eb8ea7efc957013067a8d4380e8c39dc77abcb7b60ec651b662b5572bffd80dc38279391fe72c35fea1ba64ad06832a044b207cd147a8560cafb9996f51bcd416375b085b5895b967079b9f0c6eb7e74f079d6a06de7fbf67dc39c387a9dd1f0af91fd0effe090d1f11b4ab2e33dca7d14f78260475b7c602e8ee665af5e89eba8b3c4619b01837891ef0ba72c389404e618b478b1b99dda4b2198163e895f4445981df4e689e89ad183d06f8fe4716f7f00c051f44da3535f706fbdcd6fe43092821b5b387d33ce2e16046de36db3e01bd3b50f7d1f5762dea1552d4b9f84855a80fa7db0b447772b11fff74ba1bf04f62d08ff67b2105ee3c3ab8e6c894c021344feb04314cbce299b6f662c28729b52be786de4a3cd2f9101bdc8c27279e657d8045443334ebb34e6f865e0d00687b24ca569491aeb785477de7a900aa97b19a111e2ef4fadad50e4769479bca0eb4483222f96c9de13643641aa168a2c9ec47b16fb2a5155ed054e9df464d40044aee13d778202940a7cd4d0359bdf7c689554e5a7db15046bf362641a30a84051adf275c2e47a678162108aa52ddf872675b55dbf1d675476ee2e118368a97e0ba563009c35b664700f68f4c00802ad4329fa9449b40b530f107db69dd251f93c2afdf6310c4186759ec249be1ea4dc9b30cb70310a4c4e7f4c891924cda9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6e63451871d85b67942dedaac136457432e5f34b07b990435be643e65b33574c365bbf5ff6e7545c279b106fffb8aa3da146e129c491d0e05a5cf3bcf2771a70c8cf9530ea1f44c49d6b2a91fe5e95f9372f8eeefb3aec5962eb5ca8c27869a3dea349694ecbd243ba9a32a3ff13166a3c5f8ec5443fcd0dbd7972bfb51e2d61496c38f90d34dfdac3f13e46cb56ce911f1f72e7ca5cd2472729f28c890dedeb8c99038794998dbea5a3d80942f893dd22a9872247f232725c4540fc8bddd7bbbc567c72268edd41222af5e00376bb8d0da133983d47a692585e9d0c1dfbdce022385a1d9bc26752062060d2648d9063be4a0776459a2078ddc798e7e75e0db42863b578e16f7760a3be7631d18f70117d690355b0a4324cccd342e3a42352fc52139c63efdde336074d91765ef2748af6187abe50c61f168d240dc045c73a97a894dd58b34a42270e72da8b7533b07dc5612e9826a393da582f1b4b8d5d92ccf8f6a7edf74c154b0d5e7f304348aa7f4465fe791f25efa1c2ef606175d9019ea00dfe07101b8f7732dcf55ebda90954c6606c121b61cfd21fc1fe45fe81db5c64eb7044f0b80ee999e629733e05b5f3871ffc4ab1044456c470f97509c2271fcdb2a94a4a122bb258c2543b00e5ab443e7c5037a36c22e6daaedf2c382ca002a2493f24aad35125735af8075744f2298b9f3c66f8bd7f6a3552820360476ed4fd619cba6141094b0e3b066b5e4110753c1d36f6a00d8a3fd065770d140ec8a5681aacd9a4e045b0c730edcf60ac4d771611dfeea9c4881cca4cc98310bfee4187d931b863c6cc9c84825038ff9f0ab262af1ef2ebd609f720c11b451261448db665b5a5604f9c1352d7b17d0d185133f70a10ec181ae2ddd2dd11467da72682bac09124a1a30e94e237ed0f4f7c86e9bc5b8cd2ae48f2bfc3c264a6d0cffc5e78fd3ba7e72180369020e45a4239b8ea442ee5b69e8bc2de0904af03deaaa99c6028367ba5d2089f826c6f870b39cb087dec130670880dc69435f312a8e7538fc92a8c356607a419ee8647930ad4b07cba442caf4c828bc6663d91e6aafb94df67e79323cc1fe37bb561c9021a60e78f7c2742a8748e0a56cf8cdbc0ceb2e8569b9978c9058054fa9fde2fd0e06df7d33bd6f4c0c56222ce3058be46af5a59e31ef1d5d99bc3a9e9c8bf2c59498873fdb55952494c3f4618f64bb14c5c380031f5ea2e9021a202a24b1263b8a491e4a3c4567815a0f4770f06ba7f042ca57fb9fe1fee2557fe654aca99ad7482b675359b3fe5583bc4f1b79e457c14e24a0eb7a35070a193d4685b302d1e7f3c325e5b61fb429254b918985314fe3c62d4fd06efe423c900baea5d09332b4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hedfaf7d15ba96f030950ddb4a54c2eee43cd6f46ff1251eb843766167ed39018f206c4c57b0c704f14e21207524e6a974ca41ac03e32e499bf069ba5b123014a5aed419cff47ff563e8d90cfa9e1f285d658573937cf82609eb2235717f2da908d813c138e1df33e0b3203461f618ca453bf6423fd2da65b36045b22aa4fefc8afe71d96fa6e7c6a70df1653a592a7816f3b6d296003d107b92d7db139d1bc812209fc32b1aa56c7954830159458284b45afd1af57c0402f98beb1abbb6b7e3e8bdac288ad91c82ed01285943c6f3e6ce52cc8fac82c7a06a2d7305396fb3739690dcdfa9be5a83af2400dbccd7ccf1243b807b5cc76d5c1fafacee8326adaf5dde95ced743439d95c49effe9ea5b509b0d68790df26d4b35574978fd6630898305edc3c8ffb6542738c8d8c67d487f00c0eadfb890db8ec97b8a3bbeedf94a749d0aa8c01b9175138c0b395f1cce9455ef3cad299e86357298ded0297c3dde7cd1698b49a6f00e0d6bd5360ffc288ebbb212dff3b37350137e67c483f0ec5d2538124c3af9e9c335ea0302fa4b3b61bc4377bd9e568dc8a3c7be8df363dd5e678d3260d2db55ec89482e5ca91bd338661867e9b248bb1f4bb5ed6fbcc972de2f1341eff80826903779b3949f2754ec1feb38b079d6536697d3d0f9fbb8431b2d1483b0c27634408e12761f937ce9edc7b5f6e9d78ca32ebc77db4d7798c6af71f629767a37ce236cfc98d3782b65a64f0fcfbebed00595983cc43ce8e31635282c63cf666988eb3bf7f891673365cd8ae4f2c781281f097dab6fa2c438424e38ac0f5a61df15c8bf62a90ee23b6f65a4801fd1ae56c3ee31554501848ddab8ae48b2e2bd044c0b31d7451fae84e3a2a68cb2555aa56e8407a8e65c3fcfd7b9e040d5d64ae537494f41586854ca507961f5d330662702d55ac2a9284d54c79dce9b20791ea55748466ae6e59d0aad16ea045e17a2a4d38da56136f12812c237a81dcb3b0c4b9e98cddb9fe7eda1b7e290b3a5cb07dbc8a22b4fada8cfc845ebe7085ed5094985ddacd37466f8b65f650eecec70f3e79fbdbbbd4bccc63d6fb770f2bb746486b86700a1381caa12af8f896cf40e911b9d94e9436c7942f0d80899778eb92701a0f339f4b9d74dad9a611afd6aac1fe2424025c66da3ee5fc979527a5502736adb7f09d38260837fe2ef7b50ce57b480b03cc5a9193e65aef7a5c929c18903c054d2a6bb000f9640d4c8bf43fab0cb7efdcdef0d901080da5e4af4d01819ba1478a78df12c813627671f7caf1a222c4d06d50db63f48b2d0db85009fc3ea19f1082e2994555fb45e84798d0d179ba18655cd0245eab11eb3ef60969801d496b168d84e87e7a4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h819d6600483bef241d412d1c3417a4669949210131a620875fa82ed8bf65d75aa91baa19964cda43db2fa8c9f662f689dcb76e260770d4f0f015e6d6b14832143d4a435048ea1ba8dacb84ce4902928eb948a23eb0deb99378c13617059b5ed5ca5bb0cb6e5ca1a18f6cba8d376dbd4282d32cf9c0a4c6a56a1e4b2aad942c4c985d7d1438f76c05e904a0451c9646bab6000c826d6364dc544f2850aba0d96c3e4462010d8c748cbc44e9184ed37ff399fdb86426cf7f63404a8fcae83dcf405ae8c57edf621688be9d1bebf12b5055f280bb8d9213f3716a20a677ac792c11cdbc7a6d21ee00887bd60fc7b482dc5ddc66f4f12e070e7c6b02c6293267001b79c02ce0a125e1c32280126ed79eec0a995319713a5cfe9b7900d0f68fa8a4eef48adce9084939ed3df963eac22b1dd78e3e23f3361cbe6a60a62d06f9e94a657aecaeda635977d7e823418c59a8c83c8a1e8702894656b89cda7034eb6680192f83578887127a9cb235a3d6d8dbfd686b4e80ad6af285c3b05586a461c7536722d4892751b95660aa35e44b981a85185765770034739be07778c4ad863480d05ca018d5f093aeb5800e9e1908d326ca6bbf11b3147c4fe0df8121e259b434fa1334d29aa90bf711efd2225611c3e42b054d0fa5608ce78d647f95cfd2fedc54db1c7da282aed6de67dd2c9e6e2befd4fa5130753389a9c596ac8665e0e9fd840eed546b8ab3a4fd6ed73b922b887a5e5d32cb6453c0340aea47b9eefbfbf8c2e6b4aacd3ff02a5f5d499f046ccdb2d2371b750a3bd4c034652aa899c7dbc344d6e4e020ae989cdf8c2cdb7960136cd02a121168ea60f0cb84edcb17cad921768d4914435dd8414c1593b24e677d884ed0f90612c09c77b73810e478f2b72d79caa1662f38fd4b67535a0801981db21ce8f2522b581847c0dae1ca86076bceb6d280f8be0c25b85aec4499297b5a022da110d18cc6890ef7b0b006b9f55763c09516e725265d60221747b72d944fe2c7987de78891a4e385fdf1d6a8dab0a5777adc93d061c3a408dd772137815248ecb6d260a9e1e3d48ba83c1c8df6a11998ecac28ecdda117bd0cb2d1534c76a6ad9abc765a13505a5deabdfd3291dc4e7c1a85efdc0c5001879847a56b4a2178cdafd450c15b04f00410430ed628b1f7c212bed7cc16c2545882fcc74a87853deca0733aefe25f85b83e66a976a69da2d19199941645b46498c78677f7c34e571d497d09100381df01ca6d69a7b8a7bc23a8ae3e519a94bae6a159d5c38b345cf89f509d7d37a68530fb11c1fab38e898803938adc9e8d9df791558d8914df2d7950dd39b4957fad616045903357b2854e2a0f67f4bf5b3a0456f8e8da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h53889b1feb95c53150f4ca9bf9eedbf3e3c784eec0a7b812713e452a185c04bc7ea9618b0b49180cebe8c5572977129a7e5fd032d486e8b4613e4e5bf6f7a8a8371a2b024508f5561cc0c1a649378d3d7eff8417b8da91966c34884a0bdee4274abf3ba0615125d37db6bf3eac057bad0dab4c65df44798f98d99dd638ea73185ca37b8bb96ddbe00ebbd22d69c83ddc4d5edc7ca426a0d22033d68f386746d740fe33fe3f87f10bdc47d927abc1dede2c95be0d81a11ca4b6e6e06c9c9f39454ecfe90ab31fff3c23ec103209b51b02d47fd846149730ce5db038850611d3cced7b15aa53b9abef2596c378e861c54927b6d3a2206ff5667e94db1afd9781c8b19caa1f41c6eba9d37feeadfccc1401865ccde0885e2c5fcee4f68e493bc702ef82e4882bab2c17e81e296cc432baecd475cc75445fac307c92d04580dbbac1477bb678a6ae58b0de80f5f84973a414d33a637f07eb501138143302a0d5871286dc8ed7f9d1957ab235c609d67d6f0b4096426ee8c01a94d183cfb8b0046284298abb96f41b82624f2f0fe302d2e1054feba4d97d230f29457bd96cec4a965dbcbd871e356c160e7a1fdc884a15f79c636e0c9c36e42346db62ea961a5240f28de75868e75dd752e2b868be48f874287b8ccfadb41b58cade27964467eab6684a37fe4777d5792ba672dba3bd94d9a640438969621c326131ae93f3a58d93c6ac856c26c10e8d78cf4a3369453e85f2da5f54195d77c62e67c70c7e4e6ff7b99b740d68724b47520078b2140f6c06b46ec962bc6a22aa997b8d3b46dce405992f2c573311c665455ebbfe653837b70e5a84d838bfe9acf6aa9ac531a477e4bf3f95fdbc2bd87e90c87fcb29c54fe8a09c5a09eb822a2a2b0ae5f876d6dc41d8c656e844efbcbd6992fe1c96af7f22c8811963ea51287d36396c715bb015d7a6a539c24617a2224600950a5a131a0bedf930cf98ee62728e55628602df004c239085c64f8e837749ed2d557c21198b0fdf65f207100614e155375415f1670a37b5d300b77afe1ce4085b123ebe965f31729dbf19415f41c269f655bbea13e4670c811d0e375643b241e17881166c8e0a2868341d332f065aad12a53629f12d487965d49da7033c110695ed1e01b6ff87d8ff5834a744db9d8cdf1b7b3bbd6a008a2cca9531b0d9bba10e99d124c223a9908dcfd78aca1dc8ba6aa38b00121d0d2eb6058a3a6c49bc0d1e21a27e7152f2225ae24791dbaef7c9716b548a4c02c65510ed20a460b41f9f493732d757817f31e7e21ddff366024e2d27a8b5a31dc71b8103bd74c63374dc0d39814188bb9aeab0dbb7630715d985888c55306c999d7934b72e21ffdacb7db2766f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h41bb66b887b06dfa98fc0f97e5b6a37464e85e62fb38cc0e7b31dabc618a9f39f05653e2331a07c81d6864ebee92ec6c608f2855ecbac6031a74961ec973309f6916c9fd5e2fdbab04d7edcc0e7d2d631d5d141b71766781486e0146bbc2537cb546e5a5189bdf9057a63cdde8cbdc282551e86073a422570175039817646d700d62e50d3ae1c6f0dfb3b14a0b13c7a780ad1a7c336608a30b75b34ec9843ec2e9a4939ad626896e9a38a72f87f615b413344c9d60a8cfad561eba41a0c5a70b28d723be1a317b9553520fe73a5097ef9b8fd924e9cb0cc66ef637cf3a94ed0e727d60918f28a8b39910ec5915533df1463c12c0213ffe22ceebdbc4943ee1eff3835f93bef3bc7842cc24194d3aa90659401632d344e3db36e6c1177112208e257c8b545cdbef5c7ac46dc5b9703e8b74eed039d0e6b72d2ca4e9cb849488a0baf2c8b7766907224a9ca844c99b18e1f7b75a2f0548c548d852de4cd4d092b7e47acbb5148e9218f82efcf5e80959abf00e2acec7a58b4c0e0a591a1903b0ad611ddddd725a5299ded8237190bd82a86dce3ba74483aa9a51f005e06c80b3bb5d693dfca8346f7ec4c75dac2a1c38713f97522829a6885a69283ef72b768afb7ec437ef446c966419d4bbed9c10a69fe39bd35ad70b5bc3379aa23f795b4e29fac527425c57ca120e2adb81513bfdaecd830d975790e23ff8907269f25ef452556de1ee594d0eb11a52627d16e0c7e44e919ef910affb3f701ae9550cf0849dd66dd349629c33e719b57bac243751a7833458e8850dc3108dc834c7dc2a47fcce5caac1fe5000a3ec93a9ab1ffe3181bc0523b482ef4bec96fd1f8deb0c39278132be6880a6d31dce9451147bbe04a622add031d5d9cdbbd6109d2c667f3b0f30af4efbb20c78c05343b51cce65e6da34afbf771124bd5d40c9c47bf66b9217a3ce5caf3a98c64c76ef76bcdb5055f19eaa6e263b5f67c7d5dbfeeb60ed3423ed81ea88735ec5d31a16a2d4b31690d7446a115c663950d31bbb5f04e97541aebbbc0129bc1564c806bd581c40aafbdb324c41bcb95439f6abb6c93d92fc7019a74057ba0c346cad964b164e5e47ad7e7b917fcb31a5666b2be86ec01f05125ec07ee82ea8fd9f8f0ae79bdf22402d6ed5b058ee98b29d076d7cbc587157694347a29f589a6208c38786cb0892b3b29ebbd9f2a4bb580be7404d0fc377d5a74820261b6434e8a72898d0da61b9a2632890f69a51c9e6469d7c4235be6e26fad21c313835325c82b7dc3d300455e34c76e22d2c0766ec38ba067d174adf0f0bece00f37c4f80b5373a56d759297147b6269aa0318c289fbc05d82b1c4d266b8ae7c7954768c3ee6434f7ef65e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h2290ae42cd47276a3997a01cac08eb8fd2c1f62c3d1ce1bf6e871488f89c2bc83c30bec6976a7a7e75faf9bbc52b3ca6b8f762d8b2158a965df95807746d786c618272763e7f5b937e1b2ca20be13c8ee12a4495d4a9394fd107a3a2ca003ca097ca39374941a248bc23102873d6aa326736c1ce15552778ee9384395a7adadb3b4df84e7ba6fbdeff3eff145e3b20c16911826ee27cc36168ddd6750d6e226f3fb247cff5d7018a9a7cfdfcebfe9d7b935700a21f45effb5616d1e1107a3b5e2fc18673cda97a5f70e9ebff6453e887fc001e37f2d54bef321428bd852d944bb29cbb874edabc6c2a86893e5ec255174416febeb4537a87f9880fa2b86b78b2010250502ca3e54b6fd8621ce01cfc757d0db6b8a3fcde71d1024aec5f37bf9b8a202593832c800df88cacbcc12fb0857eea3c21d92bc25dde737aebd68d98bf4a62845dca91bba9275ba8fb9b4d736880537093df37bb9d92fc3aaf679cb8831cc28ddd869df1faabce8eee868160052b55000987618136552aed33b9229aa882e1c1481797ced9c9abe882dba6340c6b4587acab1ef149f18fa160e3c50c8a48e3dd3de5d421bc832fc0a946f3e98a278382cbc46540a82ef7083e49492ad479fe9a3e288b02f2939bb56b6bb95ca9e272aedf4a5484cc544a90d40fccfe4adc76b36fd904a170a0efe86015739dd35f611bccd05c00f198b695d92fed8c990233add60b264d347c9031f18bf38b321fc5ea47d42ffc3accbc9dbef8b0d6f066791dde57e711772654f02a6e2f4c6f52ef515ab62a48c34e92482527a56183cbe08b3f6572ce672a53de1f5a75425f2145f61f151af88e376c36670a614cee7cd4534f6040cccdec53476ff5a85e56e02c9cc5821a469c9abff01050795bfe87c88ad24265502056e5dd2e13aa6bcfb64e8e4d88e63d4ab4220ffc4f88700ef1b0722a2489812ca8369205bdd87efbd84a30f1439658fa139db0f34ee619a27c492f60310366a66067a2c392ba93bc6d94e11efe9fcc28f06fc2449c0d0b98d616d5af62a300595a4e51cd630faa413cec4b72e59c35eaacbc7cdf21ab618d079e3e5bd8621797aae7124665ceada113d658d500610974266d532dbd370a02aeea0be5a8f15c7a676fe6b2d2ef113bd01bfa14f3ce42a3b5008a25d3b2258366b9420d7c7b20b806bcfce190eb7e611840b52e6367c06ae58e32a145c5192ce05e4595fcb831bf26756a9f9eba28954b45e36cee6733821ab1e34e50152720f9ff6556976d0bfe46561bb84a76f3d1405645d0a75d0008e376bc31eb86cfa44c9d91a0f604461cffe1c1febf53ae826ae7311e03ee9f9937c56154bff52522cc1c4470e34be4ff06466df6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h339b23019c4688614120569666504d88f6646c6eba1de8995e0451b6e03b90c4be40b7dfbfdf4b500494e9645007d1a9ba933fe6df889d2ba5df15af5f16cc1d6aee30de7144712ff8e83446c701adde58c4b92c7a37cb06feefa337a3040f3aeb2a4f8d411dfbc2ef672002723d19092dae3b9b0fe770ecbe61c6ecc1218d9bd3c0e93040acde7a5860eaee5c528a4f4743a2a872e251a29ceec61a77515748387620897cdd54c9d080eb4e74bb81c9fd9b2d879c6a9313c9523049a5a8d776990805375c770ab9aab7f29078e8dd0d94eb70dd57e5eec996811a1af215ba1edcb461dc4b2f3237d3cdae8d5d5f42b7a2f99f273ef63ba3efaed66b3a2a4c196fa20369a06eb146f0e4e40a943774a67292254435b1a4bca26576919b1d8cd01509a7fbb5c5c351d80057c05a3758d7bf854b6f4ebe7cd82fd6cbb091dafd15da913da72e3e9217b07e964652e849b843a7d2152cc349c25fb65285bf43824ed19283c8bda9c65fc90556476ba1caffe46e4c3fffcd21f223caa0b2427370abe970e3b0478399c60b03399db6db8d382e70ba991067065354c2a8d03348147ed65170eafd5319ab1aa1103ec0714ff328a694c97cff9c730a9d28455131cdb6263b12bc3d0cb28fd89b4c72b7ce1fccd78fac5a0533c3705a726f40a080e57e5fb60a34dc5c93c8b579051b86f06619d2c9574b9a218cf8d68749c73554a0ba075840dedf5d32fb18b840b1f802f94e3679d707a52cf3bd674a6bc3c50c8f7672859a7d08babc3190a22f93d1703489b05492b46e162742f0b6eae5466a26540de9a0fa758a2f82c30b465240bd12abaeed2c04fbd620ac326bf6d8046c9526880297f2592cb9d9f2fbea63ce7c1d7452ed518a544575292b0c25e66e961ce361c3f18d43ad523a368de0766a50e02bd5084fb3299731f886ce6200077f9078c4efdb3a7c4e6157850c85c4fb84300c5e0f9f4838ce59c5ad0e51e55841ee9a6a102dddcc83b26a7ef4f52dca48d6902007b41193931a1c92181eca62f41aaf0e7ae120cf9c22bc34a1a2c444c186403ea8c2bce1604f3f7d253df9f2e7c0d5c76d00661839b3a3d4beb163a232d3020324265a819bd5965ebe22fbf731f6c37a311e162c4f5ebf1c93f1ffdf829474abc2b3edbde3e48780b16dc9f05f1cf0a4b2889ac850ad02fcf157e164ceabb9586e17822aa62df7d20ef5cc86bc97c6cf41f1655fef41d63036a004b10aa3012702f83617138d4525b97ff9a09a07a7e13ec4de80ce90e766fee846022468a598ed002b735007eab489d56e1472ea970ae238bc56e961fed2119b6347df5b863cec75808d98f97eb2b3bfbca33f906176dc228e1272552db1385c92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hae665c80607fc7d56d8f93b58bbdfdfbe72368ca5a5dd7e5c0d4f242bbdde61a170d498a84ba40178ef05f6527af78447dcdc9c2826fc39512eae91621fda7208d20b2fc417f175630c8758590bc45dc4e2a96c9e86e4b25405c05f6608cbddb59a02b1fe44a348f9807d4fb76b9243dc19209fc5bfe68128845c5635dac22f555c6f44696e765ed287cb0012682d23bfcb909d7e1dc918b87344b435e54b24c4dbf4fa2b15f53b4f230c6279d7911bb60d879504d4f65bd1721845fec0e474c4733fcf8a538ec162d4612e29f39d0dcce88d45dabf9155f8b5dba8ea57ebef4374ab1f343177e598fc453b271b896db68907bfb23e4b6c5915db2c66b359669989dbc8e1c928162d152226aacd909dcfcba1e9b9052c1cb3970cfd551f728afbdcf2440a338a7b889b3e00ec0d56ca8fab89d85be0540da14d512f8b95cbb18777fe649abb7f261815fa99cb6a5701ee5dd2a9636c739835c1538c3d1561826423c914416bb5e1f3fa795eef463dacd845b2138ccb1323ea22dc26bde92c12491105396aae3620e0cee544e610a4f64bf7289ca96d33367e028e3ab696c064a1e5cff8119cfe53ba204e2d8c99e3d99483dfa94e958a963701b4cbb71a6e91f25d91fd9afa8247c6ec9c78b8cd215443798fd65d8232eec863d443e6bbfbbfd262a07cbce2f1f4d1f2fbebf1a377a5dfbdc7a073453f5f301516e640c8477a7787a45fc6c2326ba88814ba3766da76877ab895cfd11b683aaeeab3c04eb5563f1dde9d539b5fad083607e11aaa8850e2114a2ba83749ab3301b4bde6834b680454b83ca4bd70eec806ade258479596831d576f71cd43dedc8eebfe5d2d633262349239b354a4aff0401cbbd5d99fdb239135c717a493e979ce88e07a0e7ef8f861f38d21306a06a66d22f2d6832d5909e6fbc7ec744be8ca1c1dd0859b89daba6b1475939165c50eaa73dd71d278c323334b8ec8e6f7ef74c622ed9d14cd754b46d7bf6cd7b6a863f9eb897db52d6d4224b3308f52dc6a7ddd1472acd8b0d6146e17ad2470d9e9fa1c496cc7859f441cdbfc55c84d74bb4d171f3a44873fd9e00f081e3f8901d3f9e51b3fca81787400ffff1120cb6cfd7fefe4f1c8a83bb2fbd98d860617ee9ceaebb96258fd1e407f73c0bed775e4b952cf29ec9da815b4f8081a66cb7213bcd468da22ebfc1113c9b16b472275404040b20cc38633607e0848df6205e589e362532495a3717b1441f1d46019fcc6edecc9d88c31b86b4a95ffad1545bf8085a73b7a1b52ff83827e7cfe7d8360bfc4361d3c3e4a9358a84647f0a1e81e5cce833161128d8f39d08232956b6e79a72c61843b9106771d81c4890d78cd385960abdda91e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h182fa0aa64c19089509830b1d67924ad2aff326cb4d50e845a44a5f16ae5a7d9dbb510a493f54e6b1212b8ac5fd5ac8a9883eed41a8db10bdcc2b6fb953337f7407d941203331af4ec3eee190d78899538c771f1d34c5bca2109ad4ac9519be1de954d7d2358c742eca635dc4bda08ad4dd473324238bc0e321bace6d622e5713457450d75721c812e14476fc876fb702ee044475ec9f058ddad7ccf110424fa49bb60b0160ba4e3ec027615e72e29c04872793a7ba21ecba152de45cdeec00f057a220244aede70bb4b6dc7f37b93e9a9e0f85fc91e87c9139fd70581d03d73f83a60d22b5bc5714303ecd32b456b807049e6ea16e23ecda6440135791ea447037bfc422f712d80ffbef14230d3c13f9e97a1e37b4baad3b81d5b27fa41fcd50b3fd11e5057f1cc698f8ddcdbdfcc8b030bf258cafbe573bd3fbd018d8cb04a0ebb6de736b9e435906b92dbba78f08e6ef161335ee2057211b5b1d4af35e823b289ff3ee6f41bf486126084cbb552ba1deed12ba8cc222d8ceef4b299fed6713308dd486741ba6b6a62e90870fd8fdc84d226e7f3d4360d54f80cd6715a0e70d48f3f710de70740d38efd495cb97db66a9abf8700b442cdf06515b0d2c8575aad17a4d4695c78dbfe6b959474dbeec1cee2fb503dc4da8575c54ec1834337fbd404fcc0c49e0a843568b10123a03b7e0c3d1fc772fb3f30a5c36468c6bc065951d5647f8f6f81b55041c9231a6433e0651e822ac82e7a3840a11fe34e7fd11e2d155e322c689466958efa7336cf7bb2540e86af672f47c85a71cb7cea1ad327d3db6da8ad6421daecd96f36542d87aa3599229fe74e6c53d509f6571e9fbd528c2f4c64b6eb21d69ca25f1ae826c5c9ca60079ce1031f3d2c47c3dc0c5b495e1994612052ca8a032864838ef99dfab2fcc347c7d9c84c035e9ec6932aad8cad6779f02cdaf06572f108a89e6b56297723aa883949d3a8d8987ef49edd4eeb80d6e7174f28edd6555b9bbf5746a04b3d6f52c141c28bb355f07a08579a03ab8be108d2c6ef8f88b46d7ae3ec40b3fcd1effbb1fc63a992915b08976378a3142e592637b31ac470a73769155945c05d2a2ab0737d601485592b6af46d8152fe57e1c80a97f360d2e1376adef4ae555604b6c623f61b07d65f95924a25eaf907e0d06d4d74f778bff8b5ff4d9af6d506b584d66dcd5c114278fc60c42d640b89fd45ba2ff68f0e25b5348b97c28588d6b707544184401ef706f4b624cc6da2fdc7ca503c3ae5c0805948084f9a0961fce0cacb5505e95e5afca069fae4adbeb185dbb2614f947fe7657cc7cc6c317b6110e07787a33ab2440d5fee77ed849a8aafae23f9526b14792025663f96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h456d2121cb76c711b30874e22c7bd5cedab175c45cb97061209e9b2b24b9aba5f22bc1b3dc93fe63baa05bc36bd7b8fb1570719c48fc6a9a18264eaf425f37ec29277bee010e964f714a2a346c1002c47db2ce359a6c4f5bd3e8a60950904bd38b5b11ed322dd32804be312c124872ff894b9be37d3f430938875e2e9589d75cf873ed4c688de15db4a2ee13b1a02741aa151933d6faed67ffe0a757209ae38e4a9eab51640504a645dcd34616c50cfcd05c8b0588986e659bad0e9d6731c14abd354075f17d99724144566b75f103888ba2fe27af4c66bc841873ec4c19c75ef2605e2b1819b4beff883e87409d5a4f5796a20c278357b9743747d37f420c19c4fb9a0423cf11ac75123bdeae4323c93258c9d1dd36f6fb81fe7b1911fc156eb0740b64f553b1ae4c4da3bf584c72864809087caa0794e22b666304aed25868291ed6910ac2a0241fd0d831bff2c4da4f45d59344ef9357ab3106522c40dac2b52aa62bf102a444440f07c14b65da83d59057fd0d91e362b1665334c6cfff7c891e714a8d14a4ccac5530860ad4368befa67d635de50a81e222929b623632b4648d4a2dcf563fd45d76fca1adb7c5ef83b6e96260d9e9066e09c0faa130bef922759133f12224bf8973b642455dc96768d528e16d1f9f4a96bb1eaff21e5ee9a44803943ee6798fd32e3862ecfeeb954f5a3741c8b333d6f45ddde893c14c062252db4e4b9baefcb630dc7b73b095b0f24ee00f861ca2396c0151002591d86a0fa82eb33eb17b7b7d71f47b19d5321eb9bb7956312968507484d5fe24db50db37976110cced0b7bab4d458a7e3ad2ac73040b18f5083bbd05cdf0ab215d24a81b7c812e60c61ac7baa9570b8fa656d87884b222a6fc5846abdf55a8bb659ee54a30430edfca2b05c75401964c17b34edb1fcf0cdceb669bf240bd8d6b5dea1263d32c29fc4681e2e69d72c8f9f57a116d78df8bb1ac702c75c86e4f46656ad562553492999aefa3b7f840e59137498bcffec47d45242e8b18bd596d1b364c997eb7de2db5a91212054233bba0dbb005cb5bc6b5df582b5cba5414c98b808307c625329628c82e74799136e1d3c33df60a533ec1d51d7eb6b8969220066be0f2b4f128b71818cc2c5c4fe8869a2cf1519c13d0c45ecb660be98780c13ccf80e3335e402b84ae1d3deacc31d0d2ed57483ee1cb45d7b22f8e4b222a11072cf68fffad0a6657f287be41f4484a432c8cf068410c138b8a39b6c66be147ea93fdd274858d7a063eff1f24a43f604894bc3344d866aba1cf874d77f9fc0a32fe710523e3f2417047cbaaeb879acf25a5761f79aa3a61b442277e5d9232fc9213f1ffb4eb1d17a9e59efa7168dd07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd4acdb67f44908cbfe8cab84d39bd5754823f7ca7eefde3b1132792e28b55502dcf24c9ecdb830f356c539f5be467de9d9c4470eedcbe06ea62b2e50e45f7fdbef36dcd294574d0fdfcca69523bdabd0deec009ace86358278894d71afd40fde4d105ae09e39dcd6300230bd85bff0ffc43af8c3dd8526db73d057eae8fd666fe0ffd9f6d80f30449a422bdb68bca6d88ac0718ac564a66282c761bc22b0c4fa9cc22fd2ae19fbc2910029d1501b610186d58f9dbebbcfe3f5954774809aab9810caed73b88b6f9be9f1174e22355b36c8a512cacc94678754f407cbd130152b432940d907daf9532592f6543047c4d678b11024917b55864b75b21790c33750379eec36451e84e8e71b42d47ee6c390d2807f13b32dd256f5653b548df6a3d6a389b36bcbb21a6cd84691419828c562d7979dfaeea3b92bb33fc1102e8106b95e0b9e14ecc6a392a63a4df100d14aabe548475f5ba4579f3bb0d2e7f6836f93c34e6e48b130a2c09cfc5620d8ad302675671a2a24dcfa9fd18c6588257eeb8e7dc473e9548dae133ff7c160d9b036b2153b5aa22995b326a8ce2916fa276627e82269d4feb79e6e4e78a27f532716b1b585e473495525a6beb8e3e0349ca569429a0780966f4e65f21d1b829b87d33afbab37c983f1c311d831f5efdd8a95cd1dbc3b054a0699b6dbd7bfcd2b6e4d03b489d43639f08098baadaff3fb8698a82a73e329827f2cd5d6292ab771dc1e1469055829dc93869562cb71cb5feaa64612217591b4ddace8aeb5db56817a5764cb62730100a1b9ac66068dfcc257a368ca68d6a89623e9a4bb37b849b546cec448f6ad96514d2124caa82c99284f41ab7315ca5bb6cf6c66a1f074e83a9307d6ac059cbe7cdf9ef31dfd2f460fdbe3c56db6bf8537bac82597f535580ea9dafb2a0b4d758c57fcaa10917185dd358137b2e8342b704ac2441dd46bbaed874de21f23ca663a99018783743b3e16551de20d21ac806c5c461137f51755aa79404c228ba0caccc7a5763c1aa474a8ac0243b557723e2a0f15c773179ac67e55e132594ecd8dbf41d9ecbed61a0355d810885bd10f0a0790b3ac57f87b6c49a4446ac4a3965675785fcc9df550f0139ecba00d665a70b5244bcc6ef0f3abe58784231827e16cc0ff0188a5a8c208af1bcc92fb1b05e921ce876f8d1924bfb502eada3872c7a45dfc6077ce87839e366bcab851715d01dc3e73299f440715f19de3a27ba3a05cefe738abace460b1fb9813408b1a953b716f272d0ff744513a6e64b13ae4d626b4a05176f45c0c03ac22e7a1fd423a7b9cecdc717b145ce59091c20c98cacc9542c0b8e52f5c702bb7f6e50d9d2284c0578fadbddbdfd4a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb3579f5f583a8d0b7bd1e1b83bde0809fd30d9182068dcb0ad84760c82979652e55d244df04f8f155186a6ec11611ca3e2db6538f0d4b8a19e4dedcc9ad2e56f711ac0df972197030bb2cabea422d2b7aa907e5d7c26fbcc75b4a109ba738df5f61136b62bf35ec836770ed328a3e49e708dbe022b063a5e42b64f98a727742d21a755940d6d83976360a9c5b4d058d0fa7fcd58876e0ccbf690650bad23dd99930409448dd546454140309d6d06ef4ef666265bb68cbbf35af0d1ecfacad2629923e3e74059a3331d1397618a9e875eb0800e2130beac93b73e4ce463ab0cf89fc320b1acb93de23f72cf33a29bff94ec683ad7aad9158c423cacd8a8a69c56aacc1001ac5603fcd85e0b2fcb8e20b06513be2eac28c605c00010c7af71fb8fe1c9ce6e6fc4055ca1f150aaed99269eaa6d2170ee289d815ced958a47768adb19a397813351fdc63dea8afe16b4f6347f58a47d3747bc64644aba1caa8ca0508d170aab8ab012fbebb8256f411cf635ee48958391276748cdd18818ffb6fb28dd4f9e910cf96882b7a75aeaac3da4c6dc9f58d4c54e1f9a8d0c2267f545ec83843065f9bf175c5f9fddfe73f2c2db6ecd4d333c37846710b3bb2d76449a3affc6dd42340b039e7ce7ca3d3d22e760b5c13d188c2a82c5cab4ac0c5d9d1150eb1220f1fded1b51638088aa301c9c51f55b8783ddeb49e3f233ef6bf215ce959c9689f0cfde310d629f6536644a2de473e3bcb9b3cb171cf7e2eef5bd50fb938d32d02b03ab89aa8a24abac9bd259c9f1a12ebb95c5d7553614f0d8566c91f9825180e2c908f122737fcb984bf35487187019d668fed6d7ab3f45d811096f01d18fcffb7b2b886fc85ff353fffce5f710531a379f5d3e5e3735636e975017cee874e01e77c9880b820c7077bd912b2c24ef1b9c7a450e9b627e76f189914b00a99675b9b0ab636d6c400757cac0150a072574c85ccfeb9b1700d0390d0f6659ad247c2f62e297a83051e1e66d402c4c4c75b0df69e62a61f4113c7377974dbf53c617bdda2b9a751eeffa06d6a9cf99ea49ba4ec3cfe883194a241e042087f29fa47cd7ce1bbc4cd88d23083e40a2fd71e3b488ae8aa103550a703e2908632e89cadf8ce993ba30f2b00521e1b0f9c6e8696f3a6038c1ae3d62772f91ad717a17fddb11697ec7d934ba3446ed5089b666f0e61be17cea4fdce1772fbd4f3ee47f3a398b3a2b46caa2018e501317a358c009b2b043051a2635dcf7fda7e93537078cd95c199da6f9afe266967c95d7cb1bb08b2f7bf095c5052bb307c082d8a3a669c1508f193c4704f00fa985f6c8ffd0ed36754f62d78fc358313e4e58c6178c2b44ff140172fdbada7148d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdf7d97e2b0bd5442b54d663946007b3b1bbdc8b0ed4b275db18562430fc4fecd75fd4db0bff951434d23ad848e979bc20f666b61b4459030b9e8bcbc0408ca05e5ccac9ba6eb2268ef653f60020a28b7cb142d8200da23a83482b1ac4bbddf50798a81dc4a6ed06d558ffe19884f13c0ae377e38656b106b44cb70d21399bc5a43cc955b84175ef679ff44b4d4009b0cfcf5fe532056bf3ef8951a3345bf23f6a78022953c8488038d8c991fb498a205b9d580d21d92001c4bc67ae4af21ed07340bade5c287251843d83094ae403095978c16c5f803cb892f9b9d580ab69d0c2d61c9033af97b5111291db3f6fb3ad96a69b97b055f7f6cf92fee447d999c5ddde6ca04b36e0e414dba1009bdae8b23e2dfb17bee904f3f9b0cbc6b86fcbed3237b454f6550fefe8880fe1a16e4935ddc8d279cb1f8a46eccbc44b288fd51e34d10c9de6febea406ccaedac3073343b647890d1e1c89b44ec2964ede7a3b212a2d56b9382a70ccfb0819df06161812a6376c345297dcf313342b7e64e72458331cf3779a2e35c5ad22d3f510546e3bf2357ddb90e2edc8e79cb72b8a6bcf24018433b3c50511532365f0dd33eb3251edd1453d44335167c97db505631efb6a2e26147de7d42d8c2fb2fd7c484031d53c1ebed306ab8f3e6eff80bd891ab05eb3c11502b49b3e0597ae85878cd907d46a10b88e53f1c8c8dfc199d9c2254b8353502af729e1b9880eaf940a74e2c37de76981d52b7bb7317d725532061754ed1257c70a89ed129991cb992d5c269327af953b7f2e42ddf5ec6f61d8971f423f4724d8269841e8a7ad703ed83739aa43843088aa2470230f18976825f9f7720f759ae6d28df37699918f93b806433b0eea775db9770f4fc31434f2cc501097e20ae6f568113502a140a08812f27f6d5b97ee2d54026d7beef8b40fd3c1e7c0baffc48bc97951f04c500ccbce6263625fe5fb978de0c4e7ac1839fd41ffd18ae73d11de2a98c88eef57c7ad9edec5366191b6bd1fcaf47fd0322dd0bb0d89c9dac45310a5b7c1cdb8337b8c5ca19c056007f565e99bea80e2674dc87c001219b77e7aaeda35bde4bf272e58285b0efde3701d93245e314974560fac9b762b2afcd3dd241743694f2db19f1e5adb43feeb3edc77ad6a86a3dba980ca056faab973457260a121d37ea8305ded74b5fdd5b7926384fcf550bdd56544768d777e3914bd134d50f29d3ce0986a475cc02085004616e0ca786ae8a6e1d496a6cc9824f29e6861e0806037511d10fe272ba0c744367e8132368701af50cd114620eedb4c698e521e8a62d12c2d4963772ed4e3540443d3487cced17f5c115eedf064e62bc6a9e5055a8241fcf85785aae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdf30e252800d000d386da1ed0a1e17197dc22638b2f1f51b64a24e959a1f39af03ac99510c0cf1352b9ed3313e54c2be71756000d915f5b450062b74657c0c96699357f559efcb3e2cf32b6f2098ab1886912a56f173aace5fc6e5fd9f4d1a9d61ef5360fe542648f0bd84f6faac40e0e37260fb618f29d14404427a155c9bd1640bd093d18830ce206752207a4b51bd7d1dc4609813e2f786759144044e305fc0f9e3bf046ebe75ce3e264b8d40840674563b4028bdd2fe5d659ffa928d52fb13d5b300390d5d9fd2967959b73324333330ea0489f576a5b8ebc0351cc634a1043b3845b357427d843960988a8e470f66701204b8708511d4be70c1c8352cf1e70162589d90d7106a9727c26dd6098b4f3ba4f8070c4f49df94f6cbe6ca1b238d00ce026c43ff8d48959187acdb7f6776621e8d6e6b64339b8f33495acfcb6abb67c07b84ba91a0b43586cc2b3f2e705257148cf2db009b0cb93bbdd1bbb594bf531c059a368d89001deaf5dfa0bcd9c9c61e8e84db46105963df816a1a5cf16081a2c416af9cba16dde108a515e545e43c753dfe6779201f5594f60b0575cf4e2535c1aad16f096a719e19d222e3abfc992270636de796dfb78112a73ea34aed5a61f7172a47fbb89589ab6b2c467a991918df8c6b4edeef051a1513cacae5fad6b45db44bb8d280d5a577aebe4ef91b7a8f325d9ceb527e9296ca952fc1e959b53ee0f36ebefad838cdbad7fec5da318067e154a893b0fd353064d34174a5db0e16f7d3ed1245a0e18fc99b9c4755b14c3d1e25fbdcf61ec4e1fd98013e1bcf288a0cf3f9f91bbf2330afe5a8627faadc7e1403b3d23d5a91dfb4ff2e5324e10f136f1ff7ea9d23440d0eb76cd013822ba905ec56bc1e3b4b679e9ec904ce6dcfe615325c523457716964c54c1899cca87e5d6464430acf5954187adbf87a9c80513a10ffe73b26b8198aa3ec6cae98bdd3be8be620efa1f75ab60cd982094c7e6aafba08d323a2a569016301916bef1406435e4b21d31c54217394e628532b5f8fc840dcca6d8dcc5fc1b756029cc5a1d1c3a0b90811e1caa8681a436b0de0217ee1ab26883338e355ebc57ea6b47dc3e2a3866e6a7218892632cf169a3e8c629d29624954b5019c21b26736f4fb50a6f37f5224c8c2cc9c027fc0f7c972c3cd6eb287111f32adf5360e69fbf4cbe9488d90bfb47d704de0792464085c4781a66e3f83c31b7332ce1413e947f0850a141127b8c7d60a46cf977f1d8c0d592a8377374639195ae51ce772630b4b7cbce67bc3a2e3dfdbb83b0fcb984b11c45a2601cc0aa6a182fcd7cb01f91adc520240b45870bd0bf8a833aad712ebf4801530667253a1214267be1f86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf1fe6e3de0aaae7d8838f0b2628c64922c2fb1f821151a1de3befcda1d0046204a0b201e51aa10a1a3c574de2dcfaf3ba40ddcef556e942af2a74d3fa42b5b97e51de1b064b5cc9ea2235676f798898e3eb4d6f9f34c1fd0ce544b41b8617b603ce3954413c1bc9f23aa0c75ad41ea0f9705fde3c63716064889ad77405020a17398fd2b6b593c99e7cdaab5ccb594d3a02900a6c971c423e3edbe9c0b13128eed35addd750dd9533cc8c9df3ec217922ce80afeee5f6f313a85fe227f94f912283aa5f191ebed92039e9f97618225b7e34c659dad547e709524fe1a2b3bada17841756404b66fb466fe58ace5f35019823f25d9ba6e804482440c0eba040bb8ee14df41fdfff2ce93c410fe3f3eff125e40549598e9e1666c0389d42a33c788d5b9b1a75dac64c40ecee6ce1ae3abecb091f02f3ed9d833301b34285c2ee4f9085d7e49960415b22ad455fcaed6708c65e09a97bd3fa84e5a7e66f9286e1cff458acee1b65aa4416fa03fb3ea6a43c9603c657c80313df606a56da53614a341c39b6a1ce17484b2bdf9d520f950ebc6e6394ce94148115f40a6361c79a7a2a01791bbb034c10b9ead4ab7fa6269d21cbad95990c74b77206ed96f4dc1078e50ed4f1a97935b785fe4fa95e42b9371c87e95807ebc98423b725b84362de691b6acd0c1e9ed7330d9c756eac936749147c77651d26dde9c15ca49e50540e551c3d0e4c27e5b1e73bf74af77ff67945c31f133fbde169f7d5090c9e989ab5c4f3e53ffdf7a2baa46533de99e5f5df48e2cc8661917dd8234b2b78521c09733c82f1e18dd18ab463891f4411907df9314198681eb43cc69d2dab37bca4ac12540f86b812db158cf8a8e16d7dbb689ba00acca74e3a765848aad5ffbb66d59a66216d04797659ca13da30dc1381631f20c1242af068de2507828e6faf25d9cb004dd36372d1f9ccacda2f62e2c9fc4510085c1b34252362adf8354ea46a0016ae1919d8350d7d0a2f7fa920fdca7c6dd3d31fe28b4309fec5cbb31c53fc8457319775a41b3cffcc62719b421043e746271699dbe5bf7c7dcdcd00582c0209cb1bf59124b664600d2def70d62436de5dcf2494f0828efb40d36638f22c1a454f82dffdaad6fb958f5fbb27099af507c266f4d210a0398a5dd3a7de279af74bdb63487676cce41dd0b50b5db4b7e51724f1f197f223f57179559af9ba05db0f4dac2c7f2476564f04a418429acedaa10428e6a474e4c1e6e9df713e6f9e04da05ab9aad4f32e89cc6a8ffb77f964d6aba62f038088e7d7f08183628cb9f003aff740062a6106ab94e7cd4d01caf7e0cfe18dbf7dd88d821463768909e10107f9ba4720dd720baa26f8aaadea3c940;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'haace9379b8a4e3cbab86ea51688db174ca71e8cce2d774bedcf6878a331c39456d9378c800afb08d06cb090b71f7413aa4948b01ce31767a16f2d6e7a548d7a6919bb3c97899ede5132859b06582a0c349d1239117815ce7d8ffd6f239eb4914d6fa43c14124cf0743d4464abdc55ea055cfb3ea5cdc3e17d6331f3aebae85260162e2a89d4332ef6aeb98eb3550967b8d17e0e051b3b7ecb76deda6d1825baa5003831750e5457491f7fb8abfbc7cec846b1772998742febf5ed884d02a4dbe13fc2045613ce39630814aa05fa5bfffc86b767bf404a4f96b3b1afdaf8ae7f588dd8e54f858bb8cbc2cf5ff7f52f1328e1527b8dee49e52e0ffc6d9ad02c4c5145f727221567302b7681d8d37ca9929bf8bfe1bc4d269ec5ab307e4305fd648b323f958917b1ce10d64cc8fb0f0f39c0236157c415420e802c553af8558f6b18b6b366e89b739e71ad4bf4efc745146439f2c783f979dae4478c25204f7838bb31d5a11c6d26ef6bb34ca28173907d81ca1709d0665cf4f81eb22c44f0b3966828623d82b20b9f79a9560e056b58ca4a86ae0185d72ec7939ece8c75de46a29b8a65d0fef12938c30d539e96225cdc9a7011a44e5973a5a712dedd611cf280d512f18de0ff11932892969026a7dc9848c1527fccab9fc968a98a4c2fd74f2d2a00001369b6f5bcb2fe3b33504bd68736f082f63825f912c20033527f904d0efe06560529ea14675503bd79e7d08076bd225ae296a1592a022a78ef089a182651e7bf836206834c7a46d8ced2e44fa80e913879130276ce41120991fe81709a7c38b4ab876d4db683bd07fc0aabc85f7b4b4df3a9b727de7ecb42c8f1473d07c201321bfb830066edb671a106476ba1144194d1ffa17a26e84e14a94b8f270c6e8750ec0ee93f7431d958fb6399a56ff292a647a73fb814c1d46c4b7bc5e2d1de6cc94aea55df9275a6bdc8e8ed511d77cfca58b8463f6d8832874b302701a9a616e35e0f4953fb975f2f331ea456b147775e784e45eeb0635b66bf1f117942a04283b08b2698e1fd64e18fb4a9590c68188e017ea85b4c85ece52f033816be301fdc1bba23ee04490c40039db24561db4d97f86eb0e49feafebcf1b284a3054f43a49b181cc95b5c194e2b344a8187d58627771e635f86bc4445e4bfa63944a4815f62457e9e0a6d7a1d4153ac0b6be02d1e3901fce0799448f986dda6ea6ba009eb904edf31eae7ec230b690315eb8b16f4fb2c7936cc26eac8ea817824dfe10a85d76ae4456fe6d2fcbeff5e9601f3228da7dde8e74ff78196e11b5b4ddfeb9afb271449a47860155fc7f174219daafc8de8934806c0b65457f763aa0c31af6e198d0a6a363b4c2f4e874;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdb4ef595aa72196995e70a90cf146727bf55bec8f61245a9d520e6cb5a3abcda4445e414f7c68f4a6c698e1a7eefb181dd6f57aaf14e76b3f367cba1c7f762493fead58224afb0364433cc4e40e068ddff732dc3e0bed62a317430372c78c5e424db702a04f5868c02e1c2dce1440f4c78ab4d032672df831bb2b9bfc96f7809c3d435f476a317cd6e8a82d063308fdd2cf477b8f053c811a948bcfac6e048f69e028cdbd287c84b24bc703ebd4194d07e412818ff1f81f4dfb19b49b8311c9c429afeb864049a1a6f5f5a80df436a5f9c0527210b44c6ee682f61966cb1e34f0cfb31552446134e1623f29ebb8185cf8e0f78682f0392563148e32909674bf50bd810a34a792b40971ea06b71d2d7980d624591b7dd2b257324da2c843ccdf8d508cab48dc37ebdeb1e54e3ff07dbe02aa9292c75f4e053cfe8adda12093cdd02b1cc5f39f96b98af957f8b3160043d62fe93e9c6ca2aac67d0d0ba2d573384512be264478f4b8dc8fd881e46153b39fbd954cac5192ca37c22a0e6d68183652567a0d95d9407f2f8d5ad2f03e99ec9a967cf83e235bb04254b4c59a0cdf8722474ba49fe094a794ebe999d25d223b4910c48bf229fc48046d3e8900150b6bfc9dafaba90a9c20de8b68d89ac6ab1be1d128dc67d9d31f899cb5538270d6257d92cee707e6495d9545cf294d1ce4a639329091717ef4231f2e330a384485bf1e48d5837a4f00f6a5d57728341fd6cf870fc67066319492c5c5cbd6c7f3fe7cf389637a9e0d84141c7c8efdea3a28c9fddedb162da24176fa3b98a2e83022e7de73198d46fb62c63b9ac608c14ddb514fd51e6ff86cc73e73e00168cd9b73cca6eb200a99ebb99087e689562e33c25f4f0f957d869976b0f237f11fde76109b4dbab9aafd09e5797007dffa2cace281d350076a3e813cc88167028da4027d9e376a16e034e38301604e78224b54538bcc4e09bddc77acbe1e6264dcf7afacdfbaea2ff942e8135658ce396a515e4f47c8f7dd92e3f2cacdde9e886d585c07d34d52c236bf07277e1d410bc8178b16b79d24cd9e7d3af26fd24938da57c599095e8ed136d9f8e1bc7f75f043a0f4d96d49df74dcf204dc6b662e319a7645a4de8ea5c573be9fca456e5855ecb034eef924191d13834d55c576e655997d63f27175f5d8238092351a763188605f5030eb9564221a21f4e81d1ca7f845e34d9d1b259568b0ef288c724d38fe2d23e9b67173b05ad6fa9a2e246efbd5eed497d726a5bd496373fde0a68650b273644fc8fcef10ed59b4f01a7bbd21992b07a8b7f74e2664f1ef037382e47770cfd7da608935464bf2bd6712ec7ec2cbcc6819ad973d026203019bfff4faca3f040;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdd9ab0662a3e186f29e3c90cd7e4cee12c5d563ecfc75147a278f011df92e6d9bd3b1305bc4a4b14e48338dfbfb1eeaae3fa885999eeb28d4e01765c25f25047e79a6e148d36ed5f4bbff8e23df6a6b07b118fe90f5f1886ec4440c093e4fee5e632556ccacd9dd171cb8433c672a17c5a0b45fd68f3949cd7fa080e860dce88b187ab190f2c3f3481aab806ecb90666685d360ab3859bed980f53e6d373cb833e03cdf93b822de1121df231022c51c019c00da63ca8402693f1bfab315b7002f61f9a223215c14cdb0939ecf027ebcf3395b74c0c82f796ca2339f96defdfb219ff793961f522c472d541b30a41bccc2d6960f97009aed28c8a1c86a643ba4cfddf0144b57af4df41b3b8147c4fd7e6144029f457bc5d3bad80a365e95322e4a8c1e6f3494e2f211610653c1ce65d91fc8ac98a1bc130c086bb75c482738f8977e83406a1650e5d5a74c92a95bcf6c0f2ed670d5ffa6dca1b58325edf9d0e0aa3bd30de9dd47464c13dffbc649f63185467f383bfe87ac7e226b109d73ee36d018f44b5a317fbf2e3838b1f6245ba6aa8032ce0507699361d5591571a3b5513154137d8a7ec802838de211e769ddba2de649499fe753dd08ce5e857a5f706b375b64a3ccb888b45da775ece08188420a569eacaed60e0ec872704b57aa17d4bf9a9adc2440b0f3300bdcf80592e2814fa3a17997eeef1b33457cb3471c736cb47369db6a3a796a07afcc3037b5608d7b2faaa326c2fd2d82e0497a7ca5b32d0d8f4364b23a1121bc9f751f08a83c817552b91a7b7fae59711ac4d65d53dbdbf5137f34fca4e9d04010d6931b420c2106d1f5a39827497ef943d32004d3436485c843c73a6ae77fee6b130e8f390936e9bcc25950a7fee4d4b5e836cdef7b7d943f3fc910832883e81112bc6c719c03c9ca106acf1ee16786c1921cf51fe6c2cf34e5ec29f0ce97a6ef794c856273b6bbea0a85fde9327ed99cb39f3925f456a47cdaf503f07e5bb6377e1bd4c36bdc8e72cc9e8c336f14144f63494d6c4aa7c688fe2a0f1f0e4e7f0fe7f288c4e61f4fb04de169f16a18b189fe01f437478e8574fea43ce825f25bc2219992a56d5204a0a2a3826c6b11a281f391a6601747cdd2f8a78538deef48aa8ffae4f2580f29a6e6d03aec3db118192c5001b66e54000391ba548e476d31238c0c306c60c9b364dbb0998acbf7197cde969daebf519d6b2f715134e9c3819f650fcec10c5cbb8eb704bb24072708c8db94d6afbf7d70a5d511b06257aa46633286faaec89b4651e493a7bf8d6a4a6877dc2d65b7477b4561140f8da4f8ffe75d5cbce572bc635ce1591bb6b8c4272d37d216d157d07e04625659be9d732584ff930;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h46efa68d2ad75d5e1e21a972da523350a90c914d6df70b755be27a6bb961c3ce4b956c600365344d8ab19a7f34175db1ef9501db18976b0d45b14ed3f688331287ec6be70950e9963ab8ea9d625e77d6c32ca98e5bd552e64fd49176c10d2cdd03b485af9355fffc853ecdd89daa940be3b20834669f1978d8f9adc7f07a1ee1ea23ffc675babb89e98954f53b79401df1ea93489e6afa851e9a99618c8e73514638d370a6d6224bf439c90760a0caae67a990c8cda3812f1e089d29ad454136cffee3d61819826e0ba246a9e43671aa5e7b3075e7443e7659972de2dac681544a156adbfe323cde8051c14e8e191086b4fbd73675425a16389daf39555d6b4f9e934c0fc4851c1b6b466505bd3c2e7dedbd3e00a868241dc52fe08547df6f48aedb977a668720990c9dc9a9e084efcf876c5a3b2613a1f716d121ac96aa046713bb8d39521dc590e575fc9f474fabbad22b912e890c63b9ef01cbcaa106524542e095524c7baf3cc8d39d005f8d2028f29e3537618bee2685aa24ee25d28385a5449666c7bdb75960394192cd4d2a742b0c7b5884b1230332035a90134722ffe4ff191837a5e6cd952e178391418b5ecfbd3670da4529274df858324cf603ac43076608ad81969eed29bbf17ca22c05fc2432fa4ff41882f56794e85896083b729c4510c8225892960e86621a4334d48fa172de2168294de66992f643b87cf49063ca8e0be04152b70359241e0e5bbf03a3a9b0cfd1f69b481622df8e2ff521efe061fa655588b812674638b65b5ae2e3e5dd492e076fee293df6111996352c2583d2c4262c2d628d71f99c2f6f0b19737d4db88499dca8ae5c3ba29c2009159e5abbd837d65bfee197951931bc608bcf3988a356a1af985aed2237735303d30e178fb7798263128f5abcbd88db32d4b202805307947b235f0c86fc022447fcdfc9894d210c59066e9649c5be92355ab61561c4766adc0e808451d146bfadffb041279031a254b94c6a540dc7c8e2d46a46e6cddf2b4dcff5bc86f3aa73d777461bbb4c49f926d78b142c2bf55f8b64d045fd89bfa00f452db2f66033ef1347d1bc8336c37ac0bb94abe3fc16ed11344f9051fa83588b570b8dbc4eda7d7804d9152d0348e21c21d21aebbff3f6d3353670f329684452735f647081764bbc81cb1cf636c480ab31770fb0ddfed95779a0b29d312f88434beb7a13181440d9e36c23cc544e09833abf0cecc25c2b7780900d3c879cc93ae91ddf9e780183c5e9cc3c5ddb9e1fa21085197bf9db55a8aa0d272964759527ad7f857c3342b711119335d389bf1eff6ec03ae9b1e02499dbdfd997ee7904099c9e2d9cc5fa83f44f126dcda6f3558a0931149a3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h61d6cded8ed05343e9638b682e4533d7b292cef885251d8486cf6935fa0ccd10deb47b505c1ee13d16befaaaee2cc8c2da288e2b715c9b62eb1202f56eb4a408b7c26d70b07c0f49670f5442faed90aadfc80573673c2fbb4691160ca41e94c0b72ccc26d250502e7c0db747bf4372424c401290e363266d442d9cabdd003092a22efb9bf3cf63a7fb5f6b40cbebb97adfb7f75d20398f70819b0958269b44a5840005696a10485763b7ff30903f6c28d1a51463b1db99365d1ac3166abd0e8b7413215de829d68c5d14d92ff03316d09a3085b58f35e954d900b9f8486173c35fac8b8a2d8e871c36bbe41bb284c7a0031cf0db1e52be6bd702d3129e0d94af7a6abf038d9741156bb0464f055abfdc9b471e62dc7d847156223776abef3ace177652fdc2fc58bd08200bafacfb4c4b3eb072b9a1892da7ece5b11b98a290b2b6672fd9b4562ba286e85835ca9ab33b73f0a62042d953e852fdd881f29dec972c972e279bd452ff1c96eacb0f6409668f8bc44b17f1be2bd399ec3866c57a117fa013dc63906f102d5b7b94dc381267c22de742fca17b349d2593ff9242f45906d4d8108c44f541f08708e73689e88e5480cf678e57cf6f68807d97ecfbf10ef1af71228ed3314d203f9bef28f97aa39b60aa9c6207f2d80b01803b4a801b79f7d6c046e363618e293f2952b0be6c1201176b919cfe539ca7a58f91ae8c0b87fdb50acead6bf15c437dfb6320d98e384a4faf0a80ded44a1215552b40b994e4142165d807de4cdd9afe02ea7a299602f22abf679f5b142091a2b90d06556f89e88bacb9982af79ebd68b7b220bf1f9f5b2d27d06e5c93a227500a4e604670030502bf63fff09e3a922c46bf582b5ef04ce80c4f64c05b46c4eea550b35f05e240cccc7d6c814894a7eb42cc6846ed160c5dc724e2d8c82475f20d5499b88850eb93a8ae0838be3cd180cb20a1ca5b3af8334a77d4c8b235ef75bdcb9b64eccacfa6e551eb8950bd6f10d15f3dd1ea2d720db293f9c190d8bbc6ab918c87594558905e484a7b892b72857af35a4803e2b1c19f61448c72921af70c5a4b1fd0807b834a8b3dd114dfa00038de13f976ce51cd4f7ddd2a39819da83c91316f97de944660a431e01eacaec91de005d629ec481e6e16d0f39c2d44073c27df2b92829df20e50f3cb0dc642606179e1c63ce24fabdf0512109f79d9207bf490ab0657f7b9835c96bc35974d4ed29918c06c9b88815b14f6894338c2ee774328318acfdd722754504fb52319bedbb860ad895985709959dd4ac292c8982faf8093efaa3639ea756b0fdb78fb167d18ae349f080d7d46641b56ebdb6663d7a184917f403906744b23d3e2b5fa6cbe30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h48d7059c03b65198be0488d2333aacbe3142a912d790104b98652c999b465d9ebca07a64802e5c70e4c56568ed0e2a05026f9a47e31220e90a2a00974dfdc1f19585d74cbb7dd96656a2de698e45d4133a6f564489f5ed73706099dcd1e4b55a17cda9ebc42cf01aa9d027b2f46e11aea48f163a4b35464bf91aef46b7fa4f070531a19e27682d077fec78b90e9977d5f1dbcf12199e256c58f5d12ddc301706f0d60bc10bb6be63a4adcec1502f939a3460338dc5922332c246620f61021a64a66f45582020a44c62570398cc292c5dc0b89f066cec07fdab5d4e782c70cb9a4a269fd8c28da3e1f6e6bb2935a09781934cbcf25339c901c5e6e3a4fcb693c12e4c2b7d10f791b576454668b67869ee8d0bfb9627a41a14197ec42908779fbcb768a4f26d3ce96598e99fc04fb1fa065baff51d63eea1333b357eee5e8f8010d047e6e8fbcce0d886bd726c228dffe5d97bdd8c2fa8b09df3560d9c7574fcc558ddca8fc32e52b3569b889fcfb5c3289d403eae8d0adfe5f83842a09155a57c5afc0b190e83d818ff58c01ae5a9239209b97c0cccd5edc9e4d86179b610521503704d3661deaf07bf080fbadc166aa5f0d3a4eec31105c25705039e6ec84a1818ab50e6d1a580f89c1d13c0cd86d0c1c47c2bdded600607883160ca14d6b90108d6a9ce7aeca669b8e35a9fe18c4d588a199388b08a03d6135096274b1ec6314ce076659617002c463250f5fcc7f40347159f85da52d4f9126101b3f59a29de3c2f101b6336bd4e4b942ce7e35bc44eb238239cbe276701d5a11d10b85e2054e69e9d50ecb001b996dddc468e20b6be6524a0ef204241a76b0dc0b59d33a853fec1b677a4e1248dfdcbf854d8e480c1bb4b9dd735e558824b960639d4458d298d27bedfca81de65ae8bcb68185aca1a08b786fbdc548f942bc2e02a258d4ab2cfc04c5547fc5aa9e4ee18f514e456b62ce9683fddbb3bbd7ada24a23a61d31c27b6c61d9e7669d9d4cf45f8043c34477655f1054e027aacf6feacf0aa4c524c622bf7e0659ac910bf5a089605deae7ece3ff2e14972a44e1b6ed6f7ba3045a07e87d5975858611339a62007a12de618f68ac692b47c2c91a20bcdbcfcd3eaaed258e1e7f4a0ad1bd0fd8e911bb074c849c61103d366bfcac560129df6ff94b9758e5e491d8205e751b90df4886dafc80fa614dff7e6ff541a6f1499e99da0ce8d0ab0e5a3cc6608dd7d36009880a64e1e73a66c953fe76645c3a2dc446386ffc00951c7cae1f18daeb47cc8df7a5457a18f58cb074c8ccb286bbf44be2e699f42dad7ec99769ba09fa4ed854e5b7419662aa855e9fe73bdbcfdeb7046cd0ee8c437d8fdfb058f0afccf2d8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3680d3dcb7deeba8743198deb0e29fe2c4c47f149b971bb046d501c7e0b7f4e713d74333383a5ad3c94dcc20461a543d9bccf9df453828f5aa9e6e9dcabea06e3e5e02517c297052d340d1cc7368b42d7f9cb921bed7a0ab137ff930d0e27deb9b2f44fc935818eab03058d0b57670cdd4787eb268883659b62e707048961b56c46649d6de25f0b8c1420db7679825cc9771e3dfcae3aa4a8bccb613679da6d4c3e062ddd3b6eeade59d756ea288f6af63a800a1644cdb319c35f2fd89a0204511b65edd375451ef03dffaf65b4b603a5f232bc860579bd504ea96d838808d0e352857cd9cf9c55a17994be47ebe978d081c6a87357882ae73713fcc12a4d6c9e0899359d5f7d60ba493e47555c1dd785e6d10a729a5b3bbc40e4cc7517ce704d1dd2f57c2e95767c8ce3115ffe6c4397b7dccfce58b910503acc837fa68c1bc03b2c5a7c6f45e9b6997155e6b35011ab507ad811c72a8c7781b635c994027ec6ce94189eecb2b9e14bf6b6fafea010ea99f8f69b1c2f862075df1f3487f0eccddc534afdc6887742b85a7b3feec78967a0d6fe4e99db61e42e5506cd0d551493509797655d027fbe02b5d64781347589dc1444c2e52cde1cce1c55788fb09bcdc1bd95978b1eabd447ae23ccb08a21492f41007ccfa1cff9033bc117bea9c4537e054264d753a84de7c3ea5621b00374cf8cde1c4748c95b6d60eaaba15ef1ac76002b22aa35abf7bddc9018f14f004c2aa6b5c690b477aebd767cd01d347c86027188b7eb088951b433816c4e76d247d5a20c0fc5f50dc124fec92f3f3be1272adefc02fb21d7000a7123f0668c1a359495bf4f7b3340cdfa54161c668d5726984b3c5602dde497a0ed3513b56d3004b9f5dfc7367ad9fd18b19daff94a195dedfbed00549481c03079e315497bf09e823eca179cb3f15b664384e6d292ba428c88783afa1bb380496c9f63943f3a504abe0122b1b909f196915a80707cffc82d09dbcb06e7e17a943c6ca320044d5d2385cd283b888c35661323ccaca3ae5ca4a6e582f68486c607639258a741013f67f2ad6561fa76d8992bccddd5eb0eb3830aba27c7829e5d5307b3a1400202a0152e729b2f955eb50c78f017e7f02ff89e8f258963fd54b51381f2ef0d0ca129d999a0e50c3e015f065b08b703a36da813fdcc5312de98741ff58a8d20f0084915c7ed652926c91e7aa4555ad7c6227c782ce08003680706b7d009cec1de54f05660ea79be11dc92575fd14179c395a1cc94e1a8a43bf740d655943a76e04b231d0d4eafc62a8cb61f5616fd170757c1952ad415864822f30fe9d80abbd8f815cb80c489ca51419b96acb593ab9d699cbf13e148f480ef35dd8a045;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h137888294a1dbd6fe35b4b3cff1baa7249809a41a7e267a8afcb68f58445b5ae3e55a609a0b73ef4861f0d93c2cb8e9c5cdbf048da62229a60622828b3c53a39b34f968039393f50a633f0a042cdd15172f28e37d822f3eb3b5b264008bac81fa6b8c805fe51e5329e1bc4acd3f8342758c842e9f2c53ee79e6a41bb5d8f7c8008555f16783cf53f7c1cae411d0e5ea2da5203b2b14f44ed1330ca3f69c423e94d2d185ae29db0bec1672844d1e834ae95ac7ab830d9ae81c9892a729751d5afc76f940fda6cdb85e721bac1c4251374c84ee553c1a17411af90bf486d43ddb62a4bb5bb91f26f1625d458c747398f935109b32554ec20de634ca4ad91fed3f7e64d5ac3f1e7ef1b43a83d335cb7a897a48e46b3cda3a25d93b5cf05564ec2827b7b72bd0fe17419bd6388b7c5e9654cab3f03d6f1322770f03cbe4fc9282a7a92eb6f9fcb1d21d2cbb2bb55594708afe26537dad798c59003bb493b9c9e2ff3a89f418ea777a41df15e824fed211dd139dc96280b08d2002a499ccf95a2493345223d2ea564c73cc28e82987cea1fb13bad4137bb3c0a3c3d9a55f2cad689708bdc76c68ce2155e6902f88b9fd6f5524d44583b850159859ab9c4885ec757683e432d9cb01d52a9d8ca1bf5a99863ee97aeb4855e41403973491f061c1089955d1e11e9e02516d957e4717bc8574650cef9c377040fb14e928a95deb50f260490de3f9ce40494bb728034df16ce51162d582e932fe659269710bad01d0080744d342c0a5380a2eea6e527fd3a8481145b025ee6effba8c6780b0635db3f422f6ed2e33462b1fd9dc01af4ae473371eb123de9e3db3759586e45120efb75c93a9ee8ed3093fee08a08fc618f92ebcddfc89e4c86607b639d681a0e106b1f312af978f93e3363bbef23c9aec87836f54e0dc99cdd7f123ead6935ba9a3f13b0f43a88ad23b72ad2893dfb3abe73726a70d9177e0e14b00bf96a7eed22e80d49b68b94e2109687b47586430c0c2758f5d5be91d881a8afb29601d92af563f9af58b9acef8a8ddabbed6869d3f373dc9ec1f4e1be673fea41950a8b8a38baa083ca3b30d19c057f343caae81240df84a0d57f00d483b16c3555eeb8b2bf004fa16d9e8357aed80759c428a331ed20da9cf08608d5905b48e8f3c65ff068054159a85884e01a32a69c5cca630191c863a53973320ac629540f9cdb3bbf066cebd13590b5c3e04f23dcff637374e224f97aa0f71fe2fcdfd858eacbec297b3d719924ee5c5babb9d6a9f68db7f38ae23c7aa61161de3845a090174bdefce954e3c31ecc27d25be21e9ca5395f9be1c87d6374911e66a27ee4c8aa835d12729cc38c12793a10562409c5c26ca043ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h43857a7d0efa08db254e46f66e9fc4e2c3130d4c6db84552ab243dd4d8527c997543b25a6b0579ce0e11efcbbab512b759a37181d26b7ea9555f7a968f321f25077ba66e41f624d987bfa343b9577cf6dadecf0e1236076bbb56c1dee52b39d4a43cb4f790a965fd927d96549063aeded009d101bb18a08c7447673484a8c93aaad0449c216c0502f44e585a72aa1a9098908d954279d384e36ff74e07ef442c0c55f36f0ab2ec8ed3b6670df6f6ac6faec2a521dd6058dd8638e386410737d0a70c3fd8da5564525fd5c30dc4a99cdb2606334c4502f5595238389fa10026d862b9c09fc3e40c6713aa652ea748b534c72abbe893d68463c72389d20ff3686df438d3c938d5f352d0ea985a784034af5848b6d809df8c9ad32fd6db36a21856a1c38d95f8367f0de313cd851133e951687e26679d88c8790261b31dffcd3f5fbfe787bef01bcbc7b3d7359d0bb46b17a8e294610f900b8d3a3bd7586a284d341bc86b723c29210f6ac8ba8b5e30b05f147eaad7a5dfd6a05c6bc8f858bf33e569e1b63ad76482ca7684714ac60fccb99811ac2a3ff4c70ad894b312109ca129b115322626991494f59d300ef5f70d2c4c45092606343ea55802902d5492e0596c0f5a35dfd4c088883027838037d3c64573c7324faf8e542c9410f867cd55d74a27c75165016be7688fa911ae91e7f2a701a247860fc8c3f1947245e2bb384f2434006f2c439eb6d899ca87a6aea35b3a1f3726ff6be726cfea774dd0e3edcb889a3336399e9156523f10a25b9ad51000ca0c0ebf31f2a2a4a6c3f553c8e2bd7216d41e9f0effa9743c95053c7e55104d76f4a108a927bda610d33236dc14e7dc67fe6bb4b22e8e9e492d44b96c63ae03da725c957f6c21f70f8c66cfd923c8653aeeda345ebedebf027b11ecbfccf6b81a463673450877abed7815884c59443a5760aa90ccfaf99ccb0df675df7e06468989f79aacf17795e2278905fd878145c5de98dad4ea0213e71ba7a56dc08372e4fa9753254ef651cc06fd86041c0c88f545a480564245c41c23b7712278e6e53579f2dbb1b98b9d9957a03b6312385b67680eb610c858ba70bc65720f0e7b8ac5b36cdd9361d8f2d4f057e78b61084d2459dc078a53042b58298dde61da2a590d0edc347e7a2f7820c499c7b8ee1425dfeec3cbe0f992fa8ff1bc6a3042152d64a69a7999623fea72ee5c6f7c79f9fa46b308c3e96923c783005f4bbaebdc75c2a9be38ea38c7ab042ae8f00519a68407d15b1f82c7063379db8b82cdfaf48cc42dc6ae32b1a028c8cf57474bd007f6d7a2ebe896a7473c9c2b9d86cd39c21ba6d078df707c9be0d30faa4f4f9e2895e38aa026e639fe035ab080;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h108c76adf1cc7171e8db669d44b9b31c7cfa9ec8d60408409796f4a4873697578408bdd4487e1daece21047672396296fea5aa9846169ebdb0ad7378fa07b4fa351842492024f2194ca847351a1414f838de89c95771ca0da0778b2059e40eefa6e17aca5b5857254c49c646ba06c81a364434ea3904efbf70e5ebb7b68087cac58a4b5aa43f9f3faf811025fdf257309d4767a42f9766b9b9d6eaf0486b1ec67818ea02a8ebcaf89ce80e4e417c8413703a1d40cdff91e740578a083bc9e1565b0d4c80df1e615fe5477c85fc68e6e7a6beb647599509bbafd82352f2f413e5c74aaf7d92643a023fd503a6b823885c7e1188cc6c2880fa34952fa75052f6d4cd524cb3379ca27bec725a30c6b8fcbd181dd0153b764a99991b40467155583247195a6b2a085027453278e84d038b40b3c113c63d738efbd5c3120b902c28f585f25b63d8737a7d6eab6c96e9842d9ed151c2a49229071dca24ceeae87c60860da114e36667542b7f8288a8ac112ff60eb232ac29f4c335ecba3c032e71ca96abd21d826e0017ee4cfcbe6f4aadac9805c2b8ffeddcbd1c518613418e23bf05dfabfd4599449d94a52fd12e693c521d506462197f22522f2e526045f3b5ca0ab171e00f009ad3fa2c9d6e03c25e0803c50e0b141e2df1eb9497c7941b65e73755e87fb6ab50c1dff75433cedc395faebb541253716e1eb8e4ff26ad37aed5860e3198bf5ba4354e663030fe9c3789fb2c4dbcf6558ad84b016f6e84d21478f05035267c4ea9591a7a78da53e1898644387a6a3aee785a89ea09e0eb758cee9795f546d6c427f7acde94234279ae44574744db531d283151e38f703c4f3c732649b569a714a3b83c3f4fd5cceb3281e96872fb1a9a5c35768e0ecfddc83266f820295fa9667f8060d355892bf47a411ce9833362de9418820e3f5bf17962862981008b506031c7601eb4dc4b9e48ebb77bf65bcdd2ce81602cd06644614c875d34649379cb853ad55224c0e22097c4e5700f95ec288b87b8b326defe28a0da4c1b0b14e4c34fbc87a15275c0b7a45984df1cd1a94413a06b6330126dac8301b6e928c601fb9be38be595e354563dbf130c4258bd01f13c3f06f97ee1a3a23519e52d89d5060a36876dde1f5cf54775e2af94b96a9ba86b3c56b6296ff8df2f6565d123ed6ebdbbf5ab8532bea8672ae7046cfcb370d8b4f11ce8155041eba84b33f88a00e2af78bdb230260a556994117dbaf2de92cdd9d0aba54f4ba0f5ae19d7dff060e13010392a6cd4d17a29629eb50d0e224e7a15b28fc817e26f2045edd2c1f1ab6b589b42faec29fad4a0fec7da0ab03a79ca621da923cb4dfd62e6f344a4e4ee091e7ad7ea4a71e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6db347e02d37d17a7cf43ed345e564c957e5dc6030ab3467627fc1724b522e83f25d7948e57ff9b378dd176ede72616e77d18827d0824aa125fc8d0888eeb373df3c6eee9249ee25a7fad8e414173c0c2638d00622ff989cf36cf825579055370b08e48ee28f6ff64846c14d5d1c1e9126fad80ac7a9498afac5125abb3ae16aa6f13ee59b6b26430b9f725bfbe91bcec777ee5814a57bbd0abd16d9d8b55d615147f2387f19f300a46d0b737c7d10642321bbf67fd8895303d961d7dc7ae857b4360da8855b79abdd1771142224c35db0158ad72fa0e682e934e962cdecab5426ff665a015c5ef8ee7909fbb44b84139a58d2efe7c270599e0cd60c9de036dd02e67be80537ae4dacadb80941b730d4148993cfa3c0ebded4a988252c49bff7bd6e137e6a281aff59e635d7777d93c3b79276f5cce1a25182ea3126df244f2b902a2b1017ff7894ac5e7c273456b92664043142e12585bc5831813fb016b718763e82fbd5e692795197c27ab6abdae4be99be0cbdcc0afe145615ede98e06eaf183507dc376d0ed3e4d808a100e98ab8c6b51d4591e8fbf2e4da92e53b016c0601dd8a39f5146faa2c54ce052551b3fb2240d86884948a93de869c6eafffce7dbfe85668c28782cf66702dffdd05267f45591f08f60fed0a523300fa0996945f5a57773e8ac8bf29c2a4307f10d05777ee6ec8fa5aa63ca8cfbb3d6736707d72b9b6470755f4dc8025be97b0658003015ad74a77f021d828ad1c54ee662623c452a31c11c6f863373e8b61370e10973ac9b7bfee3ab1f64cdd9dd447f9009552d0472d5a1463538e67356add861b19a3f7c0cac6ec54d9ce1fa151bcedc216f32d575aa4e028f91261f4ae5a32db1476d4d61887e58dc586a314894c63e9f6b291c808426f584ff8764ac49e2da9a4ed1ceb4bc5644bd8eff0b74ecc2093c04a697b322bfd72b05e36313379b86bf419f4d873204dfd0d0f1c84beb216373e3d9b7d1c45ac012dbdc84de4d3d853f6b38f17df6af63796257c30c2e09d00574e154d2f6b909759e84b06b972d8a81a405451825299756ce2ac286e0831890633c8ff79bc3938cacf03c518000d1f0bc3267f133776dbce92d35e57e90278d32c51c762f260db703f01c3dfb2f43a82aefbb4d6e80d91ca2ea1510d1f01c9632eb89c5b81dd929d3f169ef8ef8ffec44d1dd92490ca85edf29d6e1ccf3a02212c30798eaecddf69c392641273cfbf3867e07365797abf22a88c5f930dd304cadce31661ac0e71b97ca3aa409be1cc332cff6a542048d0315d2f43f122a7a0a35a6491ac17f03a4531e867b981ad0098c61356d6592378c285d91d05a92b268f142b460d21dcd540f90a1e5bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5196512c9a932bfc46a7756aaee360b1354d7029ef3bed8d442abd2088d14b024c3d778b9b136e10194a4ceed37853fe06db0cb9998eb472285cb4dc9fed6c84a2036ce16a038b69705e88e31e233be0d9cf7711b5b200bf283ab6baca105d8f1b71f8b84031b6c23f8f5e3048bf6d40ed955316184d8288119304b605abe1eb917610244a058f6124fda07784e3c4516087bb3340c0726956c35ef30412af4216554b41891093387ddd147183a3740841ddcfc199a1bfa2e732e3e1c22c9df2735ba2402db59ca7e663ea2b100eea3c8eadd0a03888bb10a9ca20d81698c9899103ffc7b1b184e0387f752f8489c2124e7cecaa15bbd2c616e5e8b45c7d691888927a9ce66231bb5458e260ff28534ecc715051f196d230cb138cc51095f9ebb4d0bc7b1c39f1e7f266a69bb2eca731ec8d2fdd9dfb109a1ce50b3331af3918de3c033b904721bfa1bd22e4a0ce9fd2107394c005da8d4376538d82548ca734d18d9fdd59c358179faf0ee441aa4c616fe1fba772937b0c04c24f06259dd3ba79bf60dfda2ebfdc02465830ec3017dc0ec25efd60028a56e59c562c8a9ef11f7a75a195733da8985bc7a9b9cb259c6c5d911419907c25fbfdbdb359b24252faa6628bf36eb889771b2211af755d29c92c94b38bce20d643ea42a666f92e5b11f93373a42b7421cd0f353e73bed8ac473bf9d2291b0d9814210351a950394fadd93b84ce8f07a0c4c05dc60bf8b9c3642027159c1b5d98ce2f4123f3d2c2311b1be466309d562a4705dd3242501d311110f8984b219cc445f695d0a09454f719cdf627eee44a9b554b80323b437b5bb9c6c51275af646be11b36ae57703d7f4cb0c54bfcd5c556f20be4f553e3c4f31c6fc6d93247d6bba96b6750bdbc37174310554d555733b53766fc87d382797de71ad7a27b9b06e5ea78dfa69cf41184caa8b49a4fea35db4acc34dad7b3f7625b9b624edcae95e294f8ceafc757ee09d37671abe74268fabcaf997892f34744497ce11ff6dd39e97adbcffe6cc2bd242874378245c726a972497d05e272c57a95a45919e0aadabafd5c4a6d55d1a99747c1d703b363ef4177931a1cd92e567b92176ba6c6b0a8dc69fe64db61b9934be6108c040a366615971d31f6bb2fd803758dba9e84a4d7f6e03f516c36ac655cb5a77efe2e0873e37ac03ef5fc439c877a26feea30a2b762f6bff0999efee12f7f3f480a818bfe1005b68a11ffa13396af08387343aa61b103091e382ddf6c5e8856d716a5fe5ee733b15e54a4e49b67150b027fa9e2ddd52cb659c0f0b07d52bf8108185a1f53feb523f7b4bf2969bf6d550e71cbf8c09e9e61536cc7d10ccc1bd4f937a7170b518dd94a19cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3be4a789c11a3e2924b666505814d166eeb3812ffea9fa18a2b5e07a2da40ef275701819dbea84a57bf06d55d8fafb27edbf3f34a14ad6832a0cdc3edfc05b3bc944d5619b2c6f847c2478192c7096ee8a6ec454549dc1f0eb56fcf1a026292fbf552891f86eda77f403e3f582719da1e181323c9e62ae79534c2244599591f02d9ae7da99147beeb85c0186e30c600067720164adf67766769b540f517d022e605786035d3a52be720180bb5861bf341c35e0e7c68d90b55c1016422c1227f00bdc74bfff867609b8ae6b25dc44628dcdfda2f5dc2245a0af6e3a5e98043f6a1f9ff8b3c59cafef94e48f28d4279c41dccbbb965bb38a46e7e4e9636dc61a8567c10cd4e9cdff5166a971209ecf5cb7267b4adccf4f8ed18944f960645046dda4a19d5d282eafe8b67e1b01fec6d86b301a3acb8668d579804f5148ff90eb757fd3520ee6eb9dd7255eaf61098f5e6b07446a40418d9245ac548be913c4e279a5a0645fcd3ab803a92ef5bcc7bae16f9962038173249be118f8bd4152fc54a29fe5cf563b4cd70e6c9752cb7170048b9da8db17dcf155742cdd8f5969e624700752a0ad1c057c0945a77ef9f5abb06c0033c9ca11592987ac2f2aa26255f03649ad152f2d1f488c7d910ddac8b2a72489e0a42c17912342629bc168cb666ea4170bb83fdc84fbb84f0f7941bddf4b56ffd868ae355e486d26c7a41432335a3c0bc29dad54d889227c16367473acb7526347d0cd6f278317a76765621cccf1266af90869abd8d22a2924f96f4906b5b8dd652c547b35264f00b649e2bf776fdf2a53741170b2c6df15c4b093f7b87db9aaacb1c644127793d9e86882963a441714ca8ef64c3022e2773de5918ad62c870a6d6c16e13439d936281bad3b9b3409527ff72d65333a2bf5ff6557a3c0f0300d070b8ae7ab5cb9a7306279e415f63faa898fcba0e5d450dacf64c8b641beb21f6d8d56bc948bd5a507b1d3cc50d5afaa0510868b278400fd8e79f370e93156f19afaeca3ffb5ee33ae3e9b35ede802afa58b6e4a1370fd28d2b7a997012367e09e4d7e2fc3ae7237b18fe4b2064beb5d495d4588d55336771923eb9ae9333f904775858d59e89da073e9384ba6c1d2b25e53a019e6c1b1fee693a6602eb0293a1a1dee39eaadfee90660f4ca1a4a69fc896fd6a9fd04be897100259851559b85534b1c02fa9a7c5a09ea63fa581f1c2bcc8a910d31ed2cdc9b85527dae8f34935bcee6e0f3827675800b12100e9c73b962b5f7832edfd1505d164143e12813786700f320b63a8da1e2a22f6d935b82d9dfbae0160eea5ac436cf0f5c9c157a214fe3c6ac5efb03bcd2ecbc25d7ae6f45a892c2dd6763b2a431ff7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h44792b291e9d708d4ca58151eb6964006851be9cb483cab54cb7e23f7a56f4d7409639879034cfc0a27cf10ab86a57a0ff4103f62d1934d1c5cc17c2fdae25fa4882618b9cdd5a6011e1bae07e46e39bc40ca0258d5a8ec3846233e5df22305b3f8307225e712d88381e3d4e89daf1cf9c837340e671a883237069b68710832a3155612f7eae06f2f93040340e02ce591fc2737f2727e099d8769de8997d94113e4e24fa92b39b5034b6c3b0653960b0aa459ceae0841cb40ef5b1c78f216ad012f1730284175ff401a298c6a691d241338fb4ea9c4f904a3c797ba0f4cb67c71b77ce69f15932d66d70995005b9c7328bc934513c040f7914187093966064493299c228e08046db474f2ff1ec841b4e2da5643b24b9affc8ea628afc436c228140fe30e027b556a3bfa547f943bb5808fa8ca7e99f58db95b71cc294a7caa8b545625daec9474338eb6a9756516a69a4979408e16ef118f6f05597bf9305a6bfe6681ff965636165bfa1340883b6239c029be4da00f92221330ea08cdbb6f5ca8d101049fc97e6165d896a3282453f40c2277146aa76816f91736fd3c6ce04ed0dac76f2bd9c722da40faba2a3c02f30ceadb3697693dff60ece3b65f5ad0dbcd4a558f02500284adeffefeb1a59d23ce063f9b6516c864f7338855f8a3fd5b2394eaabe6921389bb5f738b1b16a393c8abd64fda096713454ca79a1d4707052f0208bf5e056e8a5df89c6012a135e4d5c5026a134c92b4b4ff3e1850db0eb357b1559d85f501ff7d796a0d59df78c6af4a271eab41f0c3d31e9b49d5915cc78181f9013e6f7bfb1928627335c1ebee5ba2a6711fb5667bcdbcb89956cc1edb50efceba12633d18f49c09251ed5af4b2a7dd1047f0801c4b9ad14082a31526d7079123e4dc6d92d414d55209556b772b2fcfbf864f0b874f140b596522351451e4fbf78f61d708c4eaa8f7b25c741fe6eb99fe24e51cb84662523a03e975df8df5eaf7a45a8826f91b9aa0032d9ffe1f03fbd69c5d0f25ae068d1379845eef0aeee8273aa128dfcfd4e971925251571cbb871ee25b26624152d8335757e6d0a7e2b1e09860d4ca7a6f4712027c16ac1145e889c2336ac0d5195e92d02bb71371b53635529fc971c462c78b9f21ae6faff28e17bc3573f2bf4957c716675dd913d6e0561d49d379613bf2b1fd86fb7722d9827909e69458b116c5a7266746b3fa1900209bcf78779979b2f954a073829d76baf4d149ec55791b7d1c35be34accbc5eb64f6947911935dc78203d3fd065260a78ead7b4870f588e3b4071acb27187156fe99a76aed5e0e7e58465c12a8b274fa1a6b67f6c6c3979e14b741dcec41acb618e21f9a232c8c6bf37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hbe9d853e56fb35549cfeb1fc1a2070bfa5208ffa005c8c4d34d6780b96a7311fe2fca0fa54b3a750627b96f361372244fc962cbc2e406e9ff22246794ded55244437f9f92cfe3230cbeb84c6dabab4d0dee855fe106330bad909ab30a5bc37f46dc2def67bef7c9afcfbaa9edd905696e68c72d86f8276c7669b6a2443ea51a99304dff940c74baa1d97d3da1f8e6a3eb04314f580ecf0e2ebc0b5f6766e77cccc56c77d3f5dfac6b128cf451045b7b1136953c00093efdfa5c6eaa932357c61695b72e3b55b78023565133e1a3242ade5ad647bc477eff167b8d36142afd5d846584908cd3e80a1238b3541ade8d6f52c0612b57a0be90a2d62947dba28710642c64f32f3b83785f7e5751318bab360e5ba37db1bd1dc3196a8b1620c0346f3573f71abe2488e693466e47d8436fc5aff422a7b784165dcfee010349a4cd1ebff7b1d635e769035f4d0d6642373a54f4f1e0e3c8a81349b3ab9839074787acd1c6870b9cad4da860df9c8a881729450da0a5976ff3fda0bf5182630fa02c0c6840ae3958bf8876f2d989c53c4bf0a636bfff1b866e109bedcf8bb61c0a2b7289182fa7a92e2728a292b91506b284a1add67a133aeb4fb40348c23f8ce0046a4b61dc9b98809ea3a77ad33985c86a994ae0c38739ec39bc383982967f43bc5c5a482efe3e0252ce0f3f233b142290dd152e4b83b9e66dc0368f62b343df4949ddb725107303f6b207ee65ef9f7be4419411b567927f3fe72b37741ec1d4563e475024290f60a35398aa576594856b6f4789d7ed6040d20da9c1851d29a4733ff858efe716ce0e988f16e014d660ae08bdf512b281ddb2f5338c0f5056229b47412fd65626345f5d7c498b0e4d50d8f18998f9fe2219ccd724b78c6f9272a468fbedfa2b79fc1b787992525cdd93424ccdecfe1083e7c222d6b55ecb5dde2608c24cf86ae6df2b17dc4cab16f4e6e3150fb58ca9ae362b8961dd2fbe11657de60440fbd76b84c17b4086af167c820a4af9e13a73de613415e6dc0f055625048cede2cc102450edd05c1aa44e17417bb2b7b2254923646dbc805b4b594bb4b0132801ad58104c5145dc6ccefe64e0482e718639403bed2561e3a60b1b1d211e79b5127f39411b9a78c5d5dae48d7c832831cf53539683dc720ce6c7a0e5688666fca3e29028cba9d978e9632083c60c4a1610d7f6742e61fba8d1a1c73134e9aca44b61a304914aef4305776d94c208b3bed8b22e33d260fe7e8c928216600c202fd790d59a04575d1e228a61daa908109ee760c49adcb3459985ad9356a319b4af9f5b4861021c482581d9d1dff2bd7b0dbb55e0dd450ed78cd612f6a05f61e2cdd3b6bbdd927aadd2ad0905f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h238737e4c41014beb4f4d8dbadbfcfe1b365d3746324b99c1e85ee501d7bc140fec9e9bb61fbecbb30daddab361c95b464383baf57431727fb5db6d1f0675419e4abb1c902fb400bb934ad9e9dc4ba1b29634ab095b5f59209e4e61ae24fa7d6bc1a83159f3869a8484fc088944971c9e97c6a47e1a79413000b6ea28c68668f2e265c5c5841a46bce8395763eae979d50234bde619d27f17d1066fbcd65a06dfe76ac3622cf0837554f65f8ff90e774c3232a73e6930913a213f91a752e75a0f7ba87934feba20257e78ccc56f2054a4f1ba9f1a89c4810110ee154cfb07599ea5586b63008f571ebadd1e3d028eafe7e4175b3491bddeb2d5068adeb5e7500db557d0c46f0895b7287d95ea6593da26026a04b9ee1d30c92ad5aa74d707b375ca007ca416f598e4b38106e44460b2b2f7a65eabc82bd1b0c713d27abebc5a26a73f7f8d8750a862bdd039c043e8267824d54157c2bfd9257b7c79a645557f26b0f60dad3cbb53ab962bde6a7801f8af1dc6ea10669885a09e34357d122d042dad417697b3ed45637d0ad7905f91d09e9d548175cd7ac096ceba56d800d89d6267124a1beba72719c32ec81dc599b9893c7c4474f8569c7e8f84e572ee65587dd424de6e3962ae35e74453933fc286ac845ec6eaf784d00892f200983411a826a156e4b4c125f431144d4830e5a1e651d6b0fec48bff5a346cdb4a5466f5d7999235da47ed313a745ef0371eb6cfef38e93895a3c9dbbb9ef61d7012878374b260304798cfc5f5813d1b74402667b5122bea32e763a538dbd7b57625a6de9155a78d54e058fc736e946d23b25b001e4f37ab533190b4223ce4b239f9047bb8493c4b1f7a1b6ab1f298612c8f11cf693904cc3f05342d03ba5147be4e543b5251770b6f1a18a654af2c2083dd85eb697ee2215a17ab8cc3121a5860fd762f9d4e6c59684f4b420bcb24d61ba03e81ec25e100138fbe0f9dc778581c2e18771c56ac98baf05a0715bb85e44903521ee8f12348516eb8aa1709b3054476a7699676fc0921ced35e3a4be7b27cf17e7aa58c8f762aad426591611055e0a5e9f50159705d6d6767db3cda8de9681529525bba4be96651ac2b2ac4e4babdebfb25a601abb5b0542a76df060c493c8cab9dd93c9ff2ce7578b57c9d546ca6065d71f6d74c9ef4c7ca6b66b4ab4ac46ce6658a17e8abdd9029d4b8461a6056ac61bebacb2f7ade4bcbb53d2542405502cc033c0c9487ea48212eab4a91c95a9ebf57abbd4a13911f452c7b6aa1ada6f06c7932cb4684454099f0ce5132169986a166743e5ac411bec5e43049d95d0b2ff89de1f1c67e905b93864ae1bd0dca1f782ac414c9f1409f047ce631ad6d661;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h450d17bd0e81741b0b1abcbe14e2ea0dc26b44aa3e8b326702825d547788f1194a97a80a5c2919ab6d8ccf3e4c9be2471bef84beac14597dd7a3c5b5f25d67e7dbe516a049a937065efa5d16d023bc3ea7ded62d71a8b2007febaf2ec9a6840b3510387f95e7b3528e47b6e3068506c729937570f261e430c6370380647037ba9b003181f77d58cf887282febf259b80ee39b7e4f810f835d7f699ad1e5238cae683091ab856a67086488b3d2bcf0178de560e164f0283b166e50f8ad7696b1580cdd08f295733610239f16d388e7c833d9c044b067496d0035ab8dac4b5b102a881c134a38cecf9baa7e7aa286870a5df8b719f66c74996ac9af183f9e434d623faec1867be6c9c6fd9f350acb0bda0a5e5722a6a89e3bae10acc5c4c5d898adf95961a95a265584e25946cb70d0e1412833a2356f6c1c04968380db07621024d621546e84522a322ecb5c7bcb4d93a99990a4d9668a807fdffec5d9fd4fd5b0ce032850b677c44fbfc679e4a20d6e4a25de1ba77de10afcdacc9917982965ed48a6e3f3a57761b626c55a25c35ef22b7b493fb01fa2006e68aaa548cf1dd9765c0212364cf366cdfa1472c3104e8d95a60f9994b7687b36c0148e05cf7a889f192cb9bc82ade1c37f1543f56100e9aeafba04234016213f812846fc6ef3be2f13aef6fd15c4822ab6d013e8daae261f52d6b7f07abb6c7f92e5968f6f514b3af12a62022d36f46ae7d017b53f6ac968aeae44daa0c5da66abbc880ac210bd6539af218148811e292ec0ecde2fd040a2484e3c513540c3e279f2e5bbd9f888355530b014da36ed199157f032dd8d163e6ea22cbd98a1cb7c0a2e3e15a76ce63d16fe22599eaea2b7baec506f8304ef08e6e4d38879ee7af7b74e7f24ff34bb705267bda0f9f6001975101f5dd1c44620be2258a15c5a977797394311a0f0f857c81d43e34772017ddc48d695c36460a73222ae114c1bc9eadf038392ccce3980e1dff96e011905a024c515185ebd11c8726403d34df61b6792bee3b82c5782b26e4f0c3709395628bbebe2e667470b71196d45537c40db49b2043dd934ac9af7845646f947d1bf9966f24a997fad0dbcb6b842f95f5a67e8f37cd29422af508eb8083592a4a4c1e3822bc8c86122dae3ad0f642f621121ceea76b37d6b10ae0f5e7946d798ea931126544c281cb4768b878d23a889ce50197ec666a05a5f9e879a9198eb0165c569cfebbbeaec26dee7ba6d0bec146825167acbfe5f6db5afaed8acc07361dc5d1f4350602092a14dddfe6a31d976c31a7fdf1189a2c54497ad70a17e3a5a49bab66e7a1422bd9b7ec62dbc6e0ec8a3870561b6a9b80a6c1e8dc4be9eca96724354106ec20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha1d5fd6e7cde972fba7277f96d87185f080e9ca6c1d8b3bbc15a5807b2696a81baceb150597ad6002333689a493fa132279b707372cd81dd44c61fc319aa5b059fe8c822fa426a5ab0b4d4ff5feeee4e70662ac8bd0716e3da769d20597fc9ec30724c64007d2311a964f8cb5c63c3317bb8e24fe4d65650180453f52ea26ad5ff43aa6df238031c24c1d2e50d46df98c2f28d0468f27b98a84aba8937f044abbad9acc995b2495d9c765a4b0fdba43ed07b13b23e40b1149c42b82a3ded7b9f20592797afda6d8e0df35a2b94d82488d509f4252b5670e3bfac2fc50d8d3e686f66678cdf848e90c9879f1b3d4c7ac9479caa757860bf95f2df94bc963a2691d8e9638816e7143509f1ab282707c697abaeb387cd669baa71ba84e575aab5ccbd7418aef5020e0b99dd0ad789db59280e14cf7faf5d3cc736d4d9ed7cf6316055a18149de24cb312bdd7eab411467bdd71ab17ae0c4f9dc605e0520f637dcaf8e9f1f092380525223148b03fb5d08ef0d019fa6dcf755f6a126500c76b11307876cf1bb0c273e39397f1241f00fa9d07ece4f1329c70cbb38740445216d700ff80fbe66912ca76d7f788d7c4ae5aed1b017ce6bebae8eb081d456616f7e4ed92cda6a86908e8ada4c794c650509e5bce3ea0347ceb0783a8b52ec1200495107428b9846ce37b408009827463ca3410c1c69d1e72197f654aad15a11e5eaea586024780472825a3bd0da11eeda52331ee23098091a7a8d6e282a037ce0f07c3f9a243bbbeabb8c0627ec59e0187ae20d1494c6b62085f81d5b9cec3beba133240b2e35ea8f46462cdf35444bf7001b9bc477d7ed5f20e6a05c51e89fb21713ea8f602c1123b6dd6c56819e9e0595a4204d6e3de460426b497ba3c8b509300bead517893b78e540a3fd9b93b14bb8f5c4167537aa8569424b6dc5434abcea26656f03d0030be5d048706987267831ae13a928cc08265c8a427ff331d05e94a794b9b1f15d36eb350ee8af1c89e42e6059a57439024d5602cc0b74c67598fd5c59773a0c6575bf6c9ca02808083114f64826524ef38bacd7e063f67eba4c799e14f70cbbdb64cea2eda44c7c0f9779caaa6679db3171c446ead4f7de003e7eb342d870aa97dec87d40b87db97fa4dad00ecc082571ad4b18911158bbd6bdd8266bd0dbc3031dd10eef1ef5511f0ece1cc71bc2a366f3accf5deb2e7c400f9e99fde80bc1dea037ee5b5953cf4778305d1d80d45280f13f2dac8911776912e3faedaf336d5d86372eca9e0049b960eabf05618ed46564fff65a0dda935572e6a36bd62d0c1603ad7ae95a2b712cc72c8c0f191f9ecd866014740aee2a1c81892905cfcdca8633b7d5c8e37fd4de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8e2003fbf45946c0bd3555f16783627afd9f6cab76d8a3186d0e931507704b46bb11ccc2f6f99040d30a18adb31384e616033499b82970c7b15de866453218bf8895696340ccb9c47d62eb75c2fc0f5e9d949afff0b3b77fde0c24719b7edc7934ea679ffeea5867913acf0dc71d7827e174fbe35d538aff7af4ecbe5b27854f8ffb70422f88ae38382fcfeed2e8232bd6f71bcfafa5dfc7a77a817c8804efec168907b51f4f9ff53ce590a28241cfaddf440baea0c687336b3cb1a2986c225250f65badab71a1e1d4cfe8843939376fe4bb68b3c7b7566e06a6b801dc042c81b92fc36b85a406b8532cfa62786bf7d324763f805dd8a907bc79002d609194115e825b378a561e3520c049aa691fafcdbc28bef504b09495644c725afa59f0e338b255ace375ae7dc63a4bb88b5062ae7d6594cfde0db096dcbda81a8a654884bb770668ec4c6e5d813cbe3999ff26b925001da8505e73507bc8a2648b87da42167b92ea51ecfce407f64a376ec5dd12d6cb9c756cedf716b2bbbe01c4bda4673652ac1c64daa9f06a0f637fa5a6514caa6003fa7b93a359573fe8afcf660f56078326b0845330a173eb6b57396edb5c4480ae21ccd076c128567176a47a64217661f8e85f8e5d36476248db5be0705b7721a01369c45a07d20a6f5048756065c933c0a49db6af752d2008c80c821bcacb6a8f2183e327eebd5b3484073f02b2e853eb10cac862d81f0c7850fc811764b4985e5ead933473505b58e58ac601f207e925849c524183492176bfe4e4898394b88d7236a9c26c0f1c18d71682dda49dde824c2f24dc13fa37186da618ce2c7d189b1a534ae1347e0491a4e78975ae47429d72945f963272082b8d4c3294491eae40a72f9635423c764961aa28fa53696a56cf244456377706ee506de0abf46128d4df50e6594a09d34d45dccbe0dd32727a6ef45a6822b4203863c3becd5f97c5cb62d481f505f60b1778ac163145a12b01735768a8d3ebfd350ae17f0af0b51ca490cfe5137eb7c79426a8bc0f6aec5eeaa0904ccabf0a19373aac13572233402514eef3f371971c5a652bd93bc12fca60553ba2a2885816476e42c89f17f1bc1b8541284764e6ec678a22f0cd90520f3b0e41ae40a0b4873079b07f2529c8e1aaab19cde53dc84c077b8138443e65a7fde2f838489b70d8f649d361f6c71fd73e85d98e7bcb40da0ce9946bdb82d74dc1425dbb5b26b0f8b087e11782318e50a0a58ce67a3d80d6f7f3c9fe52c12e6d38a1d9e41989b0658a277e183d342592e5e2ed6f67fab6315adbb94e2b565bce8d54e77944962db9099ab2fa3b5ea66922fd5a8b803a4977b775d440f6ad8b96b3502ffdef7ad54883a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha5e513605d1e3ea87cbc07537974566e935f4d9ea04c0a1de99644747275036cec6720313b36894c2731f7144adb76a297351ee3dd28ea204e1cd4e632d377afe9cbb8be75981f1d13084801e411c7ac59768e1dc575e9740bc56e31f90160fbb976dc70fa8964d8f6bd8021c2e4b65a70b52bdcb040ff894ab9cd69e4d8c713fc32ad1ab1fa79c4935d3962a8f06c5e5b82f9094a4d79345982149718a9a2383e4dd29e2fc172aa1ae76651387d438ec79de2b692f62e7858cbbdb4e5b1b6887417b31a0bdece1bb32d62a6590ea4365405e3c95526131415fdeb9597de412151cb90de87feb2c284ae0144ddc562bf2fd063626da5af279ff8eda00c16333b656902c7762d8117359356a97ca04b881d4c618f104099f2a242dae91562a3ac38c162c9c0af73f9ae971a266c7ea177c1858f8d0b519bd122c60a9b1b279082dda7f5164ae0b2b2b378156e543edda2b7f8a21d3377985e3f692b39841a49f7156c8c36b8a97b15eaa11aae0377b417debad2470c88d6ef87871d2398551ce8f2c29cfa16d91c3e54ad23803e5c7fb4e4c9989f3ff141fc7b77e847c06644b555f53bb354d577981719bedcd6b9913254dde7788c0f1e2d2109414e6d719bacf496d7e3fd4880b6eb9fda88704de791e0ae6ff5cf6168e4d923a1c30fd5fd34f1255efda2c05451de205e809581272000839edb690d69ca71e72e29b9a4280f15ba7c495dcd116a91b387162174dd0015716ccb1df508ea3b972d72b0666d997f94bf283bc293fe0e17ec0bbea17e2d3ffddefab757577873ffdd550f06754861b6ac8310104f10a29050ae073acb3b84fa6938ba3fce1b71ff80d648016a763d6a2bdb32b8b4952dedf4152dec10894021dea723454d970d95625cb6bd81c063a913e37cb1b9b1287bba16b59d0ba1326129c5ed330b9728adf471b922d75b72514b93934269d80c765b662ed586e5e53eb8ddde45d7c0f86860e80fb7f93d275731da22f5fbecdf93b43f12bcccb9da4a680e1893fdc043b5894f38806801ac8b55bfc59315d6b691b9c53cbd4649ee0fbf9dfdf2a2364735d502077b00e0706f788dbcab3964c5c5d7d0e656aecd80e60fb525392712005a4f45f7bc737e091411b6f166f30f9d248a4bacad08c665ab01c5d5af60b222858a480a62239099e6582d1f252856f9c9255967ef09bfd049431dce9835c238b336a18e9d51f355cd96c1ba372ed7dadd3e7619e8efdb9537eb0ba551065566bde348e6a91259cf65093bbde4e957708c7665d15e6f2f73386fd752f7ef035999f1eeab79374a90a092411d89ef10296a896ace0a90e10f2dba17e6700d605eef0d9657e6e0cbae89a1e65578d14c8be237b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf902813d3b7f6604fd7f521bed3e042566b0ad607b0e830ac9f54bc889178eb8421a70e61e16f5444be9f899ac888f31902a12c8b60ea326556b819d00a1b192f343e1d3280ea0c5f93caafcb4d459e17c7e3c569aff68758717b4604a342401d93a414ecfe9ff6391a9789e1a07264910e8d1b12c2ffea926a0e467891210b42ab64de6ad4e034acd4aa65ca2d3d6f2c59b6d356ebbe9e862ef8937ebf994ae5193a84d2884ba47589ffbc30fc7059d5e835e5a9e45f6f9fdcd00d14832fbc82f6d2dac5556c8a81a5c468b8845d02f210aaf8e74122fa2840b0c867ac7d59c2f206cae4dd19926e750130ab9d951a977d0a490b4f7083f4abeb41feb3fd94439acffcbcffa82f6eca7a1bd7e51bea13aa6211066cad18997ecb43580189ed03341abdf9754d3aaf82ce8338a5b6bc7ce329f3dde89700eed459aed6bda9235c96f2591aeea6f70241cc43d7459c7f897c50a2ce5860111329c2252ba1bd23f37135dd0ca9e759ff1a2c05c481e4da25bf75ce5ce092a63fc3155422d09fd60be93ccee015fe1a42a146964183e3816be178407813202cf07af46f725dc62269e51e4e048cb7903bdd12be7398dc81fed6389ec683090b63febb8f49d219d9f4a7f0ddcf3332c67b627eedae842f6c631a38c59f1af85c64cc7cf03a7cb761b8e2392f445bbafe7bfa78e82609a2d5f9ad1b5e6ff3b16c3c93b20245d3a7a8e286ee116fae5189e44215fd2ed3fde6eb8619aaa7b259b2df8e386adb37ceaf56b555c767406dbaf6c23bae52f4690b44e5412c4f2f7a68e07e86ce6453580e0884aa388c9fa468ca1b60400af137d4a5129e467612d5c448eaa506d102ded604a1a326e996ac89b32fa8631a53e096c0f15912d74a1590bee1508145ceb1e3c776745515a18d854a7d3fd21571f188d60c076bb164ac2122795833d133da8a4e2d610372344b21120ccc5b77386291c2712e548eb0c390ed1c79e920c674d3b4be34c4854d0ea498494a4b5f3104c510a3a288981ecd53bd5f654396222f073cacb2bf34e8e8ff6337c9af043dbdbd36ce2cb8291071ee4056af4f06f47204fa1a5843a0ea53fd7e5a8119a92953015f94391392e1a2961de83309c2fd0808c7d9feac9a2f6881de96b91b64bb5053e076355924521da9e19724c09a5b68653a25e23a8baaf97c102d7f9d3331c4ab8317d571fae7aa391b106979c026cbd1d8223c11413e143a03f7f07240bf9520363cb400e6251123d8f61cfe2e40d4a3787503282dcd5f1e49436730a5091eb9950b43dd0d67557dec7f698d05bd14bba01d9147d4beddf58842805a28f2178ac408b545d4a694d3add057a9ea6bfb21eb3a887cc3b669a1d7bd4695b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc0f833a818c81235344630f7fbfa50bb1b2214fcfd507cd74646a7e26457eedffd6e07f9ff90b239578011c9c95584f72b94035a5582dba2cce0ad66bdb41afcce97416466b951514b446df7fcb663e7bbdb2c209147792dadefa13915856680fe9bfb0ac9f9f23b8ca7a558cb4721f80058e2a34d85ce3046d00e775335cbdd926eb35b1ede805d49e3eb94f1842f5794a164c363283e9e97e44e457ecb6cf89975df6bf268d2ebbad2e0b68e638f2ccd55dfc607d0c88cdcca26d70f34470767c3938dbde42cc8335141c6135b8e5d35d9d36998d87ec7a418f704e8fa216d06d3562d66816cd000c2934fa2fe5142e586dde128d946abb02bdf5c01ae423cbf502b5749d65177c80b7fa05257ca9f07b5b16140af2e86f20ab580a1a3a2b1ec86cb9d823cd4dfc02bf282eec2e82bccd5070f318f31e163061598d157592b5f546118803587c42f8055788f40c2d68932d1644f883e66b78b81f6dc94d236c7025aa6966ec4352a872046709485a2e91242b49c1597ec4c2d7cf7474891be85283bc2a2c0146ab07c69d2fbdebe41aef17b626b1105db021760f312fe5274ee9031c703145c547d44770f3fd309fb4bf36dafaa840cbc6bfa9b61f1ff9246ef6a10686e29e96d71af38560651793d4f22fe6939ae607d6d293a491439897ef6bb34bc021fc2ad62b290e11968cc70b2b5e6d592176657e7375bc3838a7404672b7449b86e6d786e341a3b1d789724a82b900861b1c80bae2af6d38aca41c7776eccca41556691d61073c8cd3ff94ea7429fb2e025e7d0d62a5ada24b2d8dc7d8d9c5b1da21698a7b0f3d8300d5e622d0f38ebb8f3c0018c9b4eefe730092d5b7c327d4d281d48f5deeffb9102e4a766853c36fba8cd74540c050fc775c2b7929804389ed7b802d363a30d849d17f6b5117c21f855256e9667454872bb93d744ae2327fc02db6ae9d91f103571f77cadf81ec2df866d87d8a8994764f003425c04c91e6de4459f45f53c97b556bcfc9d3b447eac96ef926566def94f3e4116f6a0d4f7f70fb3b7af40e99bd9f827264a7209cdabb3cfd6a983ac619bd229869974d0203d5d4ed67434fdb821dfd21f8834afe90720c370566af2cce8efcafca5492b4c040632f465d3be87e245005f88de692cfef47aeb80c62319f1545a6abb290585c05fd09b54478e6f44d7e6082a070d67285dd6d064de568f81f66b056306b1be939019adf1a59e97f163a77b3119e7ed3de31fd1e60101ed02cb56591b4de1e58273a085bb0877361d86750226eca0e47a550cc6ea2094b7dc932d3404a42d8f6233ffe44b57ac0928975abf5c625d5616dd0818dca39acd665c7890989a4afc729ffefaf44039ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd8e25348cdad2f78111b2acd37eaabee7c82900b4f55c6647118b91693ffeaeab527e4222b4ff95949224cba88f275665e26f66ca5956e7eccd36ec99cdf5ea222aa68cf0ad2fc1f43ef63dceff8429fda2ab5577e2f2982afd737eec86059e379e12cb12be86b559bdaf8c2a26b06d0b78f982d87861fdba82fe70900346f3ff150e7300991912d4f9ee331d7b69840b3d83782a4d17ca4dae83b6003c64702516cd82bf25bae2b7f21083a836e552bbaf2009f8a96f4d312dc260ff72d96e3d86d54ff3406b3687726e149862cbab08b5d687a311c0971c997556aee91424d1e0059cc4fd1082bcce28bbf9f38c1b46a82c50539d99858c434f0c69206fbfaa4fa74484952de37a3075320d9e002d50fe5565b0727b03a510fdcd919b91d4fad51ff511ab4ec22a2ab0ca6a5521f189ba294a3d52a2c6a1380f8f327b0275d525cbccaef537fd095a5448ed852e30bf001827d1460f1a3f3ad8f52bdcc5cec6eb865ed6df462a38dddf546e36e25d91602b1ccef379300dff58b9e45d9f4b012e496e08ee8ffb295992cbe0e3bb20b4b54d2288c2d9a95e30907df0ce9894845daa0b44922b074c04caadfeb044271c2c0f4c69fbcfd513ee3d4e68a4e6997c44c0e83daa8d3a87b2b7f7e34cb667abe09abc6e571886ce4a28a83f02d5eb6992e09d0021812c3fa315f65ff8e01fe3d6de65506149b7bc1f08f24145865f0dc4a6296a18b06bad578144b2f9b23abaab218e5a60ec51f78401449187c1efc4b0af967bddfcddb14219bc357432b5e7cd56de12a67e0758e4cc0cef9948261e81544b86ff764aaa44e3be07fcc2280070d62211617a0426febafe10a8a43f1c90dfdff91b3b77bd4dd6ed8695a7346276dcd239ef71ace539f12a1a9279c2e63b75b5a483344067c28348254f18479ef4ac852ffb8572cd5ba3b2589b2d70a9d9dd36b59c824e5327f3edaa013ee878d8ac675ce77260377b20779f4e1bbd3c76aef1f6ecd07299997f7a554cd1487e44ae5b8b0c1869527f19ebb9956206349f83c9cb2080f3c2e1e790856a6b4113d3b9e83c15e8ac56e10caaae76b009a1522d86b4e66717020e97e6d23766cd9a1a4f59b266b1e4e653a27d9b31944635e5d9c552a02a45a70606006813b3ec7944000ba88e199da74ab50f698378570c1c0aa1e4860374bf39aff70177427c2b165e2029590b8bb168eac3aee510fbe8aac331f71d030b1b73b711e452acb0ed3c77f71d3e7623a5cfd08921119dfe52ac505eaaceedbe7439a917d7bbbc54211e066b3134eb5c6727a333c290564d1d36b9583e002a9c07c1ca29c67b45110cab6e56a7d3b47451fb27fc0b0d1925fecbf782b549b1e557f7b0e68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h74ef70cee638e0ed6652d813e3499d66250f18a678c10f57a6a41e98c0ca5fd05a241a5d50ff050758363db3cbb46bae0d1acb3ff6198d21d2e0c22d0a9aaf2c91d47cd4fc2c60aad2e4fa623f7d691231bad3c9b4ad750be3532463df179b93aaaa90c31f892e0f46eb602bb28939b35d98cf140230e5d2587e75302acb262e0b34c0a40c7c7b7c232b9cd4b9d54328f87ab26fa1ebdc7973a8cb19a3b01a01645f6253028c78a5fbe69cece4c5dc39a2d7d322078e49b5541844a7ed1cfd952917585bf86fe410c62eadb1d55694663ed92bfe51e0a3ad08fce9b2740626d2b3e930305bfb9cf0255aae22cc2e59e35c3397c880fb31efb69d63c4e38be938281c9dc5a51b1a6405a0fbbb9b9c80174ae2f12dd46bebb31faca0bf85ebdaa89e7e40a965c7a35a3577c7c499260ef153fe645bfee7cf2675a474e43f6a50847b63b81f348e792a2688ab25f11f7e10aa346e38c5a40c9762e1fc16661474693db372b1f515821208390ccdd208417480cec2c7433456a0755cb99eaee7ad7572e06e480e75941369f2f5cc0b0e5c03b662a103d2ebbe60fa6d053790e8cd78a1a30ab4621b64283e89675b3881eefc9f4b7ad6cc3ca5bde37630bd07d95a37ee134c3e483a3e78f47a2afb0b54fa9761a8b7987ac9f67fc4b6e193bd0008e52c4622e3a7a86680b831176b98a7b20f6e970201a21cb7f99d6899079739b8098109642c48eb4c4eb6aa8a040929e06c757f9918ee04c445969b769aa151088553010350de9de770c158650bb3a5bf6e932ceae72a6965b873b26317ec2b5a1c42c29ef5a541e63d0227c6f2009688f60f41e8b58ec1e7ad7725b0e6f084b98abb81797c08ad31f3a05aaf473a2ab25952d12fd8f836e222ff5be68479e80d60cd5cae85f196b577b398b62b5df0f24d1f936308e6c430606f916f8ae4a378956011b37883c6eaff089f9678d481c4de761dc592aa242be83e35ff333153e258ea32313179d5d317c327fb571f8f150c43aaeb440f934223727f32a2399067331f86f726d99d4d3a6d3a3646e8c0b5abda34a4afc5c52f0342e217c36855ffd4ae19acd36fa70782201fc1ecac6925a97fc139116b5e6b772712ccfd3a003f94e1758db02795860b94b907697ac21dd19a5274bd1782350888bae1ccd82a8e94e0ea3a3672f374de921f57ef57a38531ef01cb657826aa0853170f8043297d9df1eaaae1627967064a4cd594a8eb196ae0733b77b332234ee4980251aec3264c8946078ea3328bb3f5a358e4d70714cefe2bea2151d95f93115093c6d53ae1eb451796dac1376999e4d6e036586edb7e0c159fa116c48fbe31cce063b48ba162a4b9bd14bca1d6aa94f2bb5b;
        #1
        $finish();
    end
endmodule
