module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c9daba261107e3fe15aafe07b8d2266bf74cb5cd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1141531a1221f58c922e6da71cfba8d61105656aa56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3a677361c5d200fc53427963ebc6d0fb2e801365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a24c6410076ea5e2572bdc8e8980a21fc8dd35c25b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha75f4e4693db254684d2158ce39a043d2e4891407e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f0eded78b8253563afd161ab0d411f41e11cda8ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1834b8d6f496f31b03007f56c2b6bb2611e96ef2941;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3887f039f82cd46c780eb78190a55e6c425f81fd51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135ac5de337f822867fe9ae2558b0e8335de0968cd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1415daa507eb1a6787c125808ff13298742b4a27c01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40987a515119da9c317953f41a2ac9215cc989732f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62a115b97b366b16dde24289fc92eb1c13987aa667;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12cf7fa67c1bff8a6fb83deb45e4d5c803a6e44e04a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90111f4cc59209932499ca657d57977449d6bf614a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c73e07b4db08b4438d883224459f7cdd917e29dbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e438379f362098c08d5cfb5e1b5ab20d793b919f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6bda5f213b3a49503f3bb507beee76be2992435cb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1524c85fc6820292f86e8a9c7bd732b21e5621f81da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd00f26fbcf5a8b52037a277fda45a364a3c09ee9bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc650eef40082993e9291fc25fc77065ce18a780df8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11711457d07aa5687f315e3b4cdf6d83824276455a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126575237124d58edb9c0e3271bdf180aa149ffba27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd5860c188c96731dcd29f9ff9dcf27c9221abae76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c17a1e215dcfa70f5e636786f7148b301cbb3fc80a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dbc56ac77324327e62ce85882e813ba1c9b57dc3b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba0534bc71b2dd8b648541f02fb6a0377b4d83361b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1efb9e2c8bce4ed1718d9031b3e9047f57f914b0f59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6ba973afbb389dee64395bd5880442e5642d3728e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17932ddfd4c3db576f426b09e16abde1e99ec07152;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19891dc0326730ce275a759029e3474f672b6693daf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40f7b74e7f1c561cd883bfae5caeb088d23d90fc67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bdf96793f58fa0d09a54271df5b7b8f57fc48aae2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9cbf29327b7644485e288819da11c16b6ffff8189;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fddc3e81ab0250e7a07a441b645aa908cbcf68c3fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119b5cae1d6843e63635313270ea16851ac683cf350;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe451781bc11b817535c7832db3ca63b1ddf6ec6ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89435c3ddaad18416a0145856a42e7b292353c696;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3ebb2de7fc86246235a71dc36af48d0416434be87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63dcb286aedd324b04b8dbb387ae7df4d2eafe4796;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f44208797bb932b6b3bd9dc3e60ce2b4c5213d3ef3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164bbc34f4dc9206ed89e6172c3c84d6677f2f4f818;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c83ccc1609fa0c9f81f74630d400d41c476e993d67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4d1a594150a587572c5d23afb270630c7bfaf27e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he035c7f8bd268d848953af75bdaf78d5685fd955ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6837e9b1c52ebf83296928d3c3af1a610b61a6832;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha3ae3d42049aa1b3d4bdcb3f87749b038e4f0eb72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b557f24947885072c8aa8e9c18269f024700102ad2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15fbc6fb344b5e84cfa9cc78763e95d9774bf3aa6a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc60445b2df0c5dc962167f617ff62eabd21f877ddd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13436fcd17ed267b1f432ce98b722369d37dad4916c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c565395a69bf090923a3d1f1776d7de93d90d7d37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1483ef8381d87e7ef3b5450ed176bd593a0f71db456;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h546b20e68786cc36c506993b019c029aaac66a2e54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75a0c4bc19fc521dba497093b6d75e5fa821d2984d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bb98392ca06b8bd62cf8fa119ea6db14cd8447f84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0bdf096e4fda637eaf78428210e78aa6d36f85517;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ab81e1a8450220d56dc58679985eb709c03300083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd20be1fa5fb4e7c1dfe14b89878782199e4f353024;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff4ea8264bba6e9ab05b78bac5a799ebe010d260a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78cb342e229ba7293e173d2e3c4b6da6bc90d2329;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29cff3ff3804f20ede3d559e95108086fbdfca69a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1247e4f9a61f2a9a151b7ceebebdc6a7a583b211e25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54465291719f48415a6e31876ccce67568199065ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66014bca5f88e07b2d9df46de3251651b4685f9d61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h787d40af3199961b95d58eadf50927aee0399ff42a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e55f2afdf55548dde0d44c6ab64bf777c98d0b747;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1280feaef999d7efd3e99a64eccca3aa908e33a564b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4567bfb9e2c1759a7248dba70af734dd47cdf3a88b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h567df7399a07e08c9cd71f8d5c6e42e0a6e571940f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d7d62e4258adb7e0ba09daefc913c7df986169f1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10043a2d7e09c6b4c64bd3bb6df81594d1d23cee936;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b752cbcf2e4dac528bc9355018027d663238b9b24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e92a6dbb2e23a9cf0ecc90b7e5e35862f2f81bc77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e59a975b6a08397f0ddb9a1b7b9793e4ddc84e3e25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5394b28023d465f163d45b630ed84f103ac8c99828;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d5010cceea2464505d776cdb66f715c47f878481e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e99f85d118145755b2798b90d3a8c5a878aab90f5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b3b152837d767c1586d4006fcb61d0e7eedaaadee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfa2263e5a00afeed7e43d55b21dd091bc19d74bec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd267645d20f41161e3bde9df9dab4ecd359e63de40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a17181e6c6fc901aff354592cd59cbda87a8cb04b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb02d749531027f7a8e968e4b1dffa880359c7b7da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6d9e2568bf739e5b61bfeb290ec50da10d46cbc10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf366037f7207ba3b91df6ae308f984730b9b05624a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f39120a6f46471b1caaf42bb24f3c6d56b840b022;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22be205e3408b1601ed48d516ba42fe8dfd7ef0ddc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f38cd34129164e3f85dffba5e7a835a31dec784fa6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha592cef88bccc0f1f7590da27cb975b08dc155a231;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a92657c03e5731b8ae2d39b8ff279b184e764581a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed41a0ce5c2eef4b4b69b448321cf635eac3e96149;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ccc0ba92705489ece1143fea94247baf22af2f120;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h817bb53589f8af8faab7965046fcdebe3a6da34f2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d2f23f49fe43fd5dd36fe65c67d3f014afe345d92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1552dffdaae8054750dad8f5c28f9e6cd89063ba6cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a5a804a5b8fc465567f795b3539de0de49da3b614;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12cb9f15b733f3897393020719d22d14254f15d6975;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3afd3d0332737a2719e35a2a833b81c456eb1230c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7364e390ff9c81c15ba56e15b7e784fb74b71f42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66087d7ba5b11dce56883c4a30149aa7a3bb526a61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ecd7d3c772c4f3e1f0b1d485a904c500ae7d7da22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a73590028067d9f71c98cc41f7c22d56692162824;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82bec1e15c10e667953726f2cb6b480552fd48a34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86c741b0eec137061b918d45612e588f3ef8a7884;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34a6a30f0e46d90c45b3460bed02ab60598a006a01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ac0d0ea46e2a32357532fb081f3a2ce1342e1734c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131c2fc86c81de571cb0fd41dcfceb55af4b8cbcd8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h540a544f8d2ac4ef671a7e662b333c98780523ce3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4228fcae96d3ded7a09d2c7f1ff24c44f8b91be9b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7949d8ef533c839c414793362926dad979f85b2d65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h463bdba768da7a09aa1a00c84b9104cb7dd6a66634;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df42ed099fb2b094c99af81cc7f4d690e4db65fff5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba6f39395024f167fed8b3b15d6ecd23c49740dc50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee882ef84513e71b092bd100ff33cfb225f3a05dfc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4bfa030f873aa00a39f54d3c115868ffc714007d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58f32613402a4e502a45a768e0f1fb689eb2dddb47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32c17af4db2a3439a75c057453c651a7932331a350;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbe8468dcbf25e72347c980f6a607de4ace39567c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178b844a5434c8a7e60e3acf11c7f2cbe4f57e68acf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75c0adec94db513977b7fe347a0a88253d9661fd78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb8902b8b128a026456af24d8c6cdd4eef458225b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175a4ef44d799ef1a07fa720e97c401ef0fc715786a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58711abe215f9c52e73f2fe20a02ee4502378d0429;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8436d636e370352de362d758d73cc7fec4f7a0dda6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d7fef4bb3e11f68d5a0c84e295f6805c345979cb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194712096479755a627fa6698c833b4689b5afe5981;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe72812d8268a7b18df66c4a12cc79603dce97ff6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f1a5c6f13fc321d39bea901aa8e339a7971dc5fe3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87709750c72ddc15570e999627b5ee9ca912958c01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h400e1c289f855ca1a9d0ed0b349aa872480ac0171a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb92ea8c759c74c5f67a2c18374ca09c7f1c35f500b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5e514c7d78b38442de23c505ba2f7e63acd33857c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195780a26734232a2ebe674c20a68bc272f64f05ba8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2aa7adbad0b75224eab873403c5263bf68bd7b44c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175850d9966b17b9cbb617be76d3614979d70e10f08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf8e11de460a2a6457dda27575d13b9d8f57cb8fe6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ce4749105af5f9ccfa6f2a80489dda97f9d9a5e49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9b7d9c44d25449c0efd9b7358ac3dbe9b78f3f9a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c1e240bdd424ad373fc273a4816c6623ce998b491;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8e8bc432bd875fd63dbdcd0f020b1a54a932592f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ccbdd33eba0df8ae74a2cc84704a45cadd58483b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154e582202b03acaeacab816773558bdbd2365e9adf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63229dcf19dfcfdd37db4290af22163f831c0eb3e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1948ae2b8bb7073930f19876395721425ff0da6e9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d6c4f6da70b55b9a000c065819b4c62bd3e77d413;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81f4c9b7c1a0d1e7e98b56008b0b888854ebf7fd1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b7cd3f0307e6947c3e8364ade40440d206b596575f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ac314c7d8757eceaf803aca8571f8e0d6a14d6878;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15bed3ae7b51f549949ea7791b695d21dd80b847051;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1faf9f3195c9983afea7632300650551bedabd52407;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1746545f342957251a4fec576344bed19e962be703d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a910a34f4b40d793455d187b37b41683a2d7336be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148c8d2ee7745beac25b66d46594db67a0cb00cbccd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d47e29f6eb8d3e98d2dc66434f9174b78b6de989c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h780f5bf723e739e367135cb359f3e9de93fec7e232;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h869b3bf7f4fd7ca76cf39d4e3e65b3affb44f14e38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6585716fa7acf859a1c228523cf7b49393d1c04c0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbac9c7f55ef4470816424d8f68b1674d983015e09c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e75917831acace4a7653812fc03a3c9bdb26ca52a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100295af831a806c274fe1aba977cc8d0c07c9fce0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1804553940ab3919e61a20d4c04b09288d4261548e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fafa757f81cba773bfc824b0ecdd6438fb80a13643;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21c088eb34027217e8ec9bbfee4b96975511dd596e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb42d2e97603e5e69983d4c53af12fc86bab8cd2c26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb665109325a2b24bbdd05bb424acf530b73790147;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62544cb74692056ec47fa8b2a4638aa9c3144880a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdaabfaac03000b1cc790d4fbb4e318b94041ce60c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ff85f274631b45ab90e591d03537d178c5cfd9e14;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a5c423b130c42c06ddd99ac8b795c5b7a09ed5fd1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f243940918bc00e3c4b84b5883ae0d746cb0d4c096;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h139dccf7e69033d19ccb024a6c2fbc5795ee91c5946;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f42fdfbc5452835774acb7e57e32716d0d43646cef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h850888aedeca26f873175df6afbd46366207f2aa09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e52e666621495527c4b3a65da1af1fe178d6857e5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c472211c5b96bbe55b95c4768333b532e5291c1b55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9cbfcbdfea81cb257f53b7309c26647cf41056c2a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfba06958fef64108c2f49c84f46e6e1aa257e10b6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd91aa1fa3c30571b2be2021e5711125126a3254288;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a8c03eb0e9a1f51cdf9eaa74cf4f5de3c3e5987372;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147099e7a1183f2b00d60b694ab611e6d5be755682;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132b2224f0008ecf5c283413963b2b0b85847f33054;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf51cf695aa84376165b62dbfe1b8a07d5c8aa971c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8467b66b890a119895abbf8896a533c68300de27b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b11ac09006853adcf5873e64bb11f0882251952211;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he43dc45174908d5ca1887985b5f1eabf64a2ed5979;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e0896742a700b7b49023fd4ec8d295350497fdded;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h276d80622295d867fab1e20c2695bbe372304b9e55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1335aa693699fca172c415c97dcd2688092280cc072;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123d4b62fe070eaf039951f67e8e99562e033ce93e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c245bbf41a9a616cbc4e99cb5f8993429c87f5dcb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb424f390a2a804351ab9cace68ea679e4d9c1ec1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b4efb03f914b7e5f25038f46b3baa76fd46152b2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f0b330c6d177b938012ec6eec1c2446a3939485b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f4c08db330b0d080c561ead1188a165c2ae835f04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c77ffd7a35fe14a96a523fdef508f44b3f7ae3048;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4dcde35f090b6ad9636a39e24e1f3ac86ea6955f6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16705445df1dcc78a6d825156c123b555d94f6ebaaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19bbad7ddc5006fb1ce86563136c5ac4a440fa6dbed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111cd286bc0a22eb0e43d2156b600d533042a7ba875;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc6d79f56eaeaa5b52bf98b463011dce9def36349c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157861058129b2b885d25512344d24f9ed2d92236a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4071670f7866dcb467211f4336e83a29423f1695b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c00b61e30912d88924b9a6ad5d49841562b71b10d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d95cf498b75c3205467df9964c7b131e67528dc027;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11355807f3f6fecede98684d599b46dd93601538a46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha96134116a2ccf10d7cc4277f1af2ece6dcffcfe53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h305b0a9954d807c48ee970435235139d8142d669fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ecbc6bf751c32a0890af3ec4e6e76fb749e30e524;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f9e13cdd3ecde9eff6b73b70bd422762ba281376f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119cc10a5141479a1f6b5fc61d5a27e693902c951eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a203ccdfe0a2d0cb09222aa3d45640d877b7ecfd66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1063740dfc76769a016b04bf180ea7396109ebe614b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e5fe936802c5b57a0956c0bc9912a84b8296d7fe3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb88727b4a95bf24e0a711c1f1bfa40c8dd19a7a02a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6227e91fab04cba04e365e99596fc4dc8b9bc565ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a9691830669c7c98c8117f241c35146aaf997f95e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5953ffcc65700fe18f09e7d00aaf3ea378df488fed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b150bd4f4de3d913f83b3fef25aef1c1312d1b2f78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14bb7e071b22280763e3e30b95bf1d300b2debba750;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5ac931fa785b6b5084f92f1306e053a1f0729e7f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169621374d750b485a5e6349e9564d909a1fa577733;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a831d6b284d9eed68ae5b411514699ca136b36d64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d94b08ca693895453f8d1ebb04a7d9bb8dca7058c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d58c53dd279f8e8799fa92019f4d470dcb93cbde45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122881fac21b67d51163acec5ce64455c0101910a09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9470847835f3d9efa853a5c6670df3dd1c088c721;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b1914ae0fe27967de08a71f739c5630ade1aa53cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1b035dbfa446cddfbbf67e3fa9545ac3ce584297;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110dd463424b930fc4ee5262aa0838fd29d41572e0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb285e400c644c010293f62c2d789a1ab975cfc72d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb689f5627d3ebbaecc91b6da54026b9ca4f619376f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45488a81548428ee113d3cb3ff3ee06643d32e1b53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc1da958bf3065c8c9684f37ee1c0d9ce12c6e6c5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165b12b7398f1a322caff8e715c358acae29f3f65c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f1027fe1678223200c23f683f84b7f29721281809;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ceb884d6a308621baae48b671047ad88adbf870a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c7eb576c57290fac98b21c29d9ad340ae8ffd65bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4fab22a22999afd779a3d7e8ca8dae2974876a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d053cbc0504c7e353027d462b519dc41905b9ec129;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1336a7da08d43111aea495eb2ea7a5f12bf23406d2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1bd5f0e3a6ebd3cc0bab46dcdede456cee933d184;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h212b8351bde4f79d573549a6ce0d3ce9d6dfaab46c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198c2b50f7edbf1c03809a6f97b852ede25ef6eb0ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1535ba0ddcaefabba9abbbd1e3f713b6e1cbce4bff0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87cb3dd7b6c0f4c746935a5a0abcb1fe16324114f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130de18c62b771c95a17b8a71823edbd11eb4066b44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc9d4af9928f6043421215c8ba82f3f52a255e286b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h816bd7c569747fa607d2d544e205e6268bcfab7c39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3dc83240d62edd2866aedd2627092319cffe2662a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187950393ed1a305a59ad985424989ba088486dacf1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bdad3595245c170b6bb664401688e2737aca1c362;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd24c242f277b0c6759d33b62994842c8e010f8296;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb67163951bf796cf85197e56df72acd4664835902;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140bc128224c70063b457fd96094ac73667d3f99901;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17faa87ecd2caff46b697f735a78a63bc494b03da6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7f0e3303343e0ebdf69c5fa2ad669131c137e73ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db5a41209c7bd474a348a32c6319a52e063af02adc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6dad3764a64831d568124a937322eb0b691e7893d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fda707f6976713a019aa3b126548fb5fe07833b4d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a48eb687e1a5bf9aecf06e7e11bd87ecfe3605bae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5e1333198b984aa4b248762258ebec8e395e51e78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73c4eadc9853ac4eba8db8c0b274ef8d33c4a2b61d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fcb4fc20fc272e0a7c204906e6e54cda0057f2174;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e4cf8ace525d8b69ead421228dfc5e20ac207a3c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e65440cdd7a2179eaa319db811f090c30b6e2012e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a644d4371b76cdedeb3f890e8f05272574da9190c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h799026c71fd04cbcd737dfc62e76f264c6afc6c504;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1662f82a7ab675b4564dee5554f5f08187b4c225aa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87eca8e96df5939f3bf54ce87342fafd2d3103479f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d6d19aee551913f218e4405fc93d6360010c53b51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57b780ba5d6c6bca59064d7c31c6e031fe276c2072;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b027993bac28173c6cfd023279edfbd873bac26b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f331bbcc934e56cece77f69136c72585ee2f3946f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162faa23dbbdd2eadb78b2f2cfa2a7f91a69c9bd962;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc09f8148454b60a2690e94390cefe2cfc0db147380;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf38251e3a5603235da7dd8cb2444f4e2c1320c172d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6f8a4d6e2f4319ea06df3cb202408605dd9c99f13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae301fc25cd6388d25ec40f18a46c0a2db112909d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17084eb4c7754f4c2e42a2c20ee6a2970dddf511af9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd8c71baf3f83c15baef514c3e44a34e11e8863a9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b3dcfb978e9fd2f0294b8405ea6c851f759610977;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11c36552e9bee830af6b8e21694912c0b0210e80d42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfcf11263e995ae402eb4f2c26a8b91ffd5cfbbe83d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea5a797c881be1da872c3c977f32dc952ca8a503b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e17f0185033d6d8db23f1098669b706949392d2f97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54e2255f8cbcfa72894ab56e3594d560205190a3b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9195e442d849c47503ad2547208ab1d2f162fb64e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1837ad657ae3757b3ed3276814cca441d3e8919f2fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f361db811b9e9530fe411f3a6720177baeaf1b2ffe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha29ee4ecad284f70c1eb19469e29926307d452d43f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ae4ec6b98a9dad21df38478224bdd5dedb82d0b58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c0e720d8396e6b496bedfb94f216b4d2fb81095ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd76867cd391501183362df48298995c014658c7124;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19956210ed0fbb4a9105619398f3ae94d3241ab49fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8c8eea1662162d31e45fdfa4ac99ab61039ad79ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h191571622def1a48b97df512d548f9c9b399fe57e29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1790bf2abed7e426c5d1da2b353e1a9a0bceb84631b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142074874bc1353eea1c264bbace42ca7cb4d24d985;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c6804aca8dd4911db9ec80b461e54d989886e0b12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4636979e2d467f09825b114e9be9b6cd194d7302cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h539f2db3213f97feefa0e3fe4003e5f84b9caf18b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb09dc2b2d17ebbaa16e4c2229332d9cc6492a4783;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2833d94850d9da9b473f7cdbc16432a859c697c723;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae5b630495e3be7d09b00e0a4d84fae7a3bf2e7e12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3be98206012d11a798816f49d64a16d266f643df6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1613cf5c4df3a0af0df2b283f36b04395c28450a8a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165b57a49e8b8503672424d8463eca85ac67651bb3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c8f475b0a75f826081071a60e4560a3e68c42128e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d27c26a7088e96d4b2be6fc61aad5d9d058ae9806;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3e08448e214497af7fea1abdea40b067b54f0bffd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1592358cbc6ff49a50a5da60a0897bc8f36a18f6ed9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha45f4ab72160182cf6bfc9901ad1268ba7aff61876;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a99ac20d9710f2182d043909c0ee416866dd8524a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf680b8d7f1907ecf36116c52dc2563d57709aae41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ea363c1c3f1b0afdfb2c959266642d49895749e8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc4e5cf6da303b9ec1398ae6dab085be156ba6ae50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bad226c077ffc06e07a85286930bd32f6c92d59f29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39cbea7df9f63b3543f036f1e6dfc77b7fe407b196;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8863511d15abed902822284208faf7e52d02781b5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12616b3911fbe05a7f510324568bae0bfb6d745f2e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb78031d7783b80bdbab23f301f96c15451bafd527;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdae0e856eb840b8bf40ac2e12686281d0a56ff97da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcea9069339ac2228523edb4852332c9653adeb647d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14197159a07ec52bf55ba0e4a6b5a2a1f2649ede5f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb5b3c8e73640070ba7200486fd074947011df058c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdabd35c7132e55c34e06f84ab693702d969b7ee0f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101103f01079ae56309dc2e9500f113501ac0f7b33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haedb9f25e64216ae31f8757b2c58f6eeb4422cfe86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1923deaf231d97e33aa1c494e744b92e0393cc70a4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93f25027a35e3ba0d04a9942f81590898fecaf6f7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142eed95fc32339542de58b8efc06114aee86ff4353;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e2cc2d5d1ba085686dbb272af5294c68749e2721a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha3d00fbdf0c1057edd57f39b3d60ef630c7f40dc0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e2e07618f4907ecd169228807f8f5ba99823815c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2960d70eabe4dfb13b5794d97a1ce83d3d5a5f370;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123c1addef3347f8fdcd4c44226fc52ee8bb21af5ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12eec1431201cefbda2892378a8651dbf4e697366b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fa7e3c3450180a405a235c5b59a140ba626f8dbff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b5537a80b70ae97a74c8011831174065e185342c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had3e8bcf63ba25d1c2e6769dae3d3d7e8d3694d4af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c15d86f4a1866deba627f389bb71546b5886ce49b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefe18ca6bc9647d4c50485e5294a6178002f22ec3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d0b8883d88b3165170955cca5d91178f0caa4cb25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14be450e3e28da00ec402a40c4ffcbbd7286acaa713;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d641b711cd0ced5fbc01f14c7e03ba1b444037f880;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8e1991844aaeb202a1ca28fd954e08c7c60a3e6fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5766cf510afadc0b8db2ce4c8b3a916259e70a94e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15981c8e512f0bbee2551a855ba0a114889e81d0e0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he13502b61f92662365b4fc34ad25143304ce101f6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173392cc03708c65dbcd1e8c1b0998939f3131fadc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3758a43fce27988d86ebe53de1036b3eaf278f370b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6690c96d9680b657e3f71599febd0f413313c14a31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h276c8c2a02ca645da9045d1188327b519f9657668d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69d1a12aeda703ad16f435dcdbf0ca9d8f9f8ab939;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161713f67ca466adf030efe03f6bf96df1b7a117c0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5346f6273f63e3097fe8867656c2f0ac90c15a35a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed8d7569314c12b6ed60a0687e6e830549569db63e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101f5bda8218f90d69a7b0cdf2156b6a5b9561c6aa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd0def76d8c4a85bc2df673ed8e08122a5a399e69e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e34b228be9c11312fcf54986dc0e7c07e3adb6a0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72b969565d78714656c5830d4887c9ce4856d92d27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141ce72091e7fa196066cde5030df3f7068764d106e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f85c11408a9d59c16984443500df3eb259a84fb153;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3fbf21e9da8d184a84459502315811123054995c50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185c496f511c358eb79b32c9a04b9968f392175f65d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8f00c23894b14633ceccf1a5f4dd7ae6dcb9ae9aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f13c6e399c53eca247623a540b8269b6d36cc0e16e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9ff0c1cbc2df86c052a5ac826b03aac67526385fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haec291c4af5884785005fe8e97bb2d8054952bd03f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13065d7c10331418385de29b43026749614e5f04e8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11226c6f400e757b593fed880a4652b4b16a14c5fce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d956a93bb1e72543f410af4f0a06ce8433a66134d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197501341fef9686932ef92a980fcfe95938e8e3b20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc57760078948de22de33c889e5b60ac45baf2e3c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d02cd807e3c8b1560ed719d336e77a5d8c1fb5109e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f63f604e6c957fe3217948fb30802062bd2d9246ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h411a30b6c3f3e87df27dd3ce9caf7b93f4009c77f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12096d8edd0e2de87b8c6330dbecf74cd8c685263ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd86af78ba3e8a6f34ae7524897681d0767cfe2140;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9292d114a5d01a0fa7abf52d8d9f4e13ae02b1fedc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fd5c748a3dc1bfc761eded64c97f91eda7a4ad663;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75e36953b18fffdc9d1a9e1a699ee64ec5b5c57b41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12833dadc884dbfd366d8a7495199b0a196b1815074;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcb699d9b34fb03332b42af2c227b157986d77d984;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128d33b2cc843c80186106de29d6a32d4b0711db825;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha54165769542cfceceb51fdf6af912887ab3e7253a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183185e4075ef54ffc4988be977842d967537566037;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3a7053871fbff5645f594a4d7e741df14f5e5e1f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc965b6791d12b0e4e0e36a1e4532143fa0d922f4a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113158f1fe5cf43716141f5ac4eafa544f78b5149ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3cc9656cad60505b1094b9062eecd6e41d3fe97ec2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180986bd44c619df0480f4d3b9aa34993af393da77c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee4bf7eebb1e433a5cc459b66f54e5d8c931e39873;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c37dd7c8e6fe3d1ff4513ed83cb6ab791e507f9cb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a620e99141fe572ee401c04392226c618e3bb169cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1865e5035841ae89885f9aaa3bcbe6e2dde8c2bb0b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5743c1987b541dfcba627fc1e733a6a59aa5502fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142a39a977c93f3c88d9fc2ee56d9ccfb7814e2d755;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdfb89ddbf47e6d5795582f739a6873114e8351045;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114fada3cbff2b4a7e6e58f4964b4594f011f8773b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3d80dfb0447d410a5aaf49a286160e340c98516ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d536697660dfe1c2f7b7a7d740d80840f21c25b1ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f354d7cb3184148df2708037c085251437ec97664;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdea82e2020c4c4cdedcc9438bb24603cf88676297;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h317f7303117d249f89970c90f3547128e4ceb0b22b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b5ce921bab513f617053d149171c0c1e654adcfce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5eb05b5751bfecace07a2b46a133e4c507b9c1c45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2658b4215539c337dff7ce1f7b97e2db71b09d29b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4d9c0cb3abdd527305af2a6fb6d06af00f99bcbf4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118aee0660b8aa3794a56e09cf8a6974e0d2b9617b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19253d8ff2e9d7b1e819a7130d837032972b3d9e752;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he29f979e4f721573fe5ef24db1bb77df4eafade1fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c0de366c3dbeee333f7f09d3957869e891eabcb87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e782a05bf31218eb4d4a72da8bc9c81d101101869;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b3b9e6fc03d669d57591890c3e6b666eeff9e1cc5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff3caf1706414ce1b2e8d8d67404f602a2d019cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d66f0b2cdaaea969f4e2d981672bafb52571ba1ad6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78c73f62eab1b8150c7f81db8851dd7325e12ae1bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12efab28d50fe36995ea838b621451c6bb1e500026a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5a77d78ccbc0013ab986aeb00d2759c6baf05aeb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e5010c8dfea0e9d0bc08eb424d60c0c8154a8aa5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138c534fd4cc63221f71b5dee263ac6be0844dde8e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1358bcb6ca495ba6fed80d607db75532e0e736c30d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5801f474234d08dbd30f11d6b2a5e49c345a3d1962;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcdc376f602a43dba7dde627fe059947dc69266b87a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e8e2739f75383906ac0d065e90d48416148bf2c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e243cb9dc527febe188bf2098d24b86168ad039e92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa240aecdd563ac689dcc7c1af1f3d40b4087dc483;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcbf06cc3c8f61d94261a490a1dfdbb17f40a2f75a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fca65d8ac05b2ae089b0c426237e13453d68bd2222;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a60e0f6c591997aca96433ac3c99ab8056c9463e3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bdd664f10343dc2ddd295eb431af8adf0000e086c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e27b8a2d2389e2dc06a63ee233ea357e1d026845f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h790335341782b918f301e02ef17a4073e4c8acf6c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c40df370e316a0733921ee672220efb2cf5a706e14;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1f4c148319b8f1e73baebff4232bab44e3291551b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h828b3a097df923d323b44a8b6de0a88b96ed074e63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148276be208af38bd4fbf53f5320ce50c76879863e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4908edf34e9c837c30323ac083aef5f943e02df78e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1abfe833bc142d194a54d703427d3f162380d3d851a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4bd808cf01da2f627a17201166842f01f297b5b2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9380cfd48743f457db741bc977e3a63772f669eee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h273322b840fb50f2e407ed4c4f7e6f3d6ac23f554a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125a1461ee5fe9ca5013d8e81bafefb7822c39f0395;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eae9c50a1c5f0d9ba60c3ca316e8e631ce9dfdcfa1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103a7ba6b9c04cbe94cb597c7b83f518ce7788335d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4555c79c21323d723ae7ce318d88ef96a733791cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193e22342e11d35a307cc3fb3b5ff10c853ad1061fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e59d789a42657edf1718c5feb9090ffb669c2675d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81e473bad58b6252fc386c02b7bde7ad6038d25bd7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ce64beba4f5aa44c698d172714c994629e2affd43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca82ac4c3638ccc3980a3630d639217606d9c5000c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13cca74a20c553c99fe54bccd2a393beec7f8fdc341;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b6b90ea45639c0a691ddc36fc3e0b4854207eb5ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ed039e309a0f9fb66d8d1511417a92b3a0575f396;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ec3338ea6e8925788a11f7a904d9bd80d1d751bc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15aa3f92ebd6464b04aa16419f6464593ef3e6c76c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e82fa2eec7dcbd6c33c7b102661264440b6c322d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e957c1a9058fc4b90c389387b6a1e2deea76b622c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d60ed3da1a8c921f92c0bf6449c3d00f265edbca0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61f4a545789a486e99d750f4cf3535b62ccd0291bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1552ffc70bce5fcad10ac7ca15b3d9f2fcab2539cb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1125417f4969d9018ba280058e0d7b2ec15488324;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168fe4a911250b5ad593493e88641c58994a8fcdd0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a6e98015dcfcb698637be54fb9e6e9322af9a2e8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1557419a2ee33d929dbcc924114fd990eda8d921465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b3eee6c6746caa8ba35b878e7d6de80afba8c4e1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3194f9c5409643a227c6b5f95a3a7e69057508030;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6a9eec98990c663f0c654f89a2b1a562a62781f2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1effd17d58a110eebf9622f95f68a59fb65f309a1ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b8fd21d11034e1318909a5d8c0f01024a1d0183b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d8bbbee48c466d63b93191d25a57de5ba0590b115;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35477cc1352bbd4ce11cec77ffe1dfa4fba38dd286;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1584779ab46494402e59abd6f0e540939d632041ccb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b02a8a3538a8e00703023438ab5ef520e9c7a376;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee3d3d055edb6a0a321b69d78875170ec3edf9401a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf22f3d50c2ffe26f209ef4f56ba984f38cc8397bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a8a6df4a33cfb2e5c5e9f095cd2880ac142220a06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fb6367f684485c656b4e10e8539f99336d22edaff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dca34dea3ce0942db281ff66847f3b0c8a56e568e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5227d61ca0703ac7406b95d261fdc20f39d01d311;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110e8e61f6658370e8504d9be44c43490b200b01e4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b451028e9ff44fd3645655cdeb26b19b9da7a30e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10564388dfb7ecd4ccba3db292418174099d3163f69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142bfc6c4d0340fba09d17f1f48f404125a63f7e671;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd198292a688dd076e21b1fcc848e86935d0d7f4524;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4b67c565aa9ec5dd6a2ed02a6f19a4fb77ed28276;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd08ad2e7ccd5972d1d01811006f96a5cd70ee1dd1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf963f359690701c989d7b74ddbb5a80ae9aee851d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1157fa24f0367e0ee042dc593de5f2dc628f9fc3ed7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b175e9d8d59410b981a88ca92027842dd645be207;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c124a914d28dc67265d90cfe35f1d289f2abe513ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h780fc76d1feea663683f473d5d687269c7a77d9a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h105f7a07c06db30ca50d253c1fa136ac0a793b99b62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6faed12738f1d1d66aeb0edb62e28df7c4bf959d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fdb76f3546db5a9e458aadd6fde0315d04d49e8ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8939c463d6341b1373fde5fbe084b40a6f2206d829;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f1328c2750a9357498c66c7672e62eb11a72c8c9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8c646980a96da6a4802de4ff28a1db13ff78bbd53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42aec6c356052fcca1889391d7028d9faff3c4581b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b10f714ab69c5b8db6cc87936eaf6d69d0ff27a14a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b800402da22ef1bc9e2f958c32728d0fde05240a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128223e012b61c41c223bce490b97c2473e3dced288;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1594ee0209456a9b2551a8ce4eee2be5cfe4ff24284;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1148845b484960573078833caa732b790aa485abad3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1334adc9c7927337ad6485473b910eda5a403ed173f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164c2457d5e075f63445f8dd69c990e26bd54d03c66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7719ea4245fe1c662c4fbdad60b0ed0e53a9fa09a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194da18b35f7f4d10d7132c0a09827654406ff5330e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde5b0690d35cb3ec4dae3d3860ad701a717fb0c4e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a6b150dcf2fc91ec0f2aceb867f2abb575cfa081d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5376cc227c3b4cf4d8e5d6fdb7d358e405c28e1b09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36504d04b3e6ccaa7d18b821f2642698794d99c803;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h96bd3922162f1b598152434094bce019ca7473d725;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15946ee7a54a9cf8061452345c917892f3569f9d6fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c101df52eea3faa904a8c27608bfdf42211c1f276;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1935e9f615474f92087a9a507c7466366b27ebd8acd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hacbd34144ef7bbac562965d1c1e8617ac701ee0213;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15677ffbaec5bfc9b029a23d52821f29831b2d25840;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9daf8933612ff9bd2394d506375652fe82871985f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27fb3789a08866298ba6383283ccc0336d06fc07b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7ff822ce6ff7313cfab555705db4439e13ba912b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1852630a4f6a9d314219de5266fa25a1ad5fd984c41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f5e7a21da4d8ab419f14c7188d29b67f3cacd1e8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1228d9c9776252d383f6c7be7fb3ca5d20d3d6985cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4804eb8c213579542f2368e91a6344d9c7e7dd2ef8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19fe4e4dc6bdca01d3245ac0f81d4bb4b76cfb8b13a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124b3f14544a36b02069b0f595eeca4a54eb662d742;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c48a68dcc6f1602ce0e71213b99a4a4e1fce3d014;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heeda3335598624a7c7f2518b2bea1eb09417a4b8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4bd0f2fa7a46e26e69cf49e04ec1cf61237864396;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51ddeefaa6e7250497a3ebf43ff8247321b732741e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77b1eb4cd85ff753de87eb531097e913cdfa04f93b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf4167b3e7972549f0da5e87da507c3bee9c5034cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1987be8ca5f71585d5c8db2f5dc351869f9c63fd83a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d17d9e3826d440666b1d7cfec987b0d70f3d135465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb3f70afe48334a0c5d9c6a2fd8fe80473550d69bc9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b8593dafdb3cc607d02c5f1cf8ad1d3c14ea091b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1299e1bf338470e5141f961e67dc86dffb4639e60ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1223faca75434fd1afac6203a4ba6d15538502904;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1acacc176c4539bb5b66788427baf599945eb9fd0ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e1e334dc478a70bb65882d0fb2fd23b60936330d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a9004acda119ac26024c6653e200df27419f854cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff18611030edee4034922a96d98072eb5cdbed990b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190a20ca9e43e9b1d4bacd8f6cffd90aa5b8db80c7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5bc16e256d197be2b16aef1c85d863e9a2faf5a776;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbae9b304bc261e9872f2fb6115298c82a24fd79c5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a1e4329303ef1f0b8cbe0a72538b0319e59f016ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1893947b2357fdc31bb3332ac5cd3f60927a19cadf7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a61fa879cf93985fbcf44d5c176338ad5771347e9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d2fb07bd3119b449420acce4be3db0f98cf8b8abf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117d65c64b85fd09d1fdb8f06818ab67e0f6284a611;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15603eb486d132fa789cfddfd1f9fb241df481afa63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cce92d37238bfe490fad17684949867d40c82c8762;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bca5784823fad6bd4bd3b9bef1be1761606c28ec66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe389be8958018a9762d7748f1fc641b50617b677;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb3f6d7c2fc18017c2a20d5905022ab0113ab6dd36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba21f53c3c1a892be4baa4fa511a3e4e83dc548782;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd81caea7121bdc76d9a840fd9e49a43c691185e98e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12de1db3c7e22fdcc2f2b643a6e30930405c5bc4b9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ea3a3ba4a3ace85a1f865cd0f1fbe73944f1510b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb11fac6acbd5396d799d8196e39cce8f9b947d942c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b0460ff20322e175872587fdc75d4d5ae643ebc902;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa2cfb7164083e590429fa028fca94b8393b170401;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14358388ed3391819aa43ad411227f6f9d4dc42e09f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36d9935b65dc833019bfdb4602e9f573508b26ab5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde4ae980ca95bce4257f9bbe5ee4077a00edec7c03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e9d500707f16f3924efed303098e138c80f0e655;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f29f7f73f93f43f20ad86d7b11c9358e3a3883364;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1adb229c1b42f6008bc674e131c2f6e365a32ead9c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5d4e0977f48a5bb42d70b2ca2cbd8baa9ae7f8e75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf03ae99e049d533e616515be147099fdfb618f4e19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf445a6119d212b895fceea42a435509d4d9164f6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0f7beadda9c849b2a1e216e10fb224b038735bdda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3a6deb98bde5d8dce3bfe3b2dc67c5d3294b9d3e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1183e9ae05f2bc301c8ac479e854dee23c7dd526b8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e0a98cb996dcf687fefd8fad78cd0136398dbde55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55c4a0772d2c8701a389b91fe4545be24f0cf9e90e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf1976b602415fe6728950f93a0c3008404b5b62aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb92a8e2861f8fad56a9b0b90a45371e940ed8de37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he27a433dc2300a85a0ea95097d779d708f62fb039c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bce870f2ba9970d274d4f999ddecc59cb94f633a1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h346d6fe2926321fe1dabe95f87502209f40251ee82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80a24064a64bf3e859ca5b961a7d4636d170f3ee07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11b701ba57459b41a943ea0ff21268419f0d7947bb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1904232bcacae57a460d2a00d3bda245d78b7a37fc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6e037c1b7dd8996bcfdfee05377fd4365d190ccb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0293f4ef8c9cb7f2f1d1dc2ce066bf5c431132f45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b24c45fadb5230fad086388101b13f0408a4ddc38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfda56505dce69d8d9393fd58eccaf07fe4b664ebd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a93dec523431d174b760f4d07ba6e586c17c68961c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147bb4b4feeefdb96b7db4ead0f7c0c142b5402dbb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11887b3ae52c59a257aa9c6365629c18101de29804a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c997125e8277b4284b3ab64a8f732f68ec01e0a969;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e3e9b1017c9f7048b180180b262fe5c770cb3951a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11714a9d60ffddb1b08ba9cd10b4f204350e707e09d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d24ea1b95d6e29e7f1ed49f0e9b895f90217d461d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ec2479b0f096f7669048c5bbf8970c074c9edf26d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h564edd8bc90925bf19e3d763bbc6e449e19601d01f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7cf0e499c1791ac4b7f2eead0ad006768987c14a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h858b114878c15e2b9fcbe2d47582110ceda2ebf49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1404d1435ba932737e29dba05a95551dbf0b719c406;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72b1d933467b735d1485b3e95a888773c98556ee77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a09ed95b8ac9a5ec0d6c00df5b577eea85d92649dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92e795f8a30e17d0eeedf789060cc2395ec5a25260;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h218c49c020f0dfd194279d3442a5c77621f80e07cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h362dd182053035543cb7f60d027985cb701a7f9295;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd864469b6c3902129798e0b36d6818d1628913996d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h37239e7276c7936713fc9f8ff5f6469abbb39e102c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef0a7ccd64e2c079f0f20013d80317e97e20c321a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a5c6f2c12bd4f0bbd226ad7bcfe2e0cecb48180e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118b0f114fa4ee03fb333c6ff1fdefeb34facf4f34a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44571912e81050b68e4760ee233d9e306077a96a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1823bb9482c38e3870596aad08364db4f5c3e5c903f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd6eaa882ed445cb9e1b2efbce0e54d62159e1464d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7e5807fa40f14a6a0be6d8f0725701a823fe7b557;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175fddebeb1eaa17c8a8dbde4c5992b32b840b0fd70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182f5d4adb934072cb93ad7731f488d197b11194d00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb6616f331d75d2d36929487ddf4403dc96f59ec1f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10126c017bad54d32668a2da6d3d5caec13d34ab472;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124f8c212cd6a2d0f3b478c36e8234f156c59169d4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc5aa6c6615e617f3f3cca5a009b92ecaef34fa3da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd22e40d4ae0fdadaf2e70e94421d2fbee6f5bcbf87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166e4cdefe6bfcf923f74483e6991b9d9a7f6bcc737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78306c70980539539c0b59833857a82ce957e3eaa0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9570ab6ef3df4bee4de5f3eff3c7a263b94dd0efe4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d2e259685786f79b9feab17eeb3c9cb06b1494298;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb37d343d07758213b4517805e5c45fab97b16e6709;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22706951716532b212bbc0363b9c699655402b1c7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h280c360fd7c3da016fea013b44a00ad33c0cc3aa2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193a8154d7dc9b7651407b48f0558d0df8e7e507f88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1896973729b1d1396c90f8f4e217bb4ea00222dc9dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he547d6b086390eef15d530934115f181c56653637d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf15df6956f06137fb23eb10ec4bd0020c920c22c87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7b10083fba8c078070a0d65f619a017cbf3be87e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b2c4773b86602f6497b99f5a8f7a878111d06004;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa9af3c8a0c9cdbe89875fdac94400deb713017f97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1361132345973af65a589329927dcdeb6c82beecdd4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc19371afde6e3afe55612816cf18d49f3accc413cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1890e42bf5ce1e36e63410edc643d1bd84c18fc29fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144dd2458d7d111bfd7548fae78f38b32cfcb43aeb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78401d228c9cc4d3f880881e98acad7381904bcb02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1a441704a7627933eba235c4588a19ed363b4bf0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e3a2890cc9e77c0c876313e71a398bc4bc6adf893;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd761e7d59e4bccc51e507407a94b22a49d411e64ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb27972326568b3991b2853ab5324d1c8ace2067e2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f245a5d5ebba5cc80b3e2541183106dda0e6fabbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6000a073c64f59d72839aafda34b1f1b381297d240;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160366b5610e7a2972a90627eba26a9c8d751cfecae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1682bef6de037d0aed661a18295af5fa4ad495d15e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c81f0a711bd076e74486da558d75474480e6eecf4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9390a7104a443d78b058bd0d70ef83f6cf88da481b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c917d6792534527e0c36f0ad19eb6c338aba221d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1304fb274db2aa6f79e31f66a609213234f67383c60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f481f56c7b1ca1715dd08fe17a1cf89ef1166af403;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf1293926ea246ef94b578f67c9ba2d93c131fa336;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1935f6b0bc7bb24802846d7b649a83d5b22185d665e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h151e9981e16315b4818d4021e547d9b09fad964f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fe9697c5e58ddbb57c9bb356016747314640dbe28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h520783051cc8dfe79bdaa881f81ab272bffeab2436;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1862b7aa4c3bd867c966dfaad046881ef9f8614faf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d5f5c177188cca97cd9959d1f5e16c3ac8808f2ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e134aca79eb4813363c2eb6c0b34a5e14643e0720;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9bc41011fe2c395f085965a49d62f64dc0581617e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c205808e6e8d24a053c952a086c37034ec298aae8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f621761271f3bb26a6fb643eea4a10a9cccc9c398;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158e81c8a936d9bb85e35013965f2ab09986a911695;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bb2eb0204685604ecc4eee700dd83222c8d6fc977;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ec00f93eb521cb8897dec24e10515db7bc50d0b33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a6170de3042f11584ba4983c298d9e04d3d975e1ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca9f7e25a7fa5011ced2c7f567976e927faba3127a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e64146227768198ad84bb8e1d564c77cb757d1f3fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde518c28e04584cb204d34574bb7f9d9cbc1a0f712;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c4148a631101144a2d51f6f872933a878b9b8e095;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha238197eace20c72ddb830022157826eb2be8c9036;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4042e75a8c0b91687fd12cc389ea73225e817359d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11beea1a60a644507ae1f13c98641f41fdf6401ab95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e04bd5838d2c3b95efb34a0db4a59847985c4fa9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15120295ec7807cd8b63c55891a311d27ed31e4a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heeb5f92fbcadef67213d7d7a02bbf96f8e93e5c1f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11946856f356dc33fcf9397ea8fe8f08d6554345895;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163f0ed63b049182117a3a8deef4103e76d35188866;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132ee1c3749d8102567e3d1edfd068fafec7d88cfc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52ba2865ddaf9c0bb38bd2e61e8559cdc7a6968e5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d845601e1b0d3759d9f683433887beca871e1f95b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1083b3fd927967b60aabcc5db9cda659eb811232948;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee6c8b9d9637a690eb6c0b5b4c05f8ac7b46d41177;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150b8d1c74babdf4931f9d04bd639b8c82ac818edbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he98d398c4bb08792534990c8773795b58d1113cc5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a36a5c6603cb603b887179bb075a10289ef28825b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1efcb56d6b7ebb27eacd0f84e2ad5c755cb19ae3d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haefe1194fb6e6aa79ad0dcdb0e7a7388f18990d1a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f4d1be5c20015b5307d866fec24f2a81a6a56706e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16944254b6b30117eb38e7644303bc361d12490824a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1858374d8524e86bb897f698d1d0f79527c3ece186e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92bae93c3fd253088356e456b57def5ae07fc132b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d25f96fcd78d2506153acc1dff510df554ba8a4a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff15314857630295d964e1ead8816b5ed92d422e4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3943f68d19622a9382856dd1fc1c065868f1a51a9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e7e394107cced93f9dd1ab9d0e63adc3f1c2c11d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha02c9a2027c9e3f465b0330a685e4de32f09208f49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4bab93f3d912c7ea3f92359154fa2a5d242fa9d55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61cb217fffea840ddd7bc0080017ef541dd42194be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8bceaf75c0f66f414f632d1ee7c20b93033e4b0b13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1289a3e3da294a6d94e91cec78523a4067b05304259;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha78a3a59cf97c624bd350d884397674d99c5c963e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3ff0151f1e048b54658eeacbc48242dbbd5f2cbecc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1773aec8d8adfa48d0f379515ecb8aadfd44fc9fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde3be85b302366cc33c06234a3c1960630b33fb241;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137b8d4e611b4cca64291757bc525d856337544f269;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2955f5ee9189ce81a5765cc4a361dd97b8603520d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14351877c75ed1ecdcd4066425b2814213f81581567;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be5a5e535752c35c55d79b46c0069f77490a7a842;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89a1292c7d4931624151af486e927e7a69b74b8493;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha19d3d5d5b8240c841c8799040272b4a14023b52d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec38fca9588d219b55fa5174490b9d9335c9d8952d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he88723d94e7f7291989e94b182cec2cd21dfd14159;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95668e5d9a385e749dd3d6d346339e8b2119846ed3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf55699b785d75e5444393eedff67999c0e8599f252;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd16403582b93cb13a20fc390a874c9ee5fddf50c13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50dc2acba9550bce968805d6b680ec4159856cc10f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1c9287f0db1e0a0410bcf4a75225f1b194393672c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fba18cd06ad3788936ca660147ae6f411535019fb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10658f438ff91c43f09874e39c35464cd1d465fdbbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2128bb1fe26c570fbf6750dd997288739f2d3178c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2226ba8f1df776ac330d44f3d5683d00ac801ca8be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h773e172c0c8a77994fa55dbc548ad13e00d0c6e697;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19462fb3bc567b6489cc6e031d511be6a5506613f89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d3c1c0387d2cc72524a6afefbd9f6ee2208a9e86c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ee77c185346f4f6993808f73ca970f9a6a7e21e66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1241538efcf03f09acbaab4dab35f781f3cb683ad03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h799131c4dce72c4da25dcf759f0b00d2887749b4f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187c40e326d67c6e834f73ff263b5146f86e7023146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ea8cf785fb6423afbc8fed86d8eef225906dc8b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53e0f68dff395f61921c3871839ef4fe619b33fa54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17681b3e0da078e5c80512eb26f1c8404f3be1ae999;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82859df12c669b04bb75cdea40cb4bf3db762c9cc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32e0732ae5fe34c60485522af03bef73e0aafa12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1b94f9b96c52891262ae08c80f5e5ae78f276c976;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19aa808e4f1bef37fca79effd93b3b1d1a7cee7ab41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ddf0d53e198a68cffc571e81790e2cbeabf049946;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h112671602eb7c5be422250011f38426dc67dde9ed88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3389251a2aed12ccff3cd97d9cf210fd7193a535e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6165aadd8208ee1e88db64fd94c21612a9e93b0a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0882608800f4a891b7907831281fa13e636f1574b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e9709fd86f25aa0f89e4408eddfc3c0252f455509;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fd8aa57cccd00df891344f7f6cc3c2336173c80fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15bd213f7ea7f63a4d0393365cb28d3c1291a95fc10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a4923984ebd26783ee93e4020667c87bdd4ada450;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5307ae94d9aaff597ed0c07a3246399f785817d66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5998353465b128893d5c569a8e9f099ba9d920ca6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13140bfc3196ae62e5753051f064e65717e636f38c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had4bbb6040fff61e6b71265c5dcd1b0480dcee319f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3cdaca69aee3c97e759e21ab8800bd6c45f1c7682;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2353a5b2c182559b371e723baab340b5df0cbb3c9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33e91adf6c31c4b1f8cbf1adc6103bb2b71c847383;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d5884fcca12ce5747c309493e02a86fd53f0ddc659;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47f61d0d5d8894b6b3318006e3e6a50195e8783c76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5d8d918679f08e0eb36edd14efa9d7a16acd130f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74c77813621f17536b7e140b3463194de2fc7d8f84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ad21aac12cedcca3b9065234af3d193b10bac1bfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3324a0868d01b8c9a9cadc1bc9ec5448a58b317a49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159b9e36c0536c67c47738ac75fcb421acfc4bd5aa9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1898ab61b1cc4c666a593dfd7aa279f877763edb80f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc079e8a89cc9cca67e0d32075110a03f25d90d1519;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hedda071ae4c783265ecfc1d92dbb0e253dff63e966;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c6c909e85e50f6cd200c117b57e3d09e18798c9b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17c8ffcb7c59dace49fa27280b71009b7b66123185a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d2ab09499df9ec402fa279d27ef35e7fb1235f110;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc3bf0f804bb96bd6ee7e72d9f002de682aa8bcc2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19dd7ebc0b7888224fe44f121961ef2f663f0fedba3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he879b84a53e6941f0995e00098fa41b2d0f3f0390f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ce9c925af669d5e33d6386b2c587b0de72465f63e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14cad75f95d1a21ae57cfcef57857757e0222e43874;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b41645f7149ed7e1a7346ba4bc32f1dcf6ba573bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd869a93d938270903a27318c835b268e8a5a160dee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e988879ffb7d2bb5211481e376fa694bff35339394;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8e8b8ee8810ca1c8be84402b345db18f8e258ae46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e82b51572eca1346962d44b74da33ad190c0d9cb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118612ac60e34715cef78f99389510ad19a0a39ed49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h685e6e0900d586a11a88564e4a265f7cdcdc787696;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115ac71bf5b2483f54b246df43fab05857c1f024cb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68140c5d69eb1843b19ee3b648204ce8804e468fec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0d517f65e54fb219f1991341fffd3d374427c0d9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32ee69c9d413a04c2933c075888e490e06dc886278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha89c4ebf706c97e8f419781d9db4c1c3f4f84d4892;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc0058db252f29d08002b21c0bfa0ab35237ffb251;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118da22cf0f39457092bee20166cc6eec25b6224219;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1991d417240f646721decae552dd109cb434dd15220;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h663be5410f053f6660721c36d0a3783a9a854a80e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b23f85afb6cd061512c5a60f9e1d657571c3fe39e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h488cf5e7b3b44a2f6f58d78a03b875d7c8e6d18d3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1cc4985d9bc893690d601a2bafc1ba73365663d13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83b097f1180910c0c926a5544c0f8dd89a05d00b95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e82945a01858b2e33ca4725d8eb025268070b3318;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c854f6a2ba786ce9eade5f9ad1f31720f660b3fb01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74267bb3ec2af656bec00edb10c5ee19d60298c906;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68d90b6f84f030822195e7d75cd0815d5903dfd4e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d29d438ccdc7b352d2cdf0f20ddffd614aac89c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4091659de0a91cf6b68709ef7e45a7fe3282b21bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h267f30520eecd39cd22a453ed37cbf9224224976d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3c05ac164e32495a5ec41c1a0b05bd8593bdeeac1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2a4fce0cb0060af4c9e5e95e0152530b7bb63a10d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5f9a0be03559a16ff84681e38ce1f3e59e2308b6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116e60a4f20e021ac255027934c603d7b67aa7e6d03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0ae428fa1b8bee6e6b08ec002fbf0b5b2955b09d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee561191ce83ab2aca5fc282451bad63a4bd761f53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e2a87a62473ca4cbb4dda565892ca4ecc1ffc71d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha591fda641585088c901d4ef8fbebf4b4d20394977;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16005adebde04ee41889814bb0c14bcae854d6838db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e3e672d7a4111b1f3b21739be60c1241c4c32e998;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1246e61e91d092b31502f4f5cab3d4314847b4a65af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had29bc89a9ca3a8d407dc7b6ba5936b9afadc68cce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb302e19781e90cef956b20268fffb8c8894d7a0389;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h769cc2b28671136974c8b0c006efb44e01851065c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87b4040f64994277cf70f5e75889400acb8cd1f2da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fc628876a188f5b3a5bbcb59baa270cacacfbac3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee42f4fe0d0d70162cd78e3812eed3904c84d2b675;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165a6229c6ef01ce42fe2a04419f95bb85bda9428da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a1517e4845d4a03a92b7de56a310fefeb3f601ac9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ff97d483c89cc99ef0f3d10520968285a940bfffa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf9bb297a5c6bf4e71d15887cbe4dcce8cc769b294;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1507bc8b15b946a591ad5e9f2634519e9217626b3cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5572038f0dd869064da6c4a0974660932383d92de4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcdf03b4328779ec906e0d9cb241e685ff732b28c3a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8afb752a998eb617a250f282ca9b0fd5e511d1404a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7a212d7d3b8c0ac4ea5baff5b2a3358e05bdee71d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132b17971f28899af12499762518afed51cda2c7dfe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15121c95b507a681432847ef5c7d169cb58c670ac8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b06e1816cea191186cb49103bdf5383ed7581d31b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h532d42d0dea37dd01855aaf7ecc3eed94c815a43cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca05ef4c6ae74359754a525764054769e01cf4af09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12825d545a784e3c71310e965e38f0167cdedbf0d64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16384cf3b62c6dcfc786947e09d53c12ca436889a8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1786e307a0fd62584ebf8335a5648454aad5b4eb554;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170e147c67c3e366c4f1893d9826439420c4952d776;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b152f552c23029f1999394a159536921a2835a79f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119ea72cca220f31ddd54d8f541034b07315bcfc84f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfd55b03c42fd9fd838c3b1afd9ad80f0949db0805;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aea6a271548cbef309188ffc1207855d2230c666db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a1a43277a61564c0f16f87fde1e0a6d7801e39135;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb16175b2e742794eab479e7c9e9dd07a3027b725b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142ee38024949b3a13ca9e316927d48e7c0fba00528;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195e8bb05b07f24e5fc7ed1a8a37a9e552538133203;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7124e7bba663309ee846133289cd4e687e38f6c0c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b70a4a90b0b7e7daecb13c7f0a83649adb3402207d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e0ecd91c48cb19f0115b3a9d2797b128dbcb6e7fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ac4ce9ff1b8abe075d57bf878f43aa1e1ab0fca9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176e732ff87c257225f013669bbf3d9d1c4c46b03a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h449d6e6dbd30b1c94e8c473b8f1dc662eab85426f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10daef4c4dcae0be54d66d219170fac64e0fbafc7a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5205b4f81dbbeafbe1b5691264348370cfac9cb1aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182e34925470ac0be157c1538de85954595482b41fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9aecc96bb7dedc9b1fec470aa3651dea284a76e41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f4d2c7a5f37b49a4b82d2b08cbe082e73f89383db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h181cd9d3071c22e9ceb9a23fc87b0df7e681d4bc86e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192dab3e6000b3b5c2e7dad279c3ec127e18b9584ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1455273881277ed713343f909246dd96ce1e3340b3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf15340540579005dfdd316035768d290b9237604e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d16c4b5e86b438594525803b4f7596d6fb9d95f4e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e2f9219d7addcf113c978b503ee6a1798c0ea0b8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173ced41618dd8d0874a33735b426588af16370b571;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba0a0090f578786c82eec4257490cc3db42cfacfd3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1544843d8bd9e2d82dc786f2c7b20c9124322d15f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5c2c0b79f29f3e24271dd5ac6ec9f0497e03a53c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h572aec942f7caee537368b22b12ae8ca50b7ae4572;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9f5f6e70eb99abe5af8dc9a7e6c1009e4b2c908de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b594b83bffbe434b2ffc5df59f9fbbaf855ed5d01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h619abef19f311f45237d097bd1203b9b2a73022c64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cdb9ff14186b7fe800c7d5e75c821ae8a5a15786f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115d3f8391cc9afc0e63315219184026318e564b5a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1685cd8ba7a54c2e01c538509dc5ed22aea1bcbb6eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbbebad416d56cece77abaccbd96deeb10b272fdbba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea9c45d51f9d0a5fcfde5125f40c214ded4ba4040f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18594e1e10708a54dd68baadf575967b765bd1e54ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc12a1aac724557e66d6c63dc7a8afad4a6bd9dfce1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178b3449432368374b9451d83acfe5edc5377b20bb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197a61caae16508c758e31103d9fa04fd009742a09f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd4cef540e86ac1536f4174aa5949893457a281636;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13daffc6a371fd1d69115b74d2e79b78db6d30420e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1631aa4241de4bd42d900e7373bd858bba729789624;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11396e401530c29eb2e693048c57e0a86313fc482c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12395bb29267ee1a9e6130422158467308a79d83109;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1318137bdaec0ee53bcf59064c93387c5bbdb9e3ee6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4fb1c8b49f067035cb3ff8e7ff5677cfa29d090ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e1029c5a2b43b9f737310cc47958e6cd620334046;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fb4d50e51e466f11e72e7b74b540b5ef3b0898234;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h120a1bdb51d1095ef711b2b536e86ff030a15b77159;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he21e420fa10c2bfb09b3b41c0dcef6061cc801244;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24975f41f48a2c067bb13fa7f798890bd6d78c503e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16024c9a42d759227b73ee0f2c78e0e3b00acdb1968;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1189f10ac7e7aa07a51950c6a82169d3cae8cc63ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he284cd0b320adf486b872845e15a52510f308c6ce6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab1356f854c805e267154bafa9e03773926807ede6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f69285569baac4b7d93db4cdaff1413fd856bfbfa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8512d56325c69c836378bd24ffd2ec9104d4b5b130;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h330487e77c4993f1f1ee4778c95869c6d8c96bad52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a07449b20bce3a5f191067bf40938abe1fa02a939b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28942c4cd93a5a5d0e175adfe1bbc54498aa88ca29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea89ee2da706ab6b3e05d7c2308c39052b6906f808;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d967839eaa0a7ed57ce205e1f9db0d7c691dd1544;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157f48781239778ac224ed9e741a1be25300566bd22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10457aca292564ba6208bcd0d6dd8afe0c5a11797ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h907950a46b41cacf5146294e4b62921b434dc85bc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145fdd0adadf369bfc3634d5103639ba3ade36a6572;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a911aa4b016c184892f0fd4ff474ea9b4f02f98e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197289ba89e54f96def1c0b605a44d4b229786aff24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7aa3b051eae596a449bb4932b448641bf723480569;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2242da60a0641bc046295b7b320354820f7610c8d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167eb0e18d3ea2dcc1681ffffe1a53262bcca183cc0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34ab7f478891c16dd2603c31c7d6e8c40d68c77d62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36954538c1e796efdc0815e7060818869314ea321d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22559e1306aeda0c5d2320446b4a15f871a13aed8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b8a0074b1609a1db9ba2dfecf97772c200c27ba21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h835c72630c7eb21902247efc0e13393a5624b60307;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1e40974baf76d709de3506b418ddf3fb1c8bbcb39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14eba01930ccef1659fcdca233397901e44c1eb9aa5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ad515cd0d8ed7bdd5fa342c6631b879f2b0496523;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf39efa5f7e8c634d6c071db480dd870e88e06b195c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77705018da5cebf87c674789bec02354c78399195e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d89bc8a19a72fdc8a19520dd689b94cb57604aa3f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15bc582eacbe880e5392e4dfb1c78f8a23e60bd9e62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e6bae917c7e61d66a641d930318581d1b270810e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4fb651c95d0f7cde01a9df9b569aedf4f65f382097;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee182c8d602b46208c5ad8874b8011f0f904f79fdd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1abe712a85555b3f675c4fff00355b855a52f75e207;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15571dbf22586f2e37e0dc27ad2ee955bac9bd4800b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74da13f436b060d38224d63f2f4782c783c1ee438e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc2b6db906283289e06fd60f916806f57e635ff391d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176db35caa2994ffd114dda3bab50b84b0ae7465eb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ee61f53d128e1017d54064421ccf0db6a46c16483;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2b2ab2f5181a9dbc61221c773b38414d038501bb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc80f036cf2994313483266e37fb53184f7e579144c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b95a06169376ad1cc3cc5bc97885771b732b6bc253;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11edb65b833d7478cf776fe18e8cf8fddc8be06c7c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfa3fa14dc0a070357f7f35b3c0b45083904f7c0ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb6fe7e87283c71bc04269e88bf877459ec7e2b6b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h258035f0aa5f39e8448764eaf5dcc0214ab42546c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b29e364744a04e1d7cec768ad31fb11c5f54dd74d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10938a8fa2a327f4f215c018da5b6ecab4ff66e1007;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10fac665766e9aa010bdc088c036d76df3b2c6824ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f4f25e291e146b61aa77a60d0ce4f55228cd04852;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6d8d0f3c97049b54a877e386915def1eac3dcdd08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1c07dcb53fa07e540a4dbfa95bb5d38bbfdef1f11;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ca81382dc926db884cbc396a8336171863ffa61ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd947e5245fcf2f70e7edd1d5979145adf0d8dbf1e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183eddc0759657d121ff90e266b6bf6721d6ec3b081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18177c30ff7a15fa00293423af24e42bc0443efa93a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110a6739b2584914cdf573eed40010b06e982a6e44d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he20e1c05ff68f604463648c4842791adad5730e685;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110896d3cda42c745d1d58f9b05fec5381dbdedd61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1679d6f4e5aef6b9e19e8bc15d943b766424aa80688;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a38df5520f28c8dac85794ac906a4406464e08cbca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd0c7486e8d69aff1f82e38f03189ce49979ae47c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7a3447af9ed91405daa9c8ce9080e58133c402f61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12a0fc13aef292233651357b614b67d3c27cfc673e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15db58983e49561b64230bb8ac614c004231b0ac777;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e454972193e563f3663aa669ef639019bec71baa63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130919bd035e92a8101510da3c68c2e140898466277;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c450c54f266cf30a32921ff8015ccd2e658bb260c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha801ace6d36cba48d044536609787cba6bb0968af3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d8643dd0ed61522dd1ec14a79a5e29fb0278fd9de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf56cabf912e78e6b347abacce6713545c2abc1569c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132ae7b5e67303e46e916aa9028327311b3c4aae540;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1baebae09494a1b6d5dff98865bf6302a147427f7db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c9c964b910eda4ba9f3013b0af6ee957ba722bf98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fbebe5b6ad9615444a201fd51d45ce46caadeed2cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40fc321adcd0d6d9911079c9781538a72f59e6274;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130f6aae7b5bef51bf19408f2910e1dd92492bb0c75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4afd861ddb4910f6dab99af133317ddb2338727e3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3752b837ac84024e156bac1e95a0f8015a1d4ffe8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a0c99d3e21c8b36d86fd5481167c549a695d8edb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fe621312401465166596e29eff2b51c71adc56c9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha08db89bba6f559df5db210742c84dc84b66126fd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c16337ff81119e04888fcfb63aef9acb3a4541965;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f1094c66dc225be56c1c65783648048aa2573e506;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2aceeb52fe05141d730871b49a34227df2d9ad6a72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8fdde0b6c8cc28bf4dae9e88af2ee1404e1a7151e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e4c3a51fb9afe34155c7d49913f4065d8a4a32426;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccd23eba8f821d0495ec0969e18683596b8e606265;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146c78cd08752a16e8d4ebb7b93585092bec6e1f145;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0416f3afc5f45822fa9d5535ad4f749ef22366434;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7f09cd61263e7424ae12390b8f4d7ac9cd6d3669f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10237ede5db6f89edb63dc7a2e1658bd52391ad0da8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ca4a6cdac1efff5ac1158ec4f75cf2648ed4e29f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd2be7c102a421e1a2810ffe350cd02ff0afb62b8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h654ab7df2237af7b5217f35959ca2a9141372d9017;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h226ecba8be7d97ae5bc5ce7a1a42932dad8c99e083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd11aeaf0e7e0d5b66447c233b5f23ee785e586fbe4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7608ff1081e13d7fdfb0a3cdcfdb3fc4437754e6ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d4b0e6b1e8f843cda09fa86e918f4e8d46b7be33b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177df7771d124881935ddd29577034a36c97a640342;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h610dd82a4e4dcace8e78a021613f964a3a4a10d6f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5afb61b9dc521a94516b17f93542f43c2c09966e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7f314c7ceddfddbe0aca357719db5846b6257e1d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc715dc6f91fc8801356a62fb73d9b9aa4f08f0755;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1980775916459b1c6b29ca08198ef00bae590fcd39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf262d9201d0a3ec14eadc7f2c683e72d700daae077;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47d0649842415e0bb9f000cb6958fcbed0e98b0b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f9ed9a9df5685bb555d4738f3117f3464c364cf68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9a8ee9f6092f3e4fa800c591b49c68ee69ae8f244;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11de530a14b8d124db7a6fc4ec3e8c978d58442afc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ae590e95b2eba5d7da7849383ee9f84e7c5c4c56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef722ff4a795d3ba7444227e67621f91d5e77a009d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d0b989ed7c8a5b1df60ef8a8122310292c6d4e132;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63cd8418fbe5d90871cb2a8a51bc52ccb945afc3b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63df6e49a50a4878c88437a18e3c168a7692f7bcbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e28610ec44667cbce570725075a5efe16478403a7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19fc1061a0e259b566ae14916985b0031afb4b9ac6d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b125e4fd00ff48a330fe8d0147c7b70f0d0418819f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176f83a33123beb62d3950ed9c6affe92d18f44ee82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f28cdcaa0917023c61dbfa6a4ebfd0b6a12b6f5f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108b64fed52e55a36c84df4ede80183c35a33ccfaa7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb214ae4c5fe178f5cc515981e56529d5585bf4be2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130f4fcf3d786d56b04486aae39f57230cd97b5c852;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cec029395da116c7e75d076c7ad046acd2fa49f450;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192a4a26c4fb5aec20ca88574559a516a66654af8dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53585ad0f2bc7ea241ee6923f2ab643b6d4ee0e9e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fd379cee46b1714270ac160c5fc1f4c0788829a24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e7e8aa2ba1e42b51d694ae2462f6c251c0d189a97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h486fdabde5a305d09fe53b5fc7f818ef6438e05ac0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73e6fb65d7133a52cff1c41e613c60a665859fe4c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170af0b2e6d033366bdfd881e03596a1006a50a0700;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ddb9ad72aa25b64d478331ae1147693993d5d5a96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87c2f1c1fab254546757b2086be694a80213156579;
        #1
        $finish();
    end
endmodule
