module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [18:0] src20;
    reg [17:0] src21;
    reg [16:0] src22;
    reg [15:0] src23;
    reg [14:0] src24;
    reg [13:0] src25;
    reg [12:0] src26;
    reg [11:0] src27;
    reg [10:0] src28;
    reg [9:0] src29;
    reg [8:0] src30;
    reg [7:0] src31;
    reg [6:0] src32;
    reg [5:0] src33;
    reg [4:0] src34;
    reg [3:0] src35;
    reg [2:0] src36;
    reg [1:0] src37;
    reg [0:0] src38;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3])<<35) + ((src36[0] + src36[1] + src36[2])<<36) + ((src37[0] + src37[1])<<37) + ((src38[0])<<38);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9980408e5713b8b2a1332616c249111aa2338d2b1ac5b5a6db35cfd578f4fd1b0d92d593bc87a11b6559d6725b656be99457;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf037d99f3c5c0ad135e75b9c44f84748ac7545a2fbad87e07cc2071697696246ac52931c2e336bea26b263c0f4e0b44df05f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2750b44fc973586c251b64de7bac97c7c06bb51e7a94c3ef689840cadb768e5c33771d195ab2b6d09a8b6a182755e6e7c57d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha052eb63ae4895ad3a0b6fd801ca70829048c21df5693465bce7b362425b49e1701750c26d8fdfa16ef727477d3fc3a6513;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5367537100d75e0b10a53ad28d72b74d7f09eab3f9a0aa229db16d2d8b996c35d7cdb23fb27830314f721b95ff9d0b72e062;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf25fa3a99315d42994659aded461082c8c2c7f589f7ba4d41ddeb6ba6e08eb62958dc83e044bb72b559c357cad82a33f0625;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h106bb507230cb42b491ec83a39d91b63bc1413ef9c2033e9a7c94194e18685df9c56df9f38a5a1229f6c051f9e26c6664004;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52c4f38bc1935309b9a6b81b0865942da2b0de12976fe9c2caba0d20e5769e1ec70773d14b3fa91362c1f2b6db94e1898247;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34e8ddb22e23bd13c6977a8afc21b23b948b4640c39125df8552a995a3764964f07a69ae59089457176dea537b9c0f5aff86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6740e76174c0e618d0aeb3dc114389dac62bd25bc11f9e03e585f872a62b2fc464e38097ecc25821be7f5f83151623752ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60aacfd619d674f425adbe5744e9e87a2af5c8387475bb113638bd8c779f6754fca3be2908d98aed2264236eb619665e7865;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc222a6eabd32a024b345797cfd80b22ff4cb786bd27a55aa1e76d1b42fe66a675796cfe1e16a84bcb54820b951bec54f7e28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa6f07650b28b1437d665fb1a7eb20f91248c21f398f63e028ba2f9e721de153ba6f2db2c0e68f9c311168a3fe5dd251b561;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heea929d9b0b0df532fae8507c2cb472fcfc2920bfdb06ca75ee06203a62215616952f356c0a246b725bcf67dc375a181b7f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d9a19439ea05fafc010d140b2b7d16c0a5627a421f622674d51e863a2454a5d6894fdf2de60c5cb1c20716ca2f80135b29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6dc0c1d6a21943ee777b2cab3ba32272699671d91fbc0935c4d71b9dc18eb585bd78b5163ccca4b0a6fd6450b8d46bcd223;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h792efbee2e77373d6e918b9689e65a4f9b3c5a017dcdcd4d2165618b4d9b20eb3229631ec2b6cc3f1573724a745e49c77bb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd514acfe259d2c1ae3d6ca9fdc1b3e11d560e19a3608bfdcaa55df212f65f6c91344d564b1aaa908d35d229ab8f1929941ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h127e363a7efecdb773f79f3a4f4e84a8b71769aae472f34c1cf481d7edc0f33ee3031525d5ed04f16ca698859c8ddc9e12c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc1334f6c0823e0f1512709dcd73adc0f6e6dcd4eca2dac6d2f87276558826656e8b9318554047b2badb7a40b6b74cfe52ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95d32d568050910eb5ff994277b449ac85f155d10bef627828ca09051cc43616090af0a204197c69bdbd6248ef7173eae235;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f8c6da8a4a2496ccc89c559beeb70faed98a3a29a42be8a9a84fb5ac040bea072a18c1564e232f0a19fa185c50480438864;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c54e729f7fdcffaa03052222190092bfdb0fea54076941afdaef990c4148f6f48118e09f02a5421b599c033b540575354c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f153a13bd7af575ec295190d2e8e0d716600bfd93f74ecf8a9b512205da37a05ea90b7d21dce4a053c03c988b89419f598f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8c5d0a2b652be75a9eac692536e9e23fb979a125e7a0f23b5b2730ff8f6d4e06419e34b601e1c35797a933266903b180781;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd289d2130dfb3b61a7f41cc403a8fb686ae581842bc473d2c11a1c99f2edc603fca452fbf1e03f5391195ba0b667472f36b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f4fe9b9959cc7cf417b448f126165cfc0a4cbad0b1a000861ef679a534878242dec3fc1da4f51a2c00f175cfa02d91582d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47c96b0bfc2348c9916006d23f1daa9d6288857961ee129c8f0ee74236dfd6dbe889baf341f7cf672ac4926cb9204fde9539;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0b0adc7f5ce66d557dffa85a4609a49af0d416882c3d3733ec1a6e7b463420646fa619599a5a596d1b4be9b76e6cddf8460;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e0be52bc90ce69f00392a67eb6b17c57162fd963f8b3610da50ee1c82583b5aeb99b29cd0f588d62f4a5d28ef238dde1f5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8575f19fad335c0704e9ea1d760eea708b52195a5c28ca4b984eebd48a696ae302089f7b42e9a4902b589a9e07968629f0ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h537f949a0b6442bfdb8ec4f2731a52b7e8aef518fa01a5d32a2049caa4f8f96808f2e3653c1b436c3d93f1b9795c6fc00f88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h843a02d9dce19f28fa84a71c4697d0d85cb3b9981523fc92f61eaa2d50a5df7b843ad6135d31ff80bbf14a005821cd051edb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8b95675398305228d49d9a0874ec1f425234df63b14e339f8cb50bda13add5e9081d048954dbc09b8d59b70c363ae68f4c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f8e702135d4b506bee924283c4c43c0643aec5316e4ddb608f858139caa0c6fa2db6be59f1cad8993778a22359393f16c49;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7c9ceaab413d604afedb1a5ac9b858fb607a78d13462cbbc289f11c1f9a3fefd559b66821f6d6d2b9296c76c89fa8f67806;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h457462bb73ea9e166d60e60add138191c88eece3477806b09682ce26f2d6fb524ae9b39ad2a61206c8cc28e893f1a455c9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7cb9e7e04bf9c18e5b04c03d2fe1e0e38b1f752d278bd18a1fd49e6508eb579f1d4039183f72d0b19d8d4a1200e9e6b961e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc767be0e6b187f327ec748d7c9bdf8bc35ae2c5db35dc8c63db4c28c7da3c94a5bfd379b0ee2c51e3819897a4a53c392fe0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h839be23ef722aaa1a51558f45e5ec076cd212d0ebd321930403c567da1bd713a95d321c9acb712859c889bc69fd65a2e5543;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h121c3e5b550b9ebca54bd7e65052c967df75735d437238c97e64a625cbd813e7ab228982c41f71fdead77bf5fb448679c742;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6064f5c66e281a60a2d785b11619a2c1dc5d6de3461b936227d98ce028367cbcdb46f427d2012c8a018f8361b8be8fa3d4eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfca2ea4ba377ca78510adc17feb357af62e18864f6fdd60964e59421d65f7f4e1e52d16a6d8d52c28d425e594500b10e3c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3ed1b15ef4eea37abc97220889fd3770ae96a4e4f02072f670209bb96c444a4b4e4381af18aa33e885396597ab5c2e0a527;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b2dc9d7a8ebcd8972c871eed82be79ac667989a297128a1a69e593e3bc9679389ca2d059fe10b2fd11976bd1e1adf2ada7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12e201d5566017ee93da25f7ccbede630b9dc01f30f19bdd799e2f8a6d317bda899bc6a3f50c87c825e3f349750b7e85d5cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25fe3b2e24b84e0f4722e061a60468d4cf16eb4ea4b9c55b468068574cdcba9edc7aa2f236245d1d80cb78e5e92403b67f4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98057274a10cbac246aa5d24bacf6b5cada70d05a9371d92c5fdbfd5790536635816d30aafcef24ec839bdb8d7efdd58ec9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9059ef36f201f68df06f6d43f7117bb4bbab8be455be70e5e01215d940d205ba87193afcf824bd654baa2cf36749072efee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b1ecc11110206dca73c292c65766851add662bf97f864dd48f831d66740c62bfc02b51dc20fabb5a83ecd48a06aa126877b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeba1192d53430a663316a19b87a3108f1250e63627f37e6b0cb6c83d6752b58374bf5e518f611e539fa1d26f297b3b45e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26ec6c181df9705298b012e1c4e4ac6c299a50ec0ddf785a891b5d7312eb9629e92fa8dfaa4c28b4ab8e6f69635cba19e33;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h884cabb938882fb36a31e7ab1095ae87652128b1f588ec24eedcd75c2c5ff0f538c0a777ae05c5a9727e7906d3a05742a28c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89ffcc3eb9ec890c039157e28a5163f1e8dde002052f006e69cdce3f167da50e462c73d51680b1a12414adb30cdf20d7687a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha07f142330cc1b3eafc0a26fd6ce34366b0041066d595b08405b058998660dcea1d8e86902f155b22e0aac0a216755b036d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a2d2ea0967048653b53825044e8176454a54fff40f542c3327ac8c582347ae25f787debdedb4af3fefa2ea5bac632fd539b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b62fd020552ea747b1487233e3c398b030ed04720337d72eb1f682bbb0c2dfdb8716a0bace385be0d4c6f4615ec2e8af701;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5fa5b0638527c6aa5119e47178e1713859886dd7d7b27f2ab631e59387af165009a6a8cae27635eb10883a5d03cd794d7c66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40a15031d37c4534f7d64d11a69202283074faaad01c066d0d0277ea6f2df5227a75e4422d9bc506011f79db57ac75e30263;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h282c139c7f2749054daa9b34e6d9d463c54a3d3b6cfd96f152bc804dd49aa02d77741136d1acc2f7ea7b933dd503c2910654;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7abc1fe8e20304525fd2e9ec83f29dbb930c9ed71227c26ff038c13138f5630196268c0b15afaaa0187c850f795f01543d0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89a68779d08c1063743b5b2630763467731970f8230dcc06c5582eba5db91d2e73d4de1e76d4f05043e048764a0e2dbd6a57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1e09dcf71f591ace8e40cd147bb3ef0f1359e346786a8d363bd959fa448b52b07b3140ababc6512814c7ad7c5ec05fdc4d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h262a4cb9d3a9718d0413c8cc96f364605cba5630f49feeb459341f483ede8378acce4ad894d698f920aeaed3d69a230bc87c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heac5c916b60d5bb3f68477de3a483e70614ba3f3abf830374cf27ee3928820493f2a3f5a981cfe4f4d4dd320757384952c57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17aa29c13cca3f047e96ffb7d1ca45b24e9c66d2788e369a7afea723b766774c7c09f2b73b25f44654d18c64efda06b0260d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e24647e04ef3192b83f806ada42a247fdbf25100ba18a057a0c10be89d217ba1b33669ac8ef3ff8ec6927a61827fdf4bf81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3331adce39ae86f185aced30cc960d2a7ced94594bf1cbe75dd5155278d2708b1f6ae81cc1a35d2e55414e8fedbb0c3bd2c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf19fd9d18386e12d30ae056fdb9b99d0a09437c74c91e9059c268c10bf43d845d4224607918d5d72d09eda1781af4384706a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34d98378c76aba6a10a98b846ea2810d4007a0014bd6be9da296a57725f2bdabdf86176fe0e6fd9f947731b59c946c5be7b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c8283f709bdd65888b829832856d67e6b12526d690ee014621a3059c5598d84b1dbf27aa3cfd4e9bbaa4977ee1f92acdda3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0e34850a80618c9fce70259229561e400e5c24b028aacd022be4b3f220ab066e50ee9dbee19deff7719fbd90b07001e8b9f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h630702a85b159832bbb1b958b928a7593153af6712911020abc9df2e1569f6e474ec60bf2ae10f8e8c75d858495b4cf80499;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40a99bcaafda979296e03c136c9e7d5368c8485025c4feec5023a9be3e4a19dd62f03f9c8eecb471cf79dcdad62700755adb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17abbf736748aee6bfb24a56b46cf893a090b18537d1ca106ccfe12a77155d12fd618069ac5c1c8ede99da7027c4b7ac3021;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd371246be3ef34f347e6c9b66f034da3c09d8f73557129a3376791fb393ad845ce0c77b5c69dd7e9d19c02d1299cced9bcd9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36d0f67a5565f0b0bc4a28084a5baca5fddebffd3e3c0d76bb934c9211ed48de5ef9a8f395792bc13069aa9781791e43970f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2da890de65992b51c46a53bd58cc1821af0ba6ac6606945f5b2fd0aa9d14a76bee5eb4283762b1dfca4aa02c126a3d156627;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c77f10247b8cb6f6345f2bd7bbca2ea11492df1a8122ce0c4154e0a1f5a53d3745aa9bb44e05401cbf97395c835d64aeb54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d2fa105d6685cf585926876451ef6b03140c9c24188bddedf9330c830eae3c243521682e5179d7147ee09ebc5727a78a1ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h736fc9c6c84ee19d22e3ab0ce3898fd2fa957d2fec85e65ed869f4f36a1dc056bc21daaa34f86f13b6ff5a58a42142d6e0af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda2a252c1d0a1364a45c1b1493e82401ddf1cb82f226d0edb9750043fa5d096ec51572aacc68ce28a1b9ec6ee81d128134f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h188738fd732e867f097f158c92e01efb685a209588897f5e85001eaf91f37a5558710931d7873d3b3bf2177a3797761b829e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80a6b08c5f2ccba408934e9877ff6a0b4aa0b794525bd2d1b3bd1099a22024356b111e10b958aaaeed95710b78f39f10d44d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fbedc5ce5ab0b38c7efcfd417623306f900d360f0fa068a3c5982fc43dcdb42b524d403e8c83d880502f14c3698286d7c1d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha950a3c6355adb09c3961e5395171a65b53d4af11f0b79634852a6af64f91a0a2329dc979a05c422ef2b47208a9797a08b90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35ff15f1d466ac9bd5371114d8d554fd7dc049584b311bfac8599d6c224f196f807a9331623d19defd6285666175d37d8bb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h579b1cadafb49e5880f1c76ea1619e4d714f932a5cd219f85866d0734ceb12834d6747f6f3709ccf3c67ec4148a9b0105bd5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacc3dff57e0c147854a5ac68738c50e30a813b6ad067750a91685ca578fbf22acb03d1c81e47e3f1941af739dec5ac71c7ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1f5c7ea1ba75794a300c0c05c126d782e9d140a5b47bd1ce3b4313fdf916161c742c77c4a40301c941aae359ef05bc3ef04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc86d7b24f1306c5c111a1757f7c151068336a2118012dc8f3d4cab0b726c135404c3f279681928a207025594f0a95806199c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d619abf390b73edf123484a9219742f659a2e725b2a6360d3560ef3c49d90c21b60af0c6ab14f477d52e25db146ea06db13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33826e8241c8aa0f3d2c49fc7de7285f64599907f68bc3afa3fea6480d872f68876d4d357c54367a785e558ab9489ae24384;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73af7e07e09e06118c7c4eee3f80aec84a2c4cd5d9f1deda2911b162485fbb42fcb4f6827f5193526fce87d2aff60fb8968f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h745d9713e949c0b0977157aa56726e3f67fcb4f819773e93300830fa34f8229afb740598efdfaee8361e733df3d80886bb40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe69b2f22c1486d312c3d330a4eac68009c3d7e9f8d4f34c4f1c172dbc086f3eeafc34eb7ccd8062cf35697d8bb0bc49b90a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f293064c998e209cf775ce2686de7a85abf1b1f13bc3343449be23009ab3c202809459b89bd56353c1188ec82b68b916f4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h274d5844cedd1d77d9383c0cc95dac7ad47a579c60cee78145967ce6dfc4d5b06376d47bebb80fbc05a9989036a38bc8a1d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbee2e8aa679e064b81644490e1853be4aae792272c221f858d9a13539862b5f09dd343ab475d5651dd411a11c5566a476e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae7694b3e839f8616bda5a41a729d9753dd7bf712a0604b6b5e2de3432bdca5a02cd37c60bfb28249cec0414a888597b625c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72e4cbbf82aff54ff018da6794cf84ff46ff6111f45785e4193bcc7c35732104258985ed5574967c33536eae454fa02b739d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h516f3611396136d9922385818ee4e5d6846fc41433414e766ff76d3345292b0edf61d46975299ca0e91833c8c0115da9de69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6047f23068f506996992387392c3a2c875f060bbb59c7b27ab20d1aaaa510debe30c6175ce10c2b6398d0bb9db27304555b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94ba93884de39a959c1ac72a7457f67b25b841511c76b1d8504cdbd27c44ff8168518f5dbca543d58efeb61a213ddc5493e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a612d9afef57ad365474d219a6cde9c4e1553461312891a126fe11d6dc4ca15d71bc9561a025cb9e1c7f934d172b82395a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d7033d83e780796c3caeb5c5c51f70ecb9b980d2fe291bd55443e0c57870b2824e6efb6b2634ed4e7a4c24e3e3f7ef3f144;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c7519d6a2a8191956c717114ed5abe7231d37b164cc6ff490bbe8dd460842f8f475385028e5733a7e8431cc275cb8aadfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1655a34b052aaba569b8446cc2cb01f65a963ca8921953fafe1f5d7bf948f38de1c178bc84a31d1ba440fd6da058e2ae3ebd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14b44822a5fec95d9bedabcb27e2d92da7dee07d862f81f7943bba35bbec3d8eb82677dea15557db447d5fee700ee9bb898a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0d570f729e0d501e43a978f8c7213e674dc5a84b30cc189e440a65d9a140ddf96292cf4b4c2847c2bd4d13651fd77973f74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c1dca352901cee3c59cc3f046c2001fbd50a79af0565451351e41459e14b3ee7c9a84a708a77f4e5611e115d8df0db3cb00;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6de5ebdf9c9f3ed1971439c6f72a67a4222d80f5ed88850ce1c4da66aa3176e42701d3cfa01009f381d17b35f81e206fa802;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2a1ef5c898cc41b2e1d52f0d541964ad71eeb3fed7448f81cf13e0c2625337ac1c46fc0b751917db1c3e112119465f329da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he508cb89e8796c27d47dea13e88400754c4d79a6a22fc1772b232c41120e4be8c917a5b2df5cdb1d88208231d1648b196723;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6d3578ca710b5f12e303b31713eef64adf5f70abfbc7df7a10b50d850ee071ea1ae5943e6b5ee35292db4e7e22019005a9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha309d9484875918c4c65c8ba32b84348befae6f3cdd046275685b6a658b376b8fad1d6d0f87405052c4e591af5f3415aadb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7233aaa2a99634e2adaada702dd385ecd06ce3e5f8ecad5795f5296da9b685ed4cf5ae163bf6428c252a71c119e30578644d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40db4c249cfe3343939d0540ad4d802e3441beb32a973b9cba1428c3e44dd8c4b97c0c2d7f1ee2dd90c89abf0097e1910f93;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d366b9ebd7fef4599594612cc13b9aa2600208c847ea616bb140a0037cee5aabaa7cfbeafafad5a256b73d282e6982e153f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82925bbf4210d39b12a2472e437a67775b6e10e5d77ceee0fda46262b908e88ea7892e8df554d4e68f329b71445ac4ad9d05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7420a22c79c09f21c0d28072f17d950d270af0592c0228dea07401ac66e138526cc0cb7831379e9713371206a3a1bb790541;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b70ccbcf58b621091fc0db139783df503ac28e741e4702ea7fc7494615d1695e742ceb485074829fcc160d6e9d895e236a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5c8dea9c87b04859314d44559402dc1b4d17bdc464829274ee5b01970874b3dec41ec4eb412622e9620f90190eecfd6d20e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe609bfd9778c2d43a4c45f26238d4f47e3700d6f087241057d207d997a9d3244945104161b83586e9542c6ba7508efeb7b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha73a39a22cfcfbdaf5728116e74fd769fbca8ba53a885196cf2294c0ba93fe386a7b73532770a6028bab90db54860583eef5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha29db9e9f7caafd68064b5a0824e1be3e3f2e639aad7e31b7fecd5fb06829d67afb78a6fe34778eedfb3ef7043e363991477;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc66bf07161b826f49e937b68cd41940064f73d8120eea185ae8e438fece741610c17e2b672e82f641a9cbce3f24abd243fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80af2b2a25bfa7a709f02052541a8e8544e6d63e3398868810730f92c5f133d2b7beaaf98fa2489137e77c49fe6fb5a42722;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5fc689dd107c5f463944756cf21da45a6bebf362bff43e5183d456ed944c6ef0d7f461145426b9049638788abe3884ec0d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7254bb92281376f06d5403a6156c1fb0015f662c75a3aa9f7e9541148d054d40a7528d0214b89fd763ea60e7b8e698d3f219;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdcf2fb4bd045921affabab688c391c82951584b7c2b7db9c815478644d57d053249830be437db3a189e98fce93d339dd9dac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17db4573d5bc5961e673786b62408f7af74a6590f7da023a981590b75095dc9f1bdac2a09ec93e95452c255a2985b719a14a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8405f21ec9ba576250484fc9e809af341cf5660d425f99e419f3a5d08d454a5ea88d9128a401d423a29d09728bda3d3340e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b5c64ff138cd35c4ad05327d7520c94788ebf8a1198b9d5d58f08622a23d9d0c7f5da016c1fb5f474de02e8ffd10e522e9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22c378f69d49eacd91993d301514e895cedb7515928785ee758760d8984a5a3315561c6944eab85caec0d0925b5bc1db2793;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h518d7048d351ccf4aae729a17309ef95b28847a53e8b1e2146ef6ac06bd73c3438040eca4818dad8a5545f8dca94d3c87cc5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9fa90f7540cdf0b79ae27409c2b4cbd02b686b4cda6aa9bceab2f72e4217312bf785d4756fe85c6e5d0a8cafea34264436c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h154d42d9892d3cbdea2c8ebc093e961c0cf839d42e0cb6da863aafc09431c636921cf0ed26f4fa5b63b2e53f3d23d11ba459;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74c516c09df24f6d0f987ff0667e7c34439af8a4b6547c8de447dc8f5dd462d10c53d79ecf5963b4b394a4dd940f02ab41c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h982794e6c69ac950cca7f7979d16366feb2165456f7341c446851acf2f94c6f0ab78bf3f29badcbe2c5b7ae7ed3ebb35c724;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80de4eeda03dd4304294a108ff7051e0a0e55d69e8911084e673297ccda3cb1287e9f35ab509ebab27b7b5944a0df92e06e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70669dbf95c640df0000e729350f9a9f29dbc3da7d26119af2ea95908f432f7ea0db81f8bfd15ce06429e78f169dc68330bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h812e77ce87b0466aa07b95e6208985b28ca836d7ae28b323080f05e81421e5dc1fbab58d942bcafd5d71065ab49493e29a73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha94040d7f44d256911c985b56bc3f13760f36f76e48d0e0015d958a27f24590f8ed7520fb5c2f486f7442bc52c63c7193430;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58efdb361303ae1c388325bba2b50db5a48c2c683d8d57234baf16af282db9689e2eec2227f795161193a45eb173fa67b4ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57e58917a527d198b51b57aa88e7182fa67b5561467b4fae6bc5545c886d14982d944b44f63054e1f04e999a48c77fd7e1c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdba196e51db1519eb4c754c15ff8b97f602757897c1df44de2b3d6756972f93ad1598527f80cb8e340e0d5b8716b112297b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8929f04169e9b5454c11726c9c00eb9e27fe4ddae0111559bb2577c886308771f510be9a3cf409f6a004b9e7e4e6592a9e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68b9f9a49e242e6264b8fde556ac985d03ee9ffc60ecc5f56583f69440d1f1b28dac4a25c373694a459b835cf0ead10e5e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b2dcf3de6790949b859850b822fd595e2552854b52acbfff9e752470a89e1cf8ce4031100e6cb8dc44af38e24e2c9a859f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6f5978190f8cfc00da488adf0d6a4f31e5c36193628802ef0dfecd70c6262b50ff97d155b8968aff70f30370ad3469bceb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadbab3d6a13287d55cd581ef8d0f822552c026c7f854e68bf065b9dddf27d4381f773c07dace65675afc9134429a5cf93921;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9af94a92ce938022bec6809ac4e0038b7ddfe86d8308f1a83ac3900db3762a59a3396353f60cea62ed3bb3d986873525f140;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h475cb9cddb5c3757b9c242e0a9c062d399d5a5d54eacf4bd4d16fda3109f44675c6bd3bfaa66706c04916ac4de86aa1f36e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1dfe90934ae0571d36186ee151c4b91eb49ee4667dca37671088a420b571db08e3f69295cb69ed27c88264a765bdc736b7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fa7f22fc1a3eedcf6428a506f1951939a5066f4af5b69a3da2ec7496a42b9fcd7ad5a89d49be64603e88f53a3c7a1bef52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a42fb57a282fa76c727e02daddbafd2d64d549f1f00a9eb0e3c5f1546fd13f31f56d1e5bb3d213dde0a5df57882b02b6cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9e2e7cddbdf1e2e49af2b1dfbefe438e56000c6fc4c84bf040115466f217481305a4bd831437b6daabef977282dcfc20eb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5084c4bd1a8d570eb745c07aae84c3d92d1340868956b4d117553b6b294a8c5527e4815fd71c8777510a591c26a3d863429;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcad0edf623a49ed5b3026b97ae04c89371339e4a7378e12935d6f157f6ea96fb6965fb94fda572607155fe78a44ffde79088;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f2be826367f672aeca6a57a9494487f114ee9059408d397a09bc905e68a236c7a919c230b6b314caf2a2e569a09880b64d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca0938cb77e7fb2eba4a1fbb0472dc6de3f4a654ff146ccfb0319726da845b4c42932c50b5fef08a051c6877e7c274ebee56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfddd0f1670e306147639c9a8cfeff08a00e3abbcc9163745ec7302b345653773e1fdafcd38b74dd4114353c8193b82dceb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27f7c737ccc002541ec159995fedbdee3932eb567f8461177984d09cef79ca2f16d97ff22456642311f1a47d6feb1620e284;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1503a585f6fa413d4954a8650145e8165a69612d9876de6ff2e977971843ed05a561797b987b8aad7eac01fd3560e92fe3b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e6a6325119b7fbddecdfc267f0551626c847c8cd68e8eaf78317e95378c609e41f8fd53f1e4d09f9a4946b29784a97c83b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1954ac70c31a87f9f3d33d750296d0f46bfe8a67674ccd3b4b2d3f42e75c7a907a6f63f300f2b503ad01ea61db082e85d979;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habbeaec02cd15cb46224e0155b3f69ace614dac59716633fba35365a80daa9d94a5c995ee4e46017d9328eca40d703cfd159;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa725be0774a6573ee2c344ed37222d998bcbfb85740335b3b26191d9c5c45feaa6e4a93419753d8f78b57e630869213555b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf942fcaf7e1863b753fbb14743f75467fa1f98988c70b74f0c9df10332cd78977bb33343d7971c564045921eaecc9a4bed8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d8580e2218216d0485085d8ec6633cb03afb31c7c88bcd3f42cae15d66d6b6b52e944c461b8a72a772c9a229b888c9bbe69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadcded0d5e5f483e351fbd3949a7cd1825ad972b1784da52894c75a6525276482dbac78976177eb1f013697d3186ad51a11b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b82076d3abd2402d22e35013fb3a94004db35a8d6c7730a4c4fab51d64a2de3047e81cc063c04c505d687f560a89234a82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h973c31b3bf74f92042a3fd5dc86a6bdd283198f3edfbb63a1b3db8db494e4a0a50c07d125a2465333141c052acf53d52c157;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c889e641762279194ff7b33a18c2731e294de1e070cf9828a4769b4d934a3b492238dad38d404cfd34fad11f444c2b57c10;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ec1b03c6dbcf1d239f30e70026fee7be9fb20299c43747486efa6f521c280d45b1b142154f657e8b74a8f90ddfd534f1574;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9eede0f8c17e5a75c1143117995ba18b0682e4a5ebda198c8be5872eb946e51307c9ce8addd2027cdb95b961dfb3997ec3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h568483721207c9769a1699c19a23b9483afff6cad7dfac3a97186b55669cd6f714a182a0bb0788c943f5b77f1f57d1d87fd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83a4439157f0b53df478144ff0c434dcc4c98da2653162e424cde172dc2ce4d98615ea1cab90d543631f400e0734626d0b49;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf6eb40b82103547c841c26e41a867edca28a4f7ceddf877f1318e4e3400f89adf16e0fdb7070f77a05d7de3d0e36fb6c692;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35a613ca86f8d282a27011093983cb869749d7e493fc374aa83cba7b0c780e11feb5129f096bbc302c35e2aea5e1c93745d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h728e3487802576186f93a49c996fce1319de8de1da256e843bb9c23c51d9eb2e53b5d66d85684185e0312c884c3171b21429;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf21315444b0ad4956f344e3f9ca8c2ed192d2b156482b56e5e0b422e94a96dba477657508990af81b6c4c5972fa84b42ddb3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfe90ce9173253360b70a84b78d953f89241d25c7ea3471f8f8a3765141fb2b3cff46d08b949a0260ebfd1954d234bbe92a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h803675d70f9efeb94dbcb3fb65aadfe83e1b47c5b3f6097dd5ca8dadc5e48073a7cd4596787fdb8cf71f3c275279f4dbefe2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55647785848a8a900c9c379fd0ffcf3e23db5d90fa417b561132daade4921c1d59795dfbed3c14c152117bfd614cd5e860c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd5647b390b163524d78cf307166831225da39042c6971a3c6242d3ccb9f02917f0db9ed39a5a67cc23e7b6e437d5e827ca6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebbd61f10a24c3d235d725882c60076af4a4a8a71b1d071423f7444e842d2a570d554480d83e96a952eaad23ae588ab33c97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde34368cc7daa3407d88b7c6d686ad5f1cb53ebc24ee72346125c54694788c2588fdbf60cd4477317da9d6a93f5322caab41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c214a0f0dc28551e3d94056b7e2048e7fceb90fb689f645366d7a14d450702468107531ca2546c53c79033626cad7e36e8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a7c8e8668d5549bd08fcda86d6fd36c43790f36647ea556eea95efc8387cfb8f4280bec623e422257d757f75fc4c61fad40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0e21c1a3ed400e258288e25dd0b8a0476e8b3f037cad08818e6264de4ae0ccb2baff7d0830f199a1eeb18867e6da136f4bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha52751973d54b4046874e9b5b71945fa8a0af6aadb29c1d0015ec49a6fba9db760371bc4ff422a480661bfed279b7e62b380;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f135cb218dac25e2219f8a0015609db0f3b493916a2c906765e06d8b6b81a96a78b3df7e5962870cc56d7f919e2483891e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5062c337fcdb6c759450061863511ee783c413bf2fddcc5b66a6f687c91f27fe306c97af30b8777a0c71d83b58ec4799dce1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e8cc52030dbef1f0a8608dc6f14e5306bf8e14f85919ea2b9479e648a79e2ae0bc4bc6f13b5e8b01d2d4360d36a5b7bae3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e7854aec6502f153dc64b46cd29a7f3cd81b2b7ec6eb753c46ebda6e3bc54223d3083def54159d4d046c373a7591bee7e99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bb99c09191b4ca0e356b5b065976d3e04693b53bc4376cf18218d95e38cfe3e5f4c7d9c283ead359b6eae9ee213c36def40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b36e91edf7c1d7d572179b971592c34c46f28e5d1250f51ae19a755850be9e2d22ce50668a0d3eae492b2aeddd26e0f338f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45526bc031355afd5b81f2b83bebd1c527b991798e35a3c412ef2aca71dfb4753244715f629f13b18facc8c1996c4c20a0b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c6db67ec472c95a025bfbcb5cca5afa6efc659ff24f55ae9147f5bacef1b98a26c370e8ecec0b6e81505b8b9f334bc9a468;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59a5d8eebbd082fd5483493e4db49d1c4813958136083e49b027d7e235b5506cac45c5d4200c25af0eb2e597c095370acfdc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51b1c59a8b9c83e124ade36b60c8eab51a402ab054b6f516ca0e669ee655335e00642afce9150f36744caea28ea24c9a42dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f4f7b84958485b2b19ec5910a6ecf5a350d4424f07b2b0a31f78c1985bb290cc05d849228d88fe312686e3012a991d40cf1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cb1047867c3a3f00514ff7c34794878f2bed180609c9c5d858487389239233b1728d742d7b6fa1dc202ab991df6d9149d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddc51f09604c7d014659f2d731bc5b42c9c9fafcfd836ddb233cae138a58b74252abdb845a07bae9ca1142176e2720ca7023;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c8d034551dcc255c06387387a2690327669031403b189725ea05cd5402ff204bfb762dbc750844cd1b0145eae4af75b5cd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e733ca088dce7bc4e537dd581da6a2b87254cded0e8881acc3f4adca8f1e90d624606c3e9f005845951da891d328fccdec8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49c9c962ea9a2785af4dccfbedb3c2c2a8f63696bff3bd51b8c3bcfb95150f9d415d871dfbe672f69416b8d957056afdf93e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f958854bda861f1bcb4d4f33c5c63a0c5759bfcf6df26fba872f62095ed1034dca3a6e6fdfbe59b154cc1ee4cdb23ff6c57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb552944d18117d87f872257f8ff152e57f8cf5b95f485833fc08c7e7d482182c0d358e2563df2da7a56f62ddde586dfe2578;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h298ad9723ecf36001194303c0457114b5f7cb164d4de3b6dc619684db74ca5f1387c13d7f8de3553729339d77ccf585b3a0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5b62a2bfc4f397017675104772ab9d6a1292e2974b995cd7f092adea2baec6a20ed5e7564bf0f65c39176fba190b951d635;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf331a9500ead7700dd1c2a994181c7ece957c67d73987f60c58680f0b2f7d57fb1ec0d6a091130f87cc5bf3767b664ae1c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7da14a2c5748237f95d8ac94cf160cfa0af2a5eb18c704501343a85cfdd1f771ed6362f348084c43facb6bc28136a0846b55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3594ce8dd801e4f83bf965eca97e2fbba5dd35a5b755cec1ea36a5ffcec511fe8b4b194cd6c414882d8c27379aa06a9a0158;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3106455ceb9a319bfadb5053b0a80ba6e6572bedbc3efe3a28996c3578c58df034f084279eb241d2234ca51517ef816d0103;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a495ef1c524809d1b42be5724e13c077ea62e6a7d6ae17177edf3a4dcc847fad745149e570a0a24e6b93032c1b0604d776c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40845852d6f006f23a48209957861288e5e9e7eca90c8dcd7db325b27a6813c758ad9dc647acf42ebb45bfdca6a17dc32e53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd724aaadd4cc21eba236a6f2b028dd6aa5691314e52577a038336f0b0bb10cb0ba20dcd636a81e2465a22e0a90163332e0f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h934304ea162ca8060b24332943190d9b689d6020e9a2745bd1c8b62a6caf65572379b3dd90456a31795b5ccef86aee340e5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89635b1accfb1c5d09e09a68f8705e0bcfa04ef2eb2f777b3c56a91851483c10be5770f98c02a48b71123afad126240a28de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb68b1016dc0fc84d3baaf7d3e018b224b9c56513900da2a5d845ece9d28a38e5d4fd5ba95d827912dabd45c868ede1e002bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54d5039da7eed28cbf43cb5ba5b460af50569489556f3b380148192e2d8b5b3f8ba5a629a576b9d0a7d6a604cb1170e48370;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaf8cbe336890d9d249a91f12efc1a65c5f78a26083e2c56059f4bea3198eb071ffc26f40abdaf588a0fbd53f0b2d77f5760;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55208713c32a9c83c7ddc409617d11bdd1ec5c178ac930d4a8538eab6218b73e4d90c6616648508c98dede79b57c58226a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2d563d9fdc9f6294dded18849640ec4ae65b2e55ebfc289f15807f4da912e4d617657528d7c2a7eb119cce0029ca51a9f80;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc7b8c61f37461e6f2490fa03dac7fb6b025e9d8f911180efe71b59f9c687b3c3159ab73ab04ce7068aad7545ddb8a6b0f4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h134ed718369c877cdb3f2ce970c4214648fe7c1d097f7003b6ed112a1bd348ab55b575300be39e757bf6531b7339233f049e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h975a820224e15e4f3a67f6dae673d4b4ea389352abddb079fa714e11946e29ae8177f2ad3023ed47a2a906b2b52a5d10430;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc781114be2e1a442cb521cde81626cacbbaf0e6d1d7fd2354c906e21a47e0a98ad184e2d82b9a6bdb5acf5b7f0c184f14dcf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d88a4c824adca893667a419206eef7c15f1be225b84036d828ccf84afa39c0573410d9390c5862f4aca3ea4d4415952c139;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde58a1b27fc37f6a62eea41260191c583775cce1582dd207fe8cbf7642a29723ef708fad0b5fc24a68885fc7df66085d9d81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bbec0639f0b4deeddd8cb0efc65d1ecfbca607a8add74d2ccf4b4f16e3533c3e20155364aec941a15a15209df2e2760e593;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb07be46a3b1a0152d4b59d8270df8ea9a9fcba2c412b9d0d13f4d128e7389412fd1bacdf901585da223c658a3ba57b92a990;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h154ab4379a736afcfa2021e6965f850b4bc026539b6e951e5ffcfaec1bb0c0c28cc489683b078b1acad5ed80c93eda6a05be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6020e7c145a028e2409beed971fc6a901cffe3b97fbc1aeb1bb524431d20f91c86604e71e7aa739e94c7ca2d0f6241999bed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had97c880e38b760ec55dcc9f3e88496ef16cd71dccc13321278a18329004715f38fec86a80abb47231481f2ddf11b9723890;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0e6adc2440b57e262a26ede5f52427cd7708c852998054cbcda988a73e416c836f89da7a2aac007ef9dd36b2142767ee14e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h286c7df80f8f738ee71613afe2111dc4d21ef26b1afd32d446c799e9d9ec76c155fad8aa40b1b706b2d7748636a721ea4c0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1244c6a8ff6290520201057c664d639e7fac5b53fb1f548468de4f7f6a6289f20d513f1ec9dd46dba8cce8a658edab6850e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fcda55c6e4b4f6053f57688e5ddc6bfb3eac40856537753c2f9c643492486a1193da1576bccb93ee184a9580bbe654abf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd34f8a6b605a700e5d8b05102d83228d1842c79779b9bd42ff3576a0aa6f52a59dc75c38295b5217377a5f0b2459ce929135;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h109282eda3bbdbbca15dac889a92d794fff837727a869b7572daa3d8585c7fbfe70006e87fe1eddd6ee04f9309d49f2441cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76ca5cb6255881062d5a31d7299fc2cc0c47cf8f0a266399d54640ab2338bf64abe81033c4cad40712949defc1aefa436c0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69010f7f57e56ea098632cb81a9ced73f1fc0cbf9f036edf58e369f4decdfd668ef72d625e5b551f557202dd40ca9045d07f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5e66f0ff50efadb6d9ed44702c3352a3414ab76a4b111535463e697a91969f626fc9c236d05448790468e1f5e240639371;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habb851f71e23c82e6d2e5af61941bbd3fedd3d137bc4ae3bbc716ef6adc2d460ecf812db83bda1ab3854bab1cb450808126e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h841f0d073d64231f32a3f1186afd6196519964efd201bef868ea61730bb24a9e3f5e2e36403e83fc240f39ff1a5685fadaec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a37445d306769a41fa078815565029c111ead015aabdb983f7280984c3a6d10fa67426f96f9c00e36c1681171d8a810917;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99ca13b321b3065bea394742f6bd69c29dcd20300821b14545304cb46fe18de2b795ec3ac754402c96c7298052f9fcfa9001;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h176daf2dd4ea1411901adfa05d165dcafacd6c31fcf7840cb7c26c6864b7babc4de3d54ad105f9d22e985dd6c0d0c9d6d360;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fddefa2e21df2d63aeed0f0ebfcf7a91cd46b719e34fac122f60d469c83faf1391efad8dffaa90fa9f17cd27a09fac5a5b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe1778c214bfe6224addcf7d129cb6fd871658e2838cb1396610231fd859f1d9d75febf9fe5091df1f8c07942b197bddb06e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f14f8ec17663cbffc71b00d3a2501e3810371d0d86661a32689a7615243de862b8c5e44fe6a8ba72e00edf4efa4cd0be97e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf95352b1002c8add8a499f73602f0bca1c0915d25ab67fb6ce1e2963c4a4b10dbdde57fd36ad8a60fc094da784ad788a45b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h504a8a233c018b6dd07ad60ff3a2d5867ca9ec2065e290c5eb59bb6c9e1693d4bb8ccc6a865569b6e1ecf2b8fd74ddb9815d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11e10ec62a1def32208d922dbcccafb35bafe1dafcea6c6b418e0ce9ea0e066bc7fbaa9879f4e9f5e8c119fa8f5bf58348c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcac48c55ff9d63b73d329be851c070ce31eb7095d30e37838b0a4a969bd83fe46a571b41ac4fbeb96e9b027e26e4c6705ca8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8efc36f3f890722d0d7e016babe3651fd6eda3e017995e6ba6e9ac15fabdfa31cc2043800ee845c6bb1cc8f91c6f622c65de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32a88b6770d431141e973b86527d8034e052a0efe563a40f73c13d3f24cf336bb0886ff3f19307bcb9fc484297c24d6d50ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h228506273c5bcc4afa7612c1cd7644ecb47299551354c4562729cbdc2ea6ed894d6cb0a6b2555090d19baa38346ac89321f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb272660a9bfee2e0831018d186eeb9eaff3e9d6e2861b993a0c629fc2661c4b9373b2dbaf920943061e8b972a1c5ee9d9706;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd242a765f89319f8b07e634923f318bc4cc2396947db0e919e8a476aafddf1a4632836ec161d24364a546b450c20104d020;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h821ab87336688baa2ff290e68c5eb4b8062d60ae18f14910cf2617e4f7767b9be62373da31ec6fd7cf7a2ddc9798674a1be1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h152e4c7679524300a16e84461b8dae4ee368aa3d93ba0caa75c72698a6450aeaaae440dc6aa0c40fd157ac6421c6de737471;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h688e475ea8cee87702ebeabe0d5c45c9fba4b7f1fd29b99f6b472efdb1741c3ccdd161ce26ac35f6393f3c7491207e80e717;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7432c1945894c21c8a48a6be9e637e4c529197293bba9c6eedb417fba426eec07767858dbbbc1041d50dd941fd36afef4843;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc90868c17b05c3a067c595cd75220cefd4a9b32a9ec83a7bc372f426429be2df9fc07c0c70318316a4c2c46f3aaeffd91528;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4c1ff956bfff7a39937788e414f8f35784c64f52c31eb9cfd20ddcce320c7ea57545c00b8e4f5849aab2a40a591a3629807;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5ba6fff90ca7d64138fd53d9688221de82e8763f81c17fad3a07e84040767fbcfe12f3a80e73fc7bc20749cb96a08568059;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2db622b637d8484b92d5e03bbbf9a85890565972a1002cf7c3b749ff998ba89b7553ac6efeebe69ebdd76c4c1cddf89b027f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49435a7bf0cd78ec152cf7c70c1e43ff09e4ab2d1a9bf09b1d07bcfb7e38e0434dd0661dd686af0c14d0d3eac54b43e78a63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a4c4ab85592acf130127294210e38cbaa334f2944ee5efd17675119e240cbec9344e0047d753e4693edd3dc3a570b4c95d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96a64ef302e4c676a002efb6ae0ccc104b475dae07cb91a689b4acb8088f7fb7cf6a1707efe8d79e648e649b21916a51fe7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h366d3b92f14f7beb49f35d9e5b24f2ad45cb086a992ee02ec2797619a891d678393d46752a26d57fa7b1421a81a311cbcb1d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc513c3b0c2322815c7c579a51f5e946dbe1a6b535231d36072ca4e5ce0090947059b6a058c152f50f8c05df745708d623bee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he15f3ccde840ab2fe5ba4cf9e2a81e6268e6c9c1e8bfaea9b2c372ac2db423720fd7d59e492695229e85f630682ea2785d21;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a4a103e44d4c38d1d859051c1dc90fed983ba7bc4fbe412c4a3b8e05e19fcfd178b080942279086f5fb85c4815739f2a4ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h302eda10c452d31c06a1a669688409e17a2ef1312d347c73fad49d8f1938df573d33402d74d06c0660aaa3ac5a3051890f36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25154932b811f2e42508c3c57296f9a06d69a38add537ba280872c8f742c0f6b2429e21af0dc448e590305597a2b0f879cc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf87c863c90444b789d2649c75cbf7c548667ffbb53f6f71823ba11b8df9292b9275eb9515dfa96f08f2882d5a5f861024871;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ae4ea9630cfcb8c9fefde241a719af74516413df66e42e84ae4ec03f76aeddbb6414e3d64a5387ab098ecc6abbb3729dc4e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc133abc6084803784311e7641c690124b09f99cf2eab0a3a4094c63bf49b730d9cc58a1f25be485cff22a09aed1453c3aab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b387a31e4019bda7dc3f26ba046d6167aa53ce3b671df010962ec43e0fec2eb457a115489e667667b49d7e30190e45c1d50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aec3391a09cff4639e71547740e629aa08d94afab5dd5f6df833a48ee64fb0ad3d7c14c255e1172b3990b53c1a6e7de8425;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0cba4a494512272bc27c02a339384fc9b107728fdce2da63ca923d885150759ad0d92547cdd2feef450fc86867259794255;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5f23ed06ab1e9edf00d2a41b678c0353f1408656cc6b2fd9bfe7148ed440c243c7a5445779815614ee9fe45982f42a3b6c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46caeffc20160cd2fdb5738bf6a24ba147d39fa1c4a4d90720014d66f26b275b07671afb2ca4e0db77b754adcbe420594194;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa9175443d5363aa581ce3d6d969c2507a91d61c31abe5af5c3f2fe562da7d0a29d0b9b85b3025311c46799b99446a602073;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e99dc0c9fc9f89a8d1b684899e535a65249935daf773efddf9f53c723cfdb2809bf233cd9a340190238225e34edeb9a4a05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f6d05800c33ee805092a4eac4704e73f84910388059cfe3ebdb133c514af7a2addab9c7e2a71063f2871f42c4b27b597171;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0e17c1937c94b991a73cd77b538b2914d2d4f75acc7474d33a5bb277cfb905963edd3564838cd3d4f6cc070d90de4632305;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61b2a1041538e8460c87692ca084df3a6ecfcf0f989c05535222b730ba31ba02aac2fffb25a72e0f89262e1edb2970d38167;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ef82fae1e15b72c84b0371ad7fdd30f0f658c8d68fbba960bb83df1a0a6ce92e267c3b897b0632f2928f9dbb1da5d7775f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf25144ee2d3f89bfbf77d8e4acc4da203fcfd5564bd8e39be24c0c1b5dd2b107b90ed524477d4b99a59870f3592f0264326a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0568a23601c10f7bb38f445b6a5166435b9d5c0130e6c74be0a391d4bdf6d31d3366f7a5fee446e60d6dcb5737e7f9d3f1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28f14a4af30d591418d91cd78e49152ebf29ef52836737281258ae633db2ea10bd7c2f4799732a2f3dfbc9166526938f92dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccde9196c980b906715afc68aeee6eba91639219847552cb52c9faad995a24ec79f3ed649d50d987c8ad711094eda8fc988c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75d2e4ee7b0540fc882808f2205f17fcb0ce1f0ed498628d10410258119b38d7b601b165b7d5c98961c28b56d8f66e0e23c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8a9f434fc1d3cfb3d4aeedb09d77880626e3608a76d6a9d19dd41a85b03a622b11745867535cbe2f9d2875032687de52b9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6723a984fd49bdc042a6e042eccacc071fa4badaebce7acaad0d4942ea7b32f82a92de86317a1c3f362d6cf8c7a279ed43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30e7a77f647931b6beb6f0c24848f099f77db5d9e499cd2a7824664e4353677a110b491ce1643d105431af324acf20bc7337;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fdff3fc4e17fe3e0d98c15cb37ca49f07ad44f5e07e87d0af6d8907c74b1e60902d4bf5a44af94781a17d88c007c627f54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a0788552cc8d4ecf60a0e0fd3e1ba32162f0d3b101c2ebf3e04d1ff22366f8707bcbaf55b5ea083ca31fa178ba9473e6876;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb73f02cc5e064de97b5e9687e34632da9f0deb52d2d548ec14075ed9ac947e561c3f812a55af18a987873a732bf4d52e4448;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h478f45988726feae83e29974042d443f6b3c64326136e5c1f9781ab0ed5a8fb0803e7071320e4438158dc2929ce9a31928d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93238398946aa403c480ac96cfa95d617491635df1e050e78cd905649b48e44e3da62905de42add32b0d696d77164f8b98ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b1c5a74cadbf4ebd1ea92f0aea4ce1e40105e2c15be77b4f0823eafb15675a14c2d9bfb222ec6c999ba27b684c77639bab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8b5b5dff7c9c3505ec94d667b00c1d7a97040d8271f24ec8eb6290fda439dfb72b783f559f1053aa68f08975715dc479ae0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0f049f58e823815e32d99fc6c10da26c22dd86bf016a8b55a8076a9f773c5c35e27a962c5510740095a1b89c336cb449b33;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5981f0e1bc642c9beb959110839d60fa5e0fcd6c6ba697654e83df315d16e4587da8ab58728ddb4b2d850141010ea9fc6881;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62adc5e5f1bce0c188d03dc39650eb1df38d252e3a7ce166e013e3ed76dd375d973a55e98b0fd3c8aeeaab3669cb25b4474b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf28781e71c1eccc4fa645338d41e90172f5856cbbe8150323895d42051c5ed6995bb50ed3bca4403501d266ffab2261bc6a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ba77bf4548f84cb1bb992dc016a3a13878557bb70f1d2bc9e2ce4b7f0953486e30e13284205ab209fafd8d618c9fbad9f9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55949c1881afcbfaea7401d25eb53f8ad3fedbd010ebee7800ffc0ae524565a628881f708d3c93f95755c2abebb6b077dde9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bcb9f58802803c264a00868fd498d982cbdc01357b01d8a6827b9886c8a1c483249185e038e7b71702e27cdb71ad1e3019b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h655e6ae56047951999ffcca0ad922a3ca4177a463f6cf3f9498bba15083a8ecc8de536d21b45cc870478a0089452bd94b092;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0c818814d4115428d0d3b1c85c71bab5b111e8285a4dff1211cc3d827532f9cb9faad2e9d23fb55f77f6f24ec4b1ade2cf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69dfa3b436418d2eeb544277fd99b74c56f15497fce1810c5f6904cb7a160722516dd6470d43358b5c2edeb3915871da02cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb597d9c7eeb44464b65e577129b85cdcf885d21272376ff33151b47b859d7e1275e05f93f337f79f4985171211b993db4abd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36f5eda89b9a8dad50c35d14c2fae88f519be6130aed7bb780690a6fdbfcbe5b4d6b5f68b3f357929c090a90dbadefb641a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40e35662163c427fa27d102fe74c19c4ad8e881cafebad37d5727de8c3140580799edb6874ffe37afcd13576728fc7cc5b9f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2398e02ee5815a4ecd489e055df5ae96d0f9781fdb88690aa740f83b8d5e2bd73e85d29680cf425313b1b550dcaf49d92180;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdcd506cc91b1aff9b1a562bd7accc5ad2aa14fa877dc6b663c4445b3e16bad2753703545af7da854165fff38de6f67e79e69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10ed5c014ff3e02d35ef5b4845029f47f21c538949c8c969bb8e73d238a85206b8de4bb8e3b9f3b9b014e67606cd7a692455;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90b4bee46215eb9dab67d585c9983d58e895591161f4be4865e3f53c42270e426c47bdd05a0ea911110f6c17442451d5f6c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69f2440793ab03fe3071a1e52ef2c6c1192182c632ffb2451b441e33ef3798faeb1c9071d021dce3ca62ebb589dabb7f582;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he97bbaa21ff2a5f289ec768f30d2e41c838fdb9fdb480d47ca969f10bb791e82c63aeb4d3d045a35bf4f1e46a9082be4b892;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cd1a0b22511377784ba464a8ee26ea6bd7ffc06b973cd3f971c56fdaefc6bb58934b880d083b914e892ee6fbcb24021699b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14c44d06e5679819eaf464e32bd177c71213eb8fd7074ae824eca53081c3a9a69319f7f38842621592f3ab8fb0a35f1d7aab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8578b6bb295cdf28d83ca9956879b543cf03a8b64c99526a7207b9d2129629d06bf3c50aba027c227610b0028b6c475d031;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ff46f9c59002d5fbc8c58fc397c616bbc0036647be4e3f6f7bc709ce801fc9d17d318649e4882f47ce6d7b0bff035ce5c15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67ff341daf227e8fc5ef6bbb4ae1a04257fbbdf63c696879f1f33de7d899a5173ea26c2581ae2011462c3573a1a6257ed972;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13b97d5f116e148e702618afff3e34ced273f92d82059d53ae0b375dcdb419608fbf3a70a30f1390b43585a825fab66852a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1b61176489825ffb517a47f37b89233d679f21ae5bc00c6d5c2103e769906fe52a34d6e8860754dea70774f556ead682429;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60b18cd2b6d99a6459b92dd9fce1bce7dd4ec1d3fa45dc3dfe3e10d3f4b8061ba22f5c08e56812d50ef633536980571940cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521745b007d14c99b6a8b7f631df4382ea859c0533387a875af9f3af3a10c022f2a9d99bb3826ee18566c1b11fb8b466bac7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec1682ca71b767c3395e3079baae5f0331450b30598e50270bf8c931e16ed7b8185d2b22236909f76e94e5de130e38e39024;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26497f8aa6025feff69d473505e7c040a68907727ed5385ed726b891e68e9c96aa7e412ff5c4d2111a8850d6a6df96a49e9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bd6bcbcf0e857ef3e0241cb9aee9033199e76f08ad25472fb98f3255aa11fe58f9a8a8c7debf6b6613a0e6fe1ccdc356c6a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd06b156e661cd526ec3f7d08cda08881c83f3c3869e06ebac748806422c1bda18fbd24fcdc0ca09cbb5a71cefc17516edcf4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a7b4abb835b0b154e9ba9d71fbad7741b27f6353a98c59da9c4cb6e2399b4038584a765b87ec4dc9f4d851ee4989919411e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8f40d57ac161e7d7c0f4ff29285663ea04e1a58f09e5868b579f0c3a6f568831d72f64a3170841766c259dd4a4e16fd81ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8923473138be1a3843ef49cdda23c8960be6487b305801fea195e07f260b75377c47c836967c9e4333e035d6b4d74ccf992a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42fdad1cd6d46d77cb4a271be04fce41a16f136b800047cee3a0f0dc45b5e5330d046717abd2ea966c3a17f87bb5d411bb79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdda6a0cc723c54640e8dbbf608511a1c634cc49b7baad289052331599d26fc79bdf74e0c4815bf3d538dfe723a6e1b9754db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87bde34ebee839172d58969bfc5e1b1eb6525a8d342ebee9bf65fbe3ece1e008a172bb2fc52a3053673f98e10dd6b2c2b044;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ba3c3d48cfd8b3e3eaf405e7146aec8f2bc419beca921089b2239e21f3c010bc094fe55d22aa6b6b78f698f87af5423fa34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he12ad63494e5160e083f363c0f83272422d5e35590a31a58325616dd567f88d655be936841bc5c9abeff3ffedee5325e9f02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55f96e57950ed3f9413f7108ca59895131ee36537b9543b91b6d8c8effaff137d7f945bbaaf18b72453ad7f49670da0ee10c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31b34501223e973a2b16c08fdcc19905d0d96f06d05014807be26cecde0c1e2715cd6aa107f1dc7f952be718555a40002fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82f0b5bd880d35bcec7b0c316715dd79b97041ba716b3b5ab72faafcd8c2c3bff910ff06f666a3381fb866990630246b7c22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3aa5246c38a9ca301cd49d2d998a19f2d2d7465530e95639a756182a373f0201f0f86f0cbd096484aed3743a82617c9276f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cbe96e6cfb18b851baf0252116fe5a564ff15d4ee7c9d650cb22ee9a9d4b59fa4615f5fbefd2ec21a4ee61e2f1a9fc6f93f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h331675deebaa2697439e61efbaeff2796249626f93bf26683766323a6955dd467b0a376392163a0c944fb3dcebd690a2cdf8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88cf178dff8db49853fa2467d4ddd72ded36cedc1050958608b1f638011bda8e101012eaf16193f6b50decb6435fdd28bf93;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81afce095555b17f73d09a07baf0e67d39f6817fcf4aad12aba1f9eb06ab2f0f7929615bea30a68d7dd7d81935b2a66160eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23a7001abb072efee0580cb945be59b9152b619f71beb2b3128489fbabfa933c39d6611b8b76d0fadcb6f981495a1a7d0665;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b04310907263a70c5a4c157f0e1a696bb3e14a2b9119e2132e7167c24f6c5b50a54c959777b1f024c5348c7439b20061377;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7922d0861b4ce1648f9607c683e2a9db0291c00c64dfe997c73fae8515c18aae3ee78ae4c580dc5ad5dc1208fa47c40611f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcec0633b8c0680e6b0cb97cf8a52df42dfa9449564ca1e54597dd7aad3f9979747966cb63172e73b50e69a99689b91610c02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64b79f2e46395ddf1e2869c60c0d2cc82b98dcfeafdc8f2034ceec85dfb3b3791ba42ed9b1373e1bfa5b04e0c666ba89f699;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h902f1d715141a6ff69ff42049b80e6193a43dab3bdd1fc39fcb1e54cd97a2c40c64f5464e0dcabfcedf1981d0e55395057ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb618bc1fd9930b4b475634a2ec905070545eeb139690b66523ed48195014c1ca99b295d1a84bf851416e8cd30bf21ead3a8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd02da32993b9f3f05a2cf8192faf5da502213299a41b38ca59552115031f7fd8dc47ea4ab58392fd8072f0958345e1a60f36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83d6f758a97b0dba8bf36211af91321869a1720bf99157e34ce67843c1cf09de2b4b2e8c8c9159878cfc780499728133f0f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfd95aecedae209f63a9f7a0f5b85be380d86385e354aba9df67a796be6427b7adab352ba24116f86c7ac154951c2e518a86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4eefd8752cdab7d2ab6ae90372dbc2a37aa91b7ca3f921e719749f963657b9aa644f6b50b6082e7103906bdda6dd14b0cf4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9b8f56a0700a6f7d0fad02db7d37fc0ca06de3956d39185d3ace9a23fedad5e158802bd9b4694985b13b8a97361fc2afb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97e5183ae60386951f5eb860408ffbc01c633ebab7821eb308e9cac23633891b442ab590f43ba71819580efe067cd164a5aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5f1f0903c0bed041ce85fa3dccdf4bd5466c63fa069afaa5a191f8c0224e8bca389279e4496ef185d771b2712405363b947;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fb05be7bb7fdc02c3dfc8befe7dc2ef8fb6330874c73c42e3e4b21fa30daa4090be4358698e74cc2be315959d8c0e9820ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c6104b7f9aacf81fdb1a1798950ad94eac99f87ef7f7b5f8540613cdf717f661cbd256f528194b4aa6510713f96cca6c636;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb419a34c928508b9c27132471d9e2b126a574d954f2dcc7d82b9a767466acbca6e06c11153adcfea4d01666a5f8ef62f3ad6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b5fe90b8a2e77166afd1b06428adc2ce97e4f13b9b09fb2cdb7a70807f5622499dbed21ccb47e462e0abdc0f3ec5e25e62d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75389ea64bf67b9caac5eae617c6829f769ef6ce7b7a7c34fc3fc8acd80abf3b94f44cc4d37becaf506a7e90d503c9a1d836;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb70af49f1a0ec7a34ae8a87c15a493db561727f92a90e05133b0279d244c4679ce59c60f04de850b5eea375bc65b8bf10be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda278a71a54bdb9805b149f0f2aad87360ec06eca86223f887a59aadedd6f982ae360e40318f9c8c9bd9ebca3c29619f4af0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d28b93686217f56145355171199c71c2b0f338db29620fcab2b10b6d1ca7af43cb79eb50b1f8f6c08bac2bfcd21f2920bac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3773ba2d1749926657a2f1c8909c7622dcc9f42aaaab9c35252c71e424bea7ff12a9ed5d9c3c25ba5428474a4ef5e2fdb4d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1e09e307c8c2d9a6e29efde9f6fd0278c0a875ae89a3d0faaf103361fcc3fadc5226aec3a6a85c38f2f059833657986f372;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h271e9086b66efc3ee85bdbb93f5b11c56f06893068c78df38fee42e3859274faddd95d9e0a93cf2ff218904c7b6bc8876f48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfd01f3f9d6a02434f4e1031c1b7133c4ee96e27851e4e02dd2b756614d2106fb69da1bed6038f220be59fd5349be6f477de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h720c14201d226c6183b560439ff8e7b29546e7dfc3eb2c219d30dbae5ba872e378ecf8202436aa1e2be5eea7687c5cd14101;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed946278a4fcc2fbbfccc923c2dde52e79e8294f5d99cb3a1bc8389a45f622d38eb3ba592272bc858868493073cfbcd500e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha36d33152cf28c1be3ae74fced860e016d69180520828777446b50a8620c440d1a3cd5610bdb5b4e09f37ee04b21fe251c81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7594fde62b4eb53df17b6ca66c3e510a784bf48732e0700e0124ff84952e291943536a8b6e94b60244dc9b0b705125180817;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf681f1c18c50107f23b71c9258076a76a9030d68d41f3f2d53e792c4714c115c7326795656a0a193165d42978b652ecdcfe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6674e5be1e6e96efc9d5f8ed007ec1a8a38455c8c333163880c2b61e0ababc4fa170d3d2845ff36ba4308a23dece2b6a79bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2412e0d8934eca930e746447b1d4d6848f0dbe5cd125eb64febeaf5a60505ebae64343f1f7314135a126d73ed3343455c75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69ccf528e76f5ce498c5b8953b4050c4b468eb3535d3ff268ecee2c3e435e70240428d64b70a14bd03fed0b69159d7ffb59c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6e9f7e1554505bc3a71806a3ee26644792e1d84903ceef856e5184698645314659283229ec4fe491a0f3368f13e24010d32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84468d90a54bb38f500556d5176ca710a12422f7327d1217b61ff299ae65fc862bc7a530b4a545b97720130402fb35bf650b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc44e366aa13890cc8afec6bfee23edcfd874476cacc730d1e22f23416bd42b8b141bec9418c2183534f99008d8e7c5f4f9c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64b97bdd0d3247c45265b2c71294b4b4db4a61957875b962663dffad9a3f893d6534042e484a8e933a85122d6795a4788d97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45a5195dcaa00d99de5c1637f201de8b2542f0b75da1cdbbf29b4bee0543b5e4b481901758087b3e930cdaa764a055cbd717;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d02534cd043346a06907419a92fb98d007e1fc7ed4baeeac8b3eab44059ac13020841a8e2af5cf710b127d76ebd52e125ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc155159644ef02811369c09e36d346cf7ae9e495c16f45ed813445585b9e0af8a25d0c4a4e67ba0df10514347a21693f89d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a0479fbadf758853e755278473fdfb56e277b56f4b2652097c1f3d36b96d164863047be848c7c4465420a7e06bf78434835;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3aacdbeaa18265cb59223082055dcedaf1ae1bed8942748364864eb3c1c6fb286bb4b6ccb016feed7051e70706146d19ab94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8b9dd649cb2fdd94854da62772ade47f5118dabdc38d1f2514c7b2a1493fab6827442a076a7509195560d9bd91d5a25f0ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf952eabba96ae29953420d546e0246c6e2ff9ee7af6d093def5ae800d268875fb086a993d6699c5d2020014228772c03181a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99b7ce0301423e8e4af1dfad251f1d6ac7c7896033486f09031eb23bee5e0d859ae93447b63a4fed19e3026f00cec2ec5fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbec1114810ae55f0da010c78cd6a94a2561bf9e3b5ad11a2b69869cc9cc49f6de4ad6b0adde937bc34321cdbfe6b1cbe11e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb313ec85598cfb74ff2a81570213f517f00502156a3f32881c1b91478f6aa3c4e9a5eca92e3b90e978c38f1a9b4c0a46f007;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f381fe4649f67a88fcf70d042077cdf4ddb1eb31e20ede99f1a5746277d9d73fef068a03c71adbc969dd07dae57c9679834;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd099b668dd52608646747620d4228490939eb50c4ad9f8029c87f3b60f7068f4c926e0a813970fa64d76b865a8747207db2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a9a3b123778f2e79f8b86e7b3fcd108e00ced2cc6b1e10071a7b2483e7c8a56d16d4abc9c9899623a28ee38855b5f2788e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ba4c51dc8d27ad7edb933fd07aadf5ac6c98f7de40e3ad3293c8bdcdca903c0ccc0488089b71816550ab9965ff3296cc263;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6609f55b9cb687b87347f007e882c49f44174ea5845a062c7fe0ba14e117c37959e847cf0f9036e09d8a07b9981599171db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36641d55521d49fe543c6772703dd1ff47dc0229eacb5058e80ee27d4cdc7ead1d814712bbea24ccd3ff51cf53da11962338;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe9fd90efb32cd4b6e354cc63304fb5ddceee7f43ee3e613400dc16a0efc39dc860e5f100adbe9616452dabdebb3e388022d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d82084ef6d25a82742ad24468fb53a0050af60e6f18ee84ebd5c2b1a64a50631483de4270cd99dcbf31a1b90af90725c55a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf32d8fcf61b3ed1a114e5f992ae2f57aca44685d78c64f59fc45c627276f0b113bc1d187d3c03bde71e0c67bc3651ab8e16c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2488842cb62c460072658d856b67c76c7fe59fb3eb169b3685f5c106cbdafd533e891bfcb20492875af42e1c90347e75ee74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2d1da7f1b030b51b36e2404bc8199748691dd2452dec9f233f727b0ed351de8d1c4ee84c4d21921eae4467a52f864d2eb74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73b303925bce95bad8e45c65242205d42cb795554716e27911a835590ffb1fc52c04719c017aaa0ce1840dea1ca63293b203;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3a7fdbb628640f741a6b324ff0ef23e99c0c3a414871dda93ab7fa14bff187bbdcb1b87ddbebe2306f30df18d1cc16ac75e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac0e715aaa63b804a6fbe18d040b613a52b2979db2dbf4ac163f4d5865905dcb196c34edf26ed257ec678872995d2fbce810;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3ec829f153aaca6be7c8875d36048027a457371a14bea8af2847ebf647890a57a1f29f8baf31af69b5bb4f6ae0e4c2f50fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc13aa050506276ecbee0d0bc20c4d47cdf956318f53dad29e1863f25b088b095f592c5be3236ee3665e778e8159dfa9de4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbd63458a3c90a1c72c8efc64c01a7cbf980a3afc1d994a801242e5fce7a3c97e0434a54fc8f6359595da7c823f5083a625c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8321b44005d7b8152b68a90319ab847038e6109e6b042f24d95b0b8f1bbb2032d182134634309ed1c20dc9674e5e1a35ad1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h844e2e31a0f178c0cdc10ced8845cbda6402391adb09aacf4fa9c8cbcd769379e84034aaed9fdd3f37ce2f0beeacd9a1adf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8af3978933bc2849a853d8cae139b2858b86eedbd2dd88e383dde39fd8d462cf9913a731524ee13193b3879c7690fcc754d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h262292517963a3bdb85b5610dda7f42e34bf0231795b9ad8cb343d8ef88db1dfb85945ba8d3c897c748a006a755b68fa1859;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85834a040ee384dc6c031740fe58ac63823da6ba6cc8af6fa93c8c477f93ae4e430b297a3a6f248415da8de95362c376c509;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9a3baca91bc5342594f779dc4a3fd8a61e8d5da9ba0fdc0d31ff2b9f097304aa6901c14cec395ececec97717ebd89b353b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccb4c56055f39a7c624e2899e3a29f3aee80de35806c62c10e33070f2bfd9316739f1a5fdb889b0fb0eff0aab14329c62f3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c85bc3c66dfa99981188bcfa387133763adaf4da8cb7d4e95a776ddeba2fc6e12fc6650f81c9b77c4a9f354eace45c8dae9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce2bdcaf17b22cd6ed15d3886c1db503e54c0858e2cc804bfa3a7f10290376120c3192766100155176ad85408ac778665878;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f0669d3fda81d35c7ac272956e42b52a1a25348181e62431cf161b5426f618d1da8680bdfc8c5a63231ae8a619e0665612a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73f9ce0e2ffe6ff8f490c3388e5a4666c34eafb9f2f84bb174db19ae820bbaab0c9e208c1dcdcc772b8d19f9292a3fe8c8b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6169a706ba0153d7509df341493912fc272e96b023d36736d585c8fa4e5620d86ab3db37adf08e71f12f4fcff75fd234919;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74d3a4dd99d988832871eb8c43f6eb9650d2fba767a4e63d8877b5a04434551069b52897c27cf752379d76d0279d61627931;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h594d8411164a0b1d8208234d8440b32156de6a753886ef582edfce9edddbc0cf91fb813b4e3604a509586a6dd420807aced0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36f688d5677bc44798484ecb9046eb41b24d6d2becb6ddd544bb95c8452ee9b91cabc8f343000ccd4064eb12d29d681df388;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffea6e20ff930a67c07ba92dee5293042063739471c908700780c562063e268acb7025acaeb2b3a22b83bba59bc54440904c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7ae2aa0ea78b4d49050a945b08a1f3aedeec2ed4dc363dea66d270e1a7f0e7b7859416b02f6806b251e8fd17e2163c7f113;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h787bdce119f57eff7501d280866bd8545de9fb4a8c196b8ce1b7400c83a6443216bad002b06596f05f64c0abba50b029c3c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437cae925373420d866c7286e65e69b233494b56f59ee22438045085c662cab419bd0a8434389a1006a393b41d829c18b21b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3498ca4d6d7ebd1f9594beffe13e629b4260e155e4ac762c96488f04410e1e3a38bd081e72f1b597392d8681304cc18b834b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha69ca284316d933450215f2f955224b1db0fc05a56a6c87401ba2a7fc80daaa8d3c194ea8258ac178521cb8d0bfa22bb46f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ce7d462c729e7314e057959e9e7ca88e88af16903db7cab9074b0d1e340fd05781e67517e3042736eafe20d860c13db7f05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94d8498a36b96ff9888fe854a24f2d5d066ca7e46d1eee53a562dea89e14a1822797830b44d19a3756a2c74f6f3602f09644;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab0184f2b25b3d5cdc6efd88cd3f397a9365f6997609783c39c3991eb51c2af459c572e79762aa7286e45538bb6b50b23577;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38435eecc20ee0357da281d105384a053ff2b1c77f1d074429cbf7b848f4ba14c7c5e0232dbd15bf42f52172bf0a82f1def6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b4fc3a3bd27a6e9915bbd0fef337bdf282e810d8c699220ed49b4a0a1d92ee60bb246e36440318b4d779c3af8480289165d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d4d89531a2811641d537434c5d1395ed62c9269b262a34a0a0fed07d66bac0384e9769c9d96a52a5c55cca6f16f2beba751;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45dee3412786a06c4b7869d8ee3227e67f5cccdccfd88dc9084101500b7d6a371ffd9a75fb92620436acfb940a8f9018088b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h412d7a7afd01196dd6b4e68baa354ad0933e8970d3de9f91177d34218a604919818519074ead42f271b495f1419b41bd2dc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3678c973d81eac92c05a557ae65e8a1c3096e2bb048fbb3ee2ef90e3a6d07a0e9f2423cbfd1234dfd372100267b5dc93a410;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h236068c317b3e69ce2b26db966259235b25424ba6264edb8a6a6bc69f1656ebe0e43ff037b808776b984a209240c2b71f3d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf37f3cf296bd9cbafe786ac8b0f462a090e128e8b91da02b2e0e21c66131905828bfe14353ee5742d00891ab94ad50d4d64c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae9086902eaa98faf303463e85942b0b385eb0afdcbf93b0035367fbbf86e0ecdaa916f58baa610df070710612e599b0ae7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b1fbc4a991702d371f2018a5aa6f7a41c911a9f66b49711bcfb7a852743c4b64ef6b45abf36be59a2f8bcdb5cb990b2141c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6133859ab6be7a66c2b6aa877c86482ce64eab088a2f68481bb89de31f75c7e5d1584ea0b7d4a440c73e8dcaa51709cbc15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9247fff2eb31c2817be88d779e20525bc5cd193916d74eb0815df72cbf2d3aa01d6253b842d8d3ad88ca56612bed52335e9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cc3686d6b923315585b0773b4adf06a686c6a7adca73b2fc0118fa6d774f6768f377533d80071d424f62be62c7046e0a2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5b220e7c570b16d710a3b954d94591be45296efc1623865d7ce87bfa9c2fc1d2522ce6f5ac7a401fad7253fcf35c1944c28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a821f0466641dcc7bcc46784a839d02513d6c46845842132ca4901c37244f06643c43147f899f678cfd29581bdb846def45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc775e81b40f391d1c6b3d8a7d2fc091fae8c542afef790e0e928661679a36a6bbd38db7f77ce8401b97811b5e73cf7b818cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2e5c4f1cecc34be6db9fac9cde8b5f0c9ddb5d705cc2db9481f41cdf156cc43631cbf5dae501527da52e93ecb3875d9682a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4587768fb853f993a3ec318595644eae0fde791306da50b434e8ec02f0cfae61bbe279dccedd7788f790689f06893de103d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h897edd1f3cfaaaedd346aa5df5214059d4dddf41d9e81640a94cf81275cadb6636bb81f41e3c684c5169277176d0fb2ef536;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h355b1cee788320c35fe3ebf91b8a61465bad7eca72e303ed634addec142645ad74984b6293a6ed08dfb0b66bf8f5bd60a31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dc39bc473f52f21c40cba7ab60abd511653a4b0c3cb5ea0ea8ac734bf876204e65c943b28662f9e951c350d5dc8c0a34bff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d175aa7a72ac03a79f995db466e457812e03dd27b413b57ff0b3cc074aa63f89e4779b79823c6141b3900dcd306b9208d89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51ba19e78cac2638c24b2341a2a87a9d808547a199bdf2065c6b162e84a2a3f20cd59032418bc44efa770bf0e218eaf8f35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc8b9c561125ca0ea9ce0cf8bd2f2b6935e60b1b2beb6143a7b4240bfb4c0735b3ad712c71c2b4e80ae30217977942f08d3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9752d62284ca36d9809e35c5b51c3232055994ab39b9dadd9069ccdf6008be1acc4221f11e741447423ef5d1b1f7aefbe249;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h710113da2034394e99b1374902eab64b8eca20054da5aca27acbcdb29d84b52dd25007fa8d2ab5ef7ef54a2349bca93b344;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee3a564f78508d3c3fc745a7cdcd8d45a82b7e58e6f8f380ae575c959cf9cdb35cee6175a7dbeded939ee7b6d03b7d176e46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb947eb098164a8854853b686dbddd42a0b7a05a94ba788e658e5f95071d53fbc1016d5823b8292ec401d32e767190a7f88a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f7db62d48dc90e984334356c5a324f67a68be43c42a9c4912e191c2205dd81521d13147cc32ac74496a706fb286d2706277;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcafd8be09c3adfff113c162acf02dcfab5c8c87d4eb40b7317bfbe279d5a3207d77cae3c47eef7316353da0238f163d8db0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0433dab7e0eb87ff830a6e60a913f9ef7031d3196db3b24784101562c07ad7d714ece7eb70ccd3e695d45f46dcc3847ff3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a6096f2a6a2dec2d3b612c651b633780786641352ed3ba962dda5a655e78fde169b6b3684966f91ded6416864d885419a1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d8faa52e12efd285af1ccad01a39b8a5e26ad390c52a06be3ade7786013a9b2527b3a228a764c283b3cdea4a5d4fea38077;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e9b667822ba658f4dcd275aac2621853dafe201897499ef494ab1bdda0d79d202a1bea12b319e3d561832a2fdadf8dab73b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d62faa898917390773d83bdc0888cf888d2e322484e099c7f77fded4d48bd6f60f75031635c011ad7754e015a8097791aee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1a9931cd455b6d0cc7971750dd5c4da07d11986e5d82e2ded881327838812fddd40f9dc997b226388df946660439b708e8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe47e7ff9c3c0a10f3cbee43f515da9373954baa91d738c988fa2f047d5d05821f57db915c005477a0a50a0a2f1b7528a152;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69c1cceed9fd4c9065e52711983e31c8c1f17758955ea435a1273679566131a123d51e63f40b2fad7aba36277ab236f19dfc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25598168ce2bb4de5fb399d3db44d48558e84c8016029777b5495350764842b32a81f1d11fa2c2edd3cd412aa73998157e85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h166d123dc9a9d5e546bc8f8504eb0a32fa9b084c8a9aea89240c3b5b5246d48ba8846ec5de1f803a3f6587d5f3774501eb29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4b5822199ffb0cec6f97dd7bbf6c46ff6b5da6d7ad96771cc31f4d2bf1acd00bdc2ae549a387f78165569d43055cd51df70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdac5f6251a99aeb035286b044cbc395abb9b4efd7e126be09c13b758783c8f19fc3dbd569e60079ad98f1a570441b521687;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6f5efee3cc6affcfc52e14ce3715cfce0c98bc807ad031528af1d677145ccd4a7fbdfcdbd5e0a6977759bb0a55b6f00624b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he14acdb55a9e1a36d6e2f09c9d44c202897044ce27bfe267dff3a87bec4a543c3cbe3c3ed895b66e8ea2fcb428ed690313b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80fa68788bf213fc3bde0ea04f5b9004832aea9c934fdcb68c37101d9ba137ce4ea11b9ab7c39c78bbba4fbd68d361187378;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc518cd34358f1d8a3a85c673c7c5399e0b1db52113df04ff8325086930de00b75668ca2135787704c949f5cf0038eabc320;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc68c8160632725c761b4ca30159f2a34a5ee0f460768cf77a80a559e7f643832a1cdca05a4dced1454990dcd7d09be237235;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e89cf1b71c7d6ebd53af19e0328616281e6a38b98d389f61169d54af4cf669ddb51db569a0719141fd80c85c4798243f30e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b7234f2cc3b69dc21b0b600015baa6f8c5aef08a18233736aab3f60e92ab26ec42c0e09d5d7d7857ee7e7e76a9d985174b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f87a7dae8396cb63c23784d8d5589ad7844a77d87a6fa4d726f31e59c51d3451a14dc79203b4c7da1374cff1089923fb11b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he66d8787d55a177d9b52727ec93546914fe2c5f227c85a78223c9ab0565383e8875abf0ab37e11895845f6497c8e77189a5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h673f2229962a565fc93d4ca8134eb0f506c4eac933e7d640ceaeefcc5dc428a09bc06a4c6a7cc53cb0f9ecd6649ce608d606;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b2b11a9b0387878d61da6e03cf5250226a425f05bce93d6a00e8a577e01fd8b3af605d38ad8b92066aa522a1fbc770c0a84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6295cf34b7e58542c2bbe51c9db341a6a90539c4f8f7dd79d95564a7de383d3fcbb198d4873d231ecf14ecd42fe39f4412f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc42ca7a6ae4072cc654a9cb20f91086ca39998261dafbe2551fc8ee8413cdc2d5f3bf3eee5a6e0636a671dafe3dbe6548b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h846263de5461d38a6107bd51a5382811a4c8ccf44845ee57e0a0d9c2336d3556caa66a9cbbbbd47485b0aacb62e19ee5e7d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b89530f0282df724d8bd6c87409bd44b38190d319ac6bb5ffca983dad62a8e1ed9907dbf560031c8406dacd1dd4b79740ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5763fc94dd06ae07f5645fc47c8c52b4bb9605d5d152dc618d6ddf6d5ac10c04286d9cf3111365bebfec7ed59f7c4f028b8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8ab17ea46d5ffbd11cf6bec72a84b03a623e852acf2d34f8ed22d272668ba573781d267ccaee46f5a0c159de189f79217d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36e11139c6b9a690881a3f30805b2c53b4aec26cff32637a029ce04a40b6e2b70711d66389ce1c955efd463ef915c6cea0c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1108a85bbe0798fdfc4ddb1ceb1b93ea638c8634bae9a709ccfbdb51e158dd99629a8fa7ce25662f40e18fa3fbefb46378a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfa9533a74b688e87013125ebc18fb06b391d17a5114ddccecb952d9dbe46b1415c29b7a264f54dc0050c3e300af050909f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80aa6da8b47cf949d5b6e01b23628d65db2048bdcf0626c5b21138443ba749ede1546bbaf57239393deb60ef1a7cc1ec883;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3e5c842caab9bc8c8f3da591497b2411d2cbf9b53a960af940e51e4b0aac15dd6676346769e71c0eaa677fabca8019bf42e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67febc82766b8cc27a8cde748711fc99c43a3b327be576fd4814c7f803765807fca73165a8dddeec6a706ad2755fe21f2c34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc68b222d2924e5230b80496caa5f33eae2066b4cdff855d06b061e5eb7c7f091415770b79a32bbf193b02c6ec5ee681a0de9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9cde7f03526985d198717637d343addb46a394ef655017a9290760743a0f4c9ec7a60502a303ced4188b1c7c6b8e6145fed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha787e69aaf224bd4ca2ceb1e24a50c9219df68bf7caf80b951a548e8c565d6a43721f42c8c80a3972fd34f521b41719a04aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haaac53c3e1af096e47e98783e01077629e4a21ee8ec9ffb3c0cfb79f4e6f5be791ca8891d9ba0b738e3071a3632ac08eb8a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb293318a2ae832bec58f44d6a8cfb455f53819c42553cbd8a55026f7588c9bd3ee95d199bf23c4234e290ff1dae232cfddf0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc21160badfbdc6e162c0d92293fbe1078f26f48b22047899cdc2ebfc9e213e888322aa8b39ecce11e17ee893f0bd0fd3d9ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a2e6480c817e4201ee193fb22ee8431e13dd1123438531c06d27b98a0148a90ae785a5942864639c24ab77d296208687e65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9735b34234b8939d9a48009874e207f83252862bba7705f934dcbe1b711669ed12075954f1e68fb3b64df17b912507e5ca1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6c0c5def9b698be5300ef03294a1005afe8c385ec055ab55ade6c29ff6e602733993ba1cf41de57eafc75ef66ac6299874a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b306dc387c1e70650a3d1bf1d194859d748023f254192b3e127879303744033f43e5b3c76c5a413e3e2fda604bf1ba8e8c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cc7696397bab5e2d0954a016cdb0ce55981c72ba57edcaf04ee770613313c5293602b409e98a32d4eb8fc5d0e056f5a291c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cdd6b0a8790ef3b09b3e93c7ec0dc70263fff02b87f6023c48ad47b7618f2862603337c5509bb65fd2b92304295bbece83b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7ecb2fca7c09ba41459184015a824981ff6bdbdf2df5ec49826587324a81ea2a8a701569f0af6683a9e0ca92c9c65b9802a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaf7f14c63b0b162f4785c3098196659b7ab2f5cb5d7b4577cfca09c90ae72131cc2da4add0c07a1ccbe304da7ce5d74eab2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b3d00cc194813ae3c265f005cd51c07a7cf9628a0135f9c18390df39b502b83750fae744f8fd9a1fae465f210458ed6b26c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39ab93c0683ba06e819a0190ab096e9e6252c33b59b418b02924c215f805dcf015985157129e444fa5354b04cf4e27073a73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb15e70c87fe582d1a7d47afd68dadd8ad28a092a5ac8a459859a7ac0869557dd7488c838342e7d6d2618b419cbab99d37de1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe1f652bb2d1bc118ae3189cc29688da3887b90e133e57d30077601e0b5a33e241665997011e22c6c6438780ed9801feb1b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c85f641cedc1d1cf29537d629a8061846cc9f66ab110812cc91052bde450f9fe684f34c383f3929595994d2f013f729a08f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb56291a71bb9397247461fdf3aacbfac4b972f1dff65f891234b3ae1a6c82eb8972ce2487f81513d8c4b87ee78147818f54d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbe0c42c39ff13c7ec0af0baab2c30503ee57e0bf1a533a2eb30977a337eb841b62bc5ad76d7aaf43f2ee4d11cfe83954b64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fbde0c4315699024aa07b567cacc479e0003a32f6d10c5bc03bb740c14a2ec76b8c25f08aa253f81654379b8adfe2e49d42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd06f1e49643ce4b5cb0fd9cbf2552b3b7506f33eb254489b83574f54d370301f058ba387e66df0c3704093c71c872b6d9f51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51937c773d88d558e54cc4192a43ec83cee46145f37569a43d7b9f68c738e73fb1dc58bab696c6672e16750db366a0bce85a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h356a35b400ba035c46a1bacb086769383d14dbfca768fac2767fb18d98afbe21cad9d4ada5b60f2534eb7c89ff2430330c5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c7bdff8c159f11ac0ac1ce443796d264ea427bcc86d573be21a2deb929bce60c19d09a396d7d581630cdeb151567daa90a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cab7e764f7cb9f0b5955968400bc289d74061f9502a8374cb2b7246b1ed184e64cdca8802547ed742ee258d19fa0dccbc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ff21260a88580a32d87d058f99f51e7cf1f099a5568b250d98fa3eb03f10c6ad39d53e5aacf4c9b7d5d4f41ce3a83223be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf18d5350586f8f6eb627b70a43bdf3ac69585212a7cf3567548a67a179a603bada85a3217e0b4f1909419fc6c15ac32fa6f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb44afca204df96356025d703172758ea1bcdc3b2d59ad78d82bc8aeb126ce855349ab68f5831011533b91f18d0580421ce4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d240754a56a92940700dbf9e618eeb66a1e66f576639b73f7ce9618ea12fa03ff98b86d2f3f7ff15ddc6e1960e98fa5110c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5410efa238bea2599f77f112decb12c9ae5dc03cb916bd1b258c5add08859239b75c8481ff6a7a1958d830ca56d7b9f4840b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ba7b526f4cd38aec1651119817fddbd19cc3660c58a606214d22d6ebfa0c3cf086e2ae5691e6785b3168bce90d073774f4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d2d3691d883015bdb9e374381df28c8b5500577c88c539c7b3f5fecbbd335d8094b28052351cf469a7da7d5767971a58123;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e8068f61e3c439d273636772b9a3ce6369f281e59e3c8230119e795d2ceb93d6aa02c794fb8c6fae2bd0d1b300e4b79fa4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c1a0bd092d6c573ea5d2b325a04d23d74b4611a2917a0bfe718d1956a8acee8550fbfa46f1d733791a55e7362a98c887317;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4373ee7de9d65e5f313ba885914e844eb0fba3ff049c4dfac4b08f406b8d916bd90ee83d35f656556bd68b8a07573f346113;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb576353fa14184155e5a85caafde139e5eaa7f8bcde7b93fbefc034677d5424b5f184096285e6d635cf04a655c98a4a84793;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf73178f0d4cfd3486399b857d81c9471a4267aacd45bbe0f7421dfbb47721fc57067a67beed967fb42e622ab78806885fd8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddd3a1066024b3d75fc9b6f2d372cf03afc507cfee6902ff0d0b5b6fa7e10acacd4d5d2a474287a4412b72dfa6b2a47dc906;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h149690e30bd07dba0eda4e17ad52590fbceb5a76fca346de0677c8321bf3919030c0db3fd8157be5c50f5ecd7f2831e099b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc70eaeb660d678b77e4f35235a5b7b69a71be7713b30c449e5e590ec403edce1713ad4bef4b1a9c81632ab7050d6ed0a3c1e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8e385afecca996ff33a88019a5d8f0dd9c25431e8686691a8a6ae73c7f4636cdb100d28efe05226155933d5932d36b6c974;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49086f6ceb57ebdb22064979c4bceb99e697714bf3514147e7d06ecfb8e486dd92c535bae3fbd1567f0a1cbcdc54b20affb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha78e3f0ff79a5c57c1fa316294c2f7278e3b05c71e4b2820b10aed38d36b2d20726decb9aac31ccb39a5ef7ddfe11977313;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63b97261b9aa127ad5ba4d5c8b8ea2e21c6dc081eb78f2c6aef5c5bf4288ac42ce624ca449fd29f2eb9c56e1a789fad24b8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5429c2611d13db1cc7d277b62d9260b6a744faf1c1e555da2583d365d6eddbf8129925f03d67927e62fd3be4629c9b05a4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e37b55bead1388719897208bd1b6ba8b1fb87e8541bf2b34a714df6a1a9f2d44a1dbcfc9db2ac1f1b48a1861363a1886329;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62f3f9cee347704a04121bea176f49c8d838408fea92f000653c2e0113b6979a60d5fec9f2d8fc25fa597b25fbf32b00841f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5fa547734549d1b0555c3a7c32e3161418c371896cd929ed3b36b50b25e643eb29712db86161a52436596814d785f856df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h452ddfee3657682f97eaf041274e4739535abe13a574ffa1b3e74dd78d3ac3cd2f53704eb2817596c20b8e0250bb9a010f81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd632fe46c2c5647ec4a7a303c6c6e36635842d2ae6ffe58d1a3f9bf6a7d63cd85627b07ea13c1f1d7805b8dc6600809287f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haca54b3b6119b511a2c361c3f3fd5f0a9b71c0dec8a507da35ddd2f21cba3b0e87e02aad1ed6ef6de987819b4581b4e6000c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52ee9cf07bcb4cc1d8ec7ecd566fb5a1d8b5a157d77560119aad98a5ff4e8948236f19f53302855b7a14249860a0634773b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haead8c4d48165c996fd2b00347cc2de4b54e9ad877bfe5e3c7d3a779ea3ac179567cbef22f27f8f68415a70a0337dff0c4d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2f1b58b1abe1948ab3ff6c3c7c9a694079b417e3c889b10eb1662f2d9a1b64f07e89fe8629feeeb9dff6322f40351ef7239;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75cd3bd1ee15cac1403ccc1465ce7fdfeedf2e8d9f304141ae21400014fc714f4a48ffbc11f6c8c675d2ec5ae944fdf9d5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h755e74fd6095ab8b03cda046e353446652c29da25bc3a2050b03074af90d3e82e45170f5782d744c8cbfad7f3cb6915f9f89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf44caff83d19e5ca6f1b3c169aa1e13db264f0e2f24be229fd0162bd4a2d868b0e098a4a73dc06bf16eec85a8e905a4e9159;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe0b97090211f7fdb95c7795f16290682acbba662b2579ddd97e7d91a8f8cf1ab0e639bb3930977921aa7b6f3c0e5ad9f788;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32f59045c881c7dc07bbb3aef0064ed05cb40e999919d3a634651bc68885cdb48b2b0077ade02669183a85c01b9594848bad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dc8b5237a69e75426b3006b55f507ee712edcac726c8397bed3459cde68741aea0b8d390d2931506bd52cf2c7d32ec5ddee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27fc6fe4fbeee9a5f4a89bfe89b841f2030734e2a40ca0bdca6e02ce8b40c55f0292191d1b4dd505e75f4b003253af0a395;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h455a2b917eb7c914ea56861ae2b0dfa1d0384eff59d80f69cb72b027fdf75a47601926f29eee49c6c00cdab9cd385e3d1253;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a53240c11df8211ad8e8ee327ed4e51b83096ec0e39c2703ed0b93bb9c04b07ef89fa9eca254baaf94401032ebe8a4350fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbbb6e8df5f662ff7742e3fe28a0b5aae3c68ff3905f145eec75555c23b930d674955d1466561bfc1400873e08e2a7c1a67d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb58d71ae6cc409655a6df80e2bc41f39a64b07eed50003550e2abb1412f4fa0de9560506fa80f645f22b02aa08089c96dac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd961f96554ede20bd982c2b3f8609c95e574e922d2d5395ce2d32a20527d559921161f5a9b6fa2275a604248275b8e212356;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65f771e30e4f95667878c42d29fb6593ff027ff752bceecef2bc4618159d0bfc1dae0fd491b9e42476ebb53465f9d797aff2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8066b0fbb33462246bb90abd74057016949469ebf1e706600a39cff288428be23eac7837df3e8d6efaa0a008e1046e02c452;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5205f178f39ffd9771bd2516c305952cdf1aa89b8100edc0e63fa7212dd0c4f7d7da99c420ff438d3264669c996d380ad981;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b5cf65b1df652a286f21ffb01fefd62329f40b011cf343d4fd37006fd2f55d88fb454dce86effcce87faa07b27cf15d0af8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h819636add3365c479dc7d7b53f5ab9d74f1490223ca7201fc340dded592b3f5f129e4dc5c4fd786d98168c01f3db76b90fc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h315ab616b202feb392038fadfa1a260ee1f6b8607c741b3990a96c9b19fb91f14aad1833bb533e15d1457fdc1fbc87eedf36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecaee2b60076dabb39d46095e30f47bc5219fbeae9040a000be81e36a762a80e4de41fad281150b56594bdc85d799515344f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4da7933b8434134fa57878f00fe4bdad4bf0f5e3ab3cd52ee47e57ece698a3b96f7091981a3b4b26e3051610752b8bf4e1ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h261c3e5e9fcb92e3450cb06ca2e0a418df24d53fa05e7358c9e2326c12858b809829b241b49350b130ab6376d3e1ca797301;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h317a3d53ef176afe550136f457fd3ef86d39e9d6d4dd906c522966fd6f2c2227924d94422a94e948170a11d26e87263751fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h785fb99891336f6d594f8e20994cb42f2564d364f03516ec03f9f813e22149e7b1d6e478aabfe8e53251bc718779365c9e5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79133aa16ae29fe488cf8b4e7131a2e14d6c21cde409697fa9389a7deec5e92c7b0db49f155bcc9499a162439abd29888912;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc916326ce2c66a2114422ba0adc59b665a6d21a0abe5d0d54fe43b9328e873c8a3cc273a79b7d7659fc3d4f2dce42618f713;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d1ac7f05551ae11827cd81a9481371bf1ccbac63dd2fe68ae895eed3cea226ec7e3d07ae35ce8210ca57143254e6d18117e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf534161a0e67cfece10fb804670bffbb324a19490bcfd9a073fb2d637ce006f0dc61e7e807b5f1c58ccb257fddd4cb03422b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccd6ce948f37a73b9406ff3178a0fc6ab9e2250ca5ff63ed4cb2612613a7c677cb5d09693b1bdd44ad374ca1976336209ffe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8defd819388da21407abf9a68ac8ca3d81e392f0003fd849b53a6429c4e1114915a1f9306434eada89c134ce27e88554df8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ca7477ae04adddade28da5bec7bb947279c5d3fd05cbf8d14176d11f82aa476209fde975733d01996ac0bc76140900a1488;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec8a35eab97b0f3443014f6efe1d28771b535b079da10d9e59956e7ee99c89be15314c735e2150e25b3ba3c7ea2d3ab3d6f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h741f13d3f37ffc91624040650eaac93046c0a7b581d6cdf0c97d6ba448a8f4b5258e791386a2e1a846f7fa4362d77bab389f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1306f2d7692d721e9a3f4cae86b56018695e7778060b3f9ca8fc61028e9727b6527cda1730abc8853eb162e7eaf01ee49811;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3768d96425e1e59126d3a128fcbb1ee78aecfb29a4171ea5331af0586e03ab276c9394474df0714b37d5cc1f0efb50ca7a87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83dc416cb00487c4ee7825ab94f1d9fc6d229c4de056b16d1636b6f1a63f1c2f3c82541bdc0cf3092316e37707c457867eb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f453d20e1223d83157a9595515abf04d26a07567239843ffe6c69c086442a92f4e85ae96462d9ccb1b24b7c416b79b9b913;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ebfed4f7507b41f000e78d45b8bf0c7d83143ca3f023e8977ae1e1a95b1cc04aa5ec3320d3bbb36f171828c1905535f82e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefddd2cc55914a10127a791ec016644cf679fb7fb56bfd82ae649447292557ee6263d2e7e21dd6c8cd98c3e8a9b40ab66012;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa834589ea90f091ee154f9ece291f15a2e6ae6274d06938aef39e88f38885aca20a868d8d45a30a34d545091545af71fc87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd5888b0962618f5db959a6d322c24218446d111020219b7622d14f5c06996e3a91681587d5c1a3f056a101ccd55893cda7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17902eda91ac6ca130ce92cb344c8335245c8f44a4598eb81da350e30edeb9337aefe0334ec5508e8056a33fbe05ace97fac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48fef4fb2048e8e3e9bdc97dd549310e73ecfe8035b2ef80ebe1a5080cc017e28a0a0b02ba4784254fe14fd3c8af89875ffb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60b0d09f6d02af3a6acde10716bb7310678ed93705fb4de6f8b99f57623ab7af0404fbdbe5f6c38cf0bcc478f3903551d607;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h162bbdd76870a18678eb2731b2290469a26036306918c62fa799da4e37d3795780f1373a769c58412d51602840080389d2d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28a5e75850ed8d6b5e5a016a03ffd5c615c05d810ffc3d35e7dd3ad9abe2c695fcc2f038a22ea4a6f8b196fadf20126440b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec8417cfdbb5cabc4dc2fcbd0065ff540d0ee93ba7ca958ce7fcb3b31347bdd13c27091f4197c54e24f93a48fa92f46e326;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h206253692a841b4484d119542431207b06f5dff3b0350f2dfe09e8e98de9a1de8f0c08d3874da441897396820fd6729a48cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90cb3983dbb6117bd70bfaa7282882f8e635d1f2f83b1812294f52127cbaee6de9d2920158c41fdef84d7e7475c852be477c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18bbb6525d7b52454d2f7f3dbd2e2e56e909791ec22b86a93d89345f3579abb5ae47f603dbf8c090f7907fa6a0ee9e497dc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fa18027c22363fbf24cd578b11ce10edeee8c0bc09ce0952f3e0d5a8803e59f8c29f9f474349b4d09d6121a8a6544bee3d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c1887a3e7290de089d905d3af1e5ab2c1babc8d27bf749edff7120f7decc5c93a2d7b5ebdc5aac1a309a54cf83248f2a522;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h433a51d69781716c048e226807f8c453b063e65024dc605e750b139cef933a9a06baed2202b16a4ddb5873e9c9e6e9246864;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd32ef09d1a93f1f1fbcc18cd75cfb140bc8cb998c72455e2bf5aad374a5ad5041c96126aeca3332f05b55837fbb4beeefca6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h235f9013e017b16f3a0649c13d58cb86b8ec6a46ad416b020b7abefc25bdfd8ab19b105d7ebaf837eb5945ae9efc61c7140b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5081ec1a312be2bcaf7f814d05fe50ebc89701ef4769454c0971d99f98254b9b303b7ac04935b97f8ef7659514a612328635;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf878da8180a1991a8d594d725e5c019e0e6584b0fade44f3830aa018029da5efb1cb076234125e077a15c07bf22d79321f59;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h483c479f8f6d46b72d9003e22e0cffcbb36dfd453056fb3c2f71e79762eb659d0856cd2c4b4da474c26a2b52b464b0d304a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he355fd297f124dc84654aad39b2d7912d789329923ac7b68fe3b9ef2ea000e034f0feee86b7fc84b437b3ceb09b04dba7f50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0373d200344203eeae8849699fa616016403b651a2facc7bee384195ca2c2f73fe5e5875fc59b42adbc2be34b2417339445;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd58c21df2aa9f49599613d045230ac4b7373c2d2fc44e1730a4232a364356489f8ce1ba0b06c4b65e7c7ddeb239100ebdb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36639ceae26c58fb265f9d9b49c06464b512ee9a188df0532cc669e6243173af3f039b2710a0981c6b7b5dd6c02b33e063fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f064dbde80e03615d187f5459ac1efd6bf19301032962d8770a9ba81d05e1946d4694778791bee04fc9aa7b7e15f36db821;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb499c244359ac15957c569b61f819273df69cd34d4819be8ccc025af65a68c45241a75feebe02a9d4fdce5e5c21a49bc8665;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f9b5c01032029bf0d9017a03aa1033f2e63d541f39bdc6987d6e197e65f19a317b09a3a70592ceb0f4f70a669bfb68e4aa7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9d246810a7113e0af35edbc1fad0e64aa78e71d642b07d1699400c18435bd4eda486477096df722fda438efc6d09023bb20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39ca8451dc97b43bd3abdf7d91de80441e27f3a71d2a317eded0d9de2dcc36f822a6c9c23722af0b9344c1dfbe3686705bc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcac31703b81759647d37192200ad7be918f3d40add1fa3a08932656b1e6f352abd9277ab46597981a4967d4fcd20c51326aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cb5dc4a7ebe1590bf80f73edb9773b1b453e9b4f44c2a88232a907ec03907ffa513009292d4ee3afe0c7b0910fa99422bd7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb09d6b1a23a836aa5587ce91f97bcae5170fbf3a671a9c4c15d9dfa25934a1b1599215436af557a1528d9df88e5498e042d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e53f759c5b5fb50ae250fbd346bdf95fc69df3edb281a94a34dc93b2aa827460fe39bcbbb73b686426e55da65f1ee690802;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ca2b60560255a32e521be8e9cab460ec2d53c31b7d2f8a987130ed81194959a728e1878fefe281f9db2de3315fce61953cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he44c561a8a2657b8120a0499e4005d57d713f9dcdf9e63c9ad7b6d2dde9e25cf8fae1bcd8a68b82c37cde18ad02439b15271;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc992ca06a85164b2121cda5db4edc552e430a58eef4843790b21e11bfa7cf95af498081a3047cbe1256c68017f784d5f2f40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51476a0cdf968446cff7fddfeb76c80a7f492b37ccb24cddfc9f89197fc20e5a407a359362d9da0d0fe26fee6cde506a28a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a7a0c7c720b42b7cb4b2d181a02059d70d10c79d911dfd3efdf7ce7bb804b658cbfaaf5beec4709da3cf0b64e5ff2355f22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfe3428f5123f349db3525402f06c948da485867776771c7a7cbb557a323177157ac35e62338cf9dd0de3fd4f75fde3de529;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9194809ef03120aee5dd60dbd375ad23f4afabb48eff113ad9c8bfaa4689e2d3f2e7bf8a45e34296f55aea2b212a3f182cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha03d3fac4b654f65283cd7cd12237d044006c30b332b44ac59c1c3e2eaf81924b21632c56212c99641c80250cd47c9ea869c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f62857fe143bea24289133f16960ecda882c0673df07b40dc20989fcd9a057096c8a51038a481edadc3b4695f3744e1e660;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5065d4230c741f77d75c3e4e04c376228551f28376bd86fc7d2cbcb08407a65e37b618c06e7dca0b4ba1a3b72a8f7b10649;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d5e7815afbba704527feca52968fe0fa6e924ddcc513da55763def827cb94d5dc71c74f70346c848ff962bef47b1e1da7f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bd92c2658804f4f36d860d6992a7530f5eb5723b33fbd392053491cde653d5b2cff1c0a96c258f11aa2a9a2f5ed9a715be7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9883a988b786dd2ecb48fb9fa09187f76bb816bb79099f3188f73f2c5884f6f579cd9df4f894f877df046ff042fb80b4bec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfa19f2a65aaeb9506a79f515e4e61e38b2f071d58f0711b0c97171449400323120f5ebb2ae4ba2ab5907f004e3d816b33cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he225a145ed3f532824a083b28e4faf9920235f82f544d2bcb80902bcc0d27facb3a3281a1cdb0df1985c8f404b3fb7a8738a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c2638505e4984d5a24c60422263ce0b581e5a855f907a42fc984b611b02217e055a9b7754c5556683d116921a52f3c824e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11b0085f54b0d76e00045c2d23f93b0673d704f6ae84aa2dbd51e22b5ff853b509918d50cc470363f553a07833ef5287a40c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bbc6bbfc35acd8748503f8c0efb33e0dd705ccadb4972bc861772186123683ee264bdb2ea6fc749e7c76f785dc38d31ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38ed365b24adfd348e0645034edf4fd5bf604ff8fc2cf7cd13fc7f7343dd4794933b221523ea1ffe3071b03a4d9ded2342fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45ab249a24adb2034d7478cf5d4919017ba5d03bfba1b654d5917fbf4ac230c30f91102912748193e373cb5189c03ef4508;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h709a081b01e175eef7bde3348dd424f5567c0f525a30eb1afe916251aa587a7f117cc5c43e827e2dfe81234e0ef223d163d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57cb943b0f648b57583519b79e8d00d4ccd5540c2c031ffd7a6724f5e4c37ba51298575132bbcb6072f989b31f19331befa7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78df4ca7bc88a3562dcfc695b7089e505f7329405dc1545492ce236767206459ebf9af470b5b222b7850e15c78aaac5e01e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3af6abfd382bd02ec74e0428fabdc80b6bd3b95b913db65e819357de674620bf7101e4b7b02ce56b97ee453e57b9becbbea0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57882f0037eac3f27c59d15a652b6c129a2c51e4e6c0b7c96f2d6cd78d3dfab055a81a4c48762f0de674f3e0aca772285eb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb796601aa409e38522a0b9ce616ef0d56c976b3a778b4bd32410eb3b98a8c3320ecf1dab7de73075342dd4713c05f141b4c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haec83ceabc4581fee1398167d1d7639ae17d58f57699f7ee99b383e09a0289271962a7d8f139abeb404d11b784ddd1807050;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h868505d1fd29c8262cee452acdf8480c5017a505ce876681ff97e981b052107a0e3a8be5fc7ad2a77b60ea51f11fdbbcc0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcca5ca48b618d1377476d59f5c326d184cb211c662eb25eeba9b3f871b1eff88c15050ade876fc1636dce15e722d7b91aadc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25096abbfb591922060ec9f727adecbe9d6f35b1ad61467b1e10d966fb0c7f23ef885611fec4782be075b9aca80cefd129d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c214ac5d100df036229c281f901d00ad2a868286a7ff8157ad738886e378a5aff802aa2a11b08c1d6500317bde4a125c5f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d56f48016e0d1bb4d4bb19cf4e1f0ddcbdb5dfdb883a97babcc9238a0ad474692e2e0265a65651563d19304bec2797793e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab6e90d742b77be651b5152fdc793b2a110cff4c673a2b397ca2a8510baf9b161a5f7d38dad070f97a8ae07f765ccfd26c05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a109aa5350bee245c4a915928465efc40dd92bc3b0836cd175fe960d62516e4f007331dbd5e3036f2ef762f582319c64a2d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62d8d29bc19f52b6c50eb3decb57432d4830df0e238cff094136960893e45cf376b6d5752723c62c18801ba73508d3219f39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87c7c6427666dd72dc4d4cfb628d4757ff760491520a37b635b33725f448be879a39df23650b3050a2f7a86dc65b1a451c0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97053d2f5f5b31b20700070387df1677070f5270f8bd9a19bc0262c1f384f45ff384643b74fc22481a0d14ac0ad0a411a50e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8601cb62c1d3c348ae762848a6103fc36a004b2419cffa19e4c4b7235970273c377034d3e578c09b8997d4417a144b8013f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1051b0cbed8f88ba268f663adc7ab5c59db6f00301d08de8b4a69427d6820d72da93bb6b6a4f9e5ff822064373eae4783e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdd62173cef68dbab50ade25738e60d7878b85a192ef7e5921c29fb9d139e58e7ac5675de410ee9f8ad0530960408bf2086e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8310465286d03bad8c8f80d80bc975cb9020a9ecc191723b4b4e603ebd2171a4d60dced18f14f2f418493a173a14d348701c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h781ce172341b60955d3a3c0daa17c79379e86fd8143e71965e1ad5f8f1e6b3b37cd05803b396ef9b661d165d2b37fd7f30f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebf1c9bb26db7dff9daad3fa0119d54f69b0a5654bbc9f4054fa80084dd52a8a069acec7380f773e3a6326e7ca0595cf74b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4483ff35a8a7ac3f0388461314b7f461169212c5c8fe8520d830c1e829ece6f55538ff773a4cfef39e73d18c2a2f374c4494;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2202b088752d51d408a58dc9b61755738fe4c0e49d86c7d6237cbc5b2bb98b0e99f9298634765c718c4bf2866ed6d6eb3c7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8486c5dbe76b48f8a952377d5b497942f804c9968cf20939b30d303f8813eca7825bb1b1b2a4d038f829f89554d55530b89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd1b71d776ce9ab6d48b3631efd4f6a9ba9980c7124bb0e489a71c9d3ad24c30c28b6e088579ffd6a1949d9ffd2f70044d9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96611f6536a46023a0e10ae4e80f6e3b4e3773f2dd09ddf0d2ab82a6a4f375bce421cbb8688cfd67c5fc6a9a92bcd9556afc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1b82a7e2910e04ae7c14b7df24cc8e3b8e8a721b0359749c59c595697751006c0f58ede5969c4f4fd6685aff97f8d691917;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha45c49bafbbdad9de9fef4ae0854c560bf49cf733c227637fa21ada9612aeff93f065e17a57f0a909cfb0a1219863f5dbc01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cfd592e5708ddedfa19f789e2b5337c5877c618586c697d43fc43604dce1c80b0e7586e4b847bf0529d74f56b48e283a946;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f66157d3ab2aa1d7bc849d0121f1a9d5b45f5f6caf7096592a80654bacd397dd0a40adfb5a4f8da66a21d9f97edb0481f1e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41796884fd3afef2b2a1e316b53046327da73fe0e336840c000204b4793a1ad8e652b6dce83f81c5fc71b9281b852be6297f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h370281ef9ad142025eadef486fc5506acac07ee028b9e64e03a10921dd11a2d1a636bed4d0a2b456c3fc92e633eef97fbcc0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31fc7aba52f6f49ff84eb73799649fdfbedbbef2237f5c71798d384aa9173534c8fc1a91677288f4d40372a0928448efe34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3deb301c86354c068e600a2489a6b2b8b8087372b138c2611e59e5bdbdc789d5c9192e31f4c1f19521946daecce61f3c389;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d919f551e76044f618ae312225034e27e96526978610ee5bf3702ea3e417f9c42337f22fc7b2db88401a4ce6b07280c928;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b7467f250fc6a78bdabb038b2edd971eda9d3e343736e4ca72d992551d25bd48c15f4b6748000e7ebe3f0d6c95229a966f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h934b880fa22740308119314a37fea95cdab20ff20dc074bfdeeb14056b11bb017968e40f6f97385df27e490dc1d592f3205b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddf00f1e83b2769a315c0f29e6ecad212ad6fe8b36406e61fa853190f5bd9ab777af1ee0225fc0c3d1f03f2e9f3c650a03f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2eee48959eac9a47d2c6dcb40ae0587e5640021d4df67d0a0193589f8ca0378c0fb5ed8b31d6ed5b0127142014718d2bac22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb521196bd6e7c1201af68b4ee148d34d6bd1aef299563671dda42637429b92c3c4a39029c269d7606435ba04998bed08d531;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb7ec86f0ab047056d667f124647b48fae8151cee93a3f690ef3b0329ba73390d006df6ff2e3cd60786f743272e8460da434;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habc3ba4517b173c6b29cd128191ccf3ae309a5c2c57893bd8e5577a070fd0c4509da9611d5ad138145e0d4e31508ff015eae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82bfb5554fd2c092106870a52a46271944f01e23ec5cda2b1649e3505d59d83804c1b3182b6ed30aba23037148554bff6640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5fd6b2a7ff93a38955c30fcda63b835c0b0903205cf53c1af841adac3d5a4a2a68e4c6f848f22c8ee74a65d880d624944a61;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8557c25a181c175fee6250168259c002f6c1a7cdc4a78dbd87d6e99d14a5aabf79fa92da09aca8b2f736ccc1d2bf8b450a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h748a5fab97738321add478b762f3d1340fee38b868e60aacbfcba7a88dd0a7266b1114250b95e4742243e8e7dd2e2ed746ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4052fd4c063226facb7808599fb8786a1b1b3c3ec70452315d91854080f75451100ad2587a26a2f188c399fc2107f7dd41b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e4501b92b30b0865a3384628f32cbe63a7371eb4fecf8ecbb712a7c52dead402d8d5a2f97775fede2dfee1e9a64ae4f29ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd041f0bb74df7dd194bf88272516345620896723e6ba61fac54b91891f43076926272f5f2370d903667aab4cdec1e7fa2808;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ec0ce562b67290568182fa743536c6745f0e0bdf23c0afa12af631decdc079d2815bb5fff0d1583b91afe06d20e88770e75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb5b14ec1e32f6534881f67326a6af6f13c008ffd076db372da86f11078465e55039c0f69ec6422c41c86b2ac876a710ab5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45d298876f38afdeb923667119d2e97b746bb1c89f5c609e404f5442790f107517e78035c94839d619d9f06a087655815996;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda4b080680f19f7f299b484606ae7589fe7e3d1bc0569d405b7434adcaca84fbac27ade7c8b7417bbd8f276c8f77bf1c4220;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99891666c1548aeee54b96a1950564d79800a779cc9dadb92a60dafa837b2cbd3c0c00f74e9cc48892a7fb4d06de720ebddb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbaa927bfa55d5ee46b2c87facd2da40906c329212b6902d147a7406cebdbf2d53510b4f688f64a2171df942ee55f78f8fe6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d903fa3e639aef8d51cea07fd78d036861ad09e3c3e072bbdf1b7a0f5d92759297c7f9f945361378727fabad5af15cb865e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd2b5e408095d8578be655a0c56f3425ea4989dc3f2f6c93d170b8df7996f7b90636fe9d688edd529a0ed53ed28044c5973e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9b4bcdbe98053404bf0d8cc15aa4f0ef3bcdee2010aa439d4d9d5a53cb025899430a0ef38537a69e284c7a687806830b4cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd28337391798a427fe112a217226cae8b487984280afaeb51acc4ecaf48109a8e753fbdb4c106fabb6d346f7503f8af7608;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a01b3f29f25fac0b569df98fb043f87cb28c34637ae3fb69c2a942ad9d3ff1df44be57b3be02d8a7e0533d7bde760f38afe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c067ab7bfdaea478a2bb5090ee7fb9ceb5d14b43f793dc844d6463c594c55a007d534029268bc18a26a27dcb652dd0dc914;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf666d156056be2a7abd4419f4e9869161e1f7bd31af49b34848f156670f77738c1fca9b68b14922be381f6e7234c34e89737;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a22512b52921a109994ed445f0d3b6d164da437210634b150057530757b8e475c84a1f4ce385fc89d37e5605aa4ff49a579;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc390a3e9e04cb0fa43e94781b4578744b50b99b0e386c8875adc937854d2d075e91a9c65f442b3db34017d7bea5a38e24ace;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha418e5c14e59b9980d67d3152ee70ee02e59d8d9f1255428eb45d40d3b60ecc71c13aa8e07205b4de89e507de69f3be4b196;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51ea5b6e89d0e263bc6ca29f4321f97591f19e00537bbaf8376a5d240ff0418419bdf451bd0540ecbbbbaf6b181e7502cae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a2bf518716b3cb551a45ee67d3a9cb6af14cf73e9fcf5f7eeba15033985b7ccd8b6d70aa9c7fc1bc2d958fa0e44687eebc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd75c002bf2599a647f8989891ba6c6681f8dee3b2142f3d199105919a82c083c43dca3253d2be4ad2ec00cda9cb46171fc72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b4c6f066bee8de517048b0ae2252528cbdf1f8bad58549561b91fd0bad9460c6ebfc020b85529fa65e52408d18831d3f90d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbf4991de627011734ec799d83ce9d6d3bbb627193a3186af615bf401cc1eb65fbe4a306178a1986fe9a611dbc9bc5c16ec7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9bdc07c921c6060e071b0bf5650ce71c14a496fef99888f65ddd3e8f2e0660fe66949ef62e4ac2caae030e181adcf229fd7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h859a37d67628eb258222f5f8379bf2420c02d28a745589e67bc7a5a631169d46d1510acb67eed1775ec02a170ed54b1569c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc007ed549c27c51b5ccd2402f89a4acba7a7b8425225bd1df18fe3523e6794138589b221e4267e12d053b1527798c1273aab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54906b023bbf06edfb830cae5438c8ae3c031d6ff82f40664a44a700e42fd5034146d152c306fe1c1b938dc674e475807ed2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3f3d8a26897007eefbdffe5a8238148c3eb73c8c27b43349a6da5e9c536f213573927f4da67ae65f04590832dd5b1892053;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h825c6fb8366d667dcaa3579ccfa3e773698a3c5454d8596a5460b74874bcad9613e416f07803db6db7ffbe324e6a8189c6da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5cc2ccd2e685213a54f533882c939fda7a6a31b6c7d326a6c68584c35f21d233bf1b0c9ff798b11e5dc2d543aaf5de370221;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h370ed6e0af40975a80fb275c75f3463b47eb91770c55c768e569fe2603316bd1dc6f86e43b870c02aff22d10014b8aa61292;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53de703b5a9269872061cfbdd1257608b83ca8dc525bd5cf7a3d1db1ce5dc0ff182d78a4212cf342919662a6b890f843130a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3ef7839ea2ef9c981825852e223bd14043029a58df02cc13b173eecc28f5e522341b82282657db0a34a3a3a424fff10f377;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb93905b60f28c654a15f63a94e745d73b58a2e438eb10652d6f1a154f59dc48fc8d05b14294a9386ace241b493bc82cf2e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h192e7936b8a34ca91a8f2a1bd3377ccbab8986224ba62d0dae81ab4b84c3626d6b0f74987f823487d7707dbfc7e3776fa95b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h718d8c1f39d28559de73fccffe4943200e9963337a8c5b6314fe697da0558e9182df45a82a8ddaaba59b501851199f3e136b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4eb0dc7aff82c7ed4fcdd65a4ddc85385ff1eae7bd1354af310b962e091b129381ba5e61ae38f5992e9c9c683f104a15d28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeac6c93db7be3ce8f526267db9f1d84daa1b87ed4db22637490b92148aefe4a28348b073115fb777f5394e9293fd529e819;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39f2633127902eac98507d3e2aa3202f9a9111b6b53c77c1fb7038c2743ee523bad9f96d80226d7cdb08a30d24a6844ac332;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdb2c3d844536136ee171a421cbf65b8188fb1cfd5236004c960a62dccdf73c947a84343b012cb8de044760305b66e3c733b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14ca2ece27fc1fa08d7cb53740614944c54c04796197d7633a704a7d9314d6a224d20ef05baeed368441a162f426073eaa42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73924c3bad78468ac7b5a7aea2a44050b253d8426e8e2673ebf22d3073ffd18011f0753ed297659ae47bbd5c429dfc35112a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha97bc0a9b5c029a7700b676f10de2528e3b67b0a87a0935b27bc78b7e3db63c8bf86d07a0a00078921d5feb850ef55397bb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f13627c0f3b78aee1f174d55eab59b869a9c7d23472badc206753644944fc2a986d29978e71e4f72b41c5231cfc7311c756;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb02328e359f2a917bd3b92da88e6019d906b7b65a5c1ad4c822b2fa1ae83855aa06073660b23909fbfcb7175c6f7c7159fd0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcc4450eb8a4b5d871d8d037f87de57cf981e07e48ff2f9a4c13ef9b0991738441de195660daa3e1c3f365386741257955f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h762620c7f455da495994991226cbef027e8a7649bbf32a6071245f050143a014b16f3bfc0d70954ad7586a77dbdb1fac496f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf7bcd265784bfc54d6ed822e493d927751969f2cd9ea01843cb4781e6cae111594b1ed939ebfff1d753546b49315981115;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc565d71f9c60f1f0442ec6ab0a39c2c8b0eccac3937f237a1677912fd299f8d8ba3215695b7cdc96f1fa420c63e9313d856e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h455199ca115be6a505412d6433430e7a4a68e9368c0071f19bea3029f40f6552de70828a0a2947fbd3f3f2a96c3c1cb20c53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7ded47827395e685b960ee26281c7a503ec16f38d6c94b7ae48fb410bc652c825ba2d8ca600e86c1b92f24d2a00cd2a349f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6bdd2cdac47d7b0039f95a594d052d5ef71c3530e6c7fa4189b280d7a9f6fad9f18f3b6743f88eb6ee056857eb7aa7e0c39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2d944809437e1e3ebed633e6a9772065c2617fa44fd84bb7b7ab5d8087f4d7b657aa167a92f9f0125ae2f09a2b9b0ca5c06;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba7cdf75690abdee124bdc129054d46d25e4b9a0a420179397a52dfba58ef014f2a6c76b49f68ada7680f91e20fb0b5bc2c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae4ad6840f696b06f35969211c4e27408e0e04a0e74b64ad8a85d20a28bb7f783985c72a6059eab24bd52abcc5665d5584fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7abef6ac40bf1a99d4335ddfb96f42dfdf2f19349ad19141791ac30b0d723831efa2e19df036fd0e11b1d0955023b801342;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heba6446704f8fcb4a0344f813ef31e1f2fa8edd7a774d445e35b634c23f6e926e9510a7f130856f412c5ddf584b131f37261;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h244a50b462e4ace958e8d70ba1fccf384a7c872bba7518cbe017b1f3e4b3a815876f64d572cb4e3c0bebad301ede59e613f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb15962e0e25ea605f20830119148dbe84dae3e9f6dbdda6e3186794b12f72da07fd6c69c6053c9b63662a6de22b58f0ba90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h501721361387d82457c49be10ee8f51c08da5576c5d78736098aa590a71d250855643a2117c6c078a6b8f6937623d9d13836;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h789df873c5f66882cdd4f3683c41d7e26d8e28438b10390b0dd24b56b3509254d9accab030ce95cad6951f40c841715e3e89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h120a1974fa51a9479514f2eef5feecf5b00abe206fea17ed35a9a42051e06e862931fff71ca65febacaf775a66a56b10498e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18e8ed96578ae753972d0169072beb45972b96c69c016cd288e3d30fe182623c6dc228f5ed6e42b0d88a5d418575d5905c45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfb81604b0b09ab3971983df652b4a373d3db2e6be0727ac67adb485573b2b83a31cc6af616abcb2863e75c3aecff7e2fa78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52c47406bf828f19ca1bf976c26d761b0fcc29c39fd862212f1082a4e36397be93cffc1b791466d558bf8cc39b16b887ba2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3f5e3856c0ac31d824a8fc75d32788db0f8956c284d4a1eeeab563bd22a12dd2dd138a914bb589e0d01a1c455b5744a3e61;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf5ea1673c547c5df4cf7a0237186bb7d88f6eb899255eaa64fa4654fba5c24fce89f047fe5dc8f809c27976300e0625422f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habf1e8409007d1683c058ce3c4e12c81e7d310602adbcba19c78ec7af47b17e17fa6301b61ad661189dbaefe3ef58507371a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h303327b2857089a58e41d29b45ca9e7bad90ddae6c481504f5ecf25219b9ceb30de6546f788aa748dcb65adf9e3878016c6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bce2c69199df9e585474f00efaff288e517e1db01b8a216efecfe5cc0fad461fea1194c769a46dfc12573f59f81d0bbc2fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb50b12cb853e8144a25799ed6b3dcb13c453898d8b1fa298b0de3fa512f474e4ff4e6197925d5372978df48a8c1481b49543;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11ea48d44f22d0f732a9cc6c892c691a8be4ab4ac257926c26208f02d67ee31b63340d0849bb1a0e4f2f5a987e8b20e32352;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e7754498746c4fe82ecbf17748f9408fe0f85e0f0807b3c11ce4ccda1ac3dfaa05b3902ed21ea08827b4ab80e47c1e5f145;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha208cfc865b85eda645840f5f2dc9deec03248c8eb30789433fba9b6c342c4b08efc8f30c7bed05cfa48b2c5d20781b6811a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7d904455b4d08cd49ab2f7b6904a9ea4a81ee5246a187044ece501376fdb387bf579a4aa82ce36fcdfc23c5d6d9db1878c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cf7e4974c7d6acca73402747238d9d0fae528697b8bd451bc818bb45a76d1cfe8d5a0a49bf419acb766d372dc800f8b3ec0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe71cc20ae79f42636cd3dc30ddc6906a393577cc357bec49166440a44c4d4ea50804c8b1c99eea8a60bb9c210c60a758dfd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d4f6bfe7485343d0264d6c96a73b583bffece53bbec03ef436770b19d7bfc6509a3a6c8d0de1340ca8072c667bc928ac8ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70b36e53e4bb0e5e757f4b50f4b9d14e76887bc5908513c4c1d7c60e706bf14c2a63dba74c51b58ddb3036adf07f52609a5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h690f9bc507c72fa098ef7bdbac09def9aa821c7f33a3b3508d1fde41768a56e96191c8bbeb54e07f686f189130c89df62501;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3373e01d25352b5dca9d4e05008e84f70512bba8e790eceb7fdf4e4e2c5ecc3b4966e70b07882a085d2332c2e7671e47f374;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecce6240eb0f6cce4a736d04063a4b23f84db13471699b2316e64af2e0597144f89a48a8c6abe9a481ca0e1b691df95e31d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h331fb88eb530b406c1b1c6cdc4a68a2417055b57b5ef5e50612633217c9addfa6540cabaa9414dd214f8ff33a526ac34463f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1497989c5fde76cee0e3907fb2cfce17784cbc36470b96982fd04d5442c3b1004a590e0ad99c21201ff548e996b4db23b83f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe416ed067baf276a42f09dbce59adad82b813e1437164cb33f71bff349f4bb5809c94251b6982f3fcd06907030475d857b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9393f6707831c832ffbb41b8cc397efda6c6d841c852740324c0fbd0b491ee5de10493063c764ff87a5bd8cf628f2d84242;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1847e42249a1b22144f9fca16d343d6db3030914708ca4dcf8eaee2af3f285b41d31b8ff829b4ff5ee02145a0ab3a7748b38;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ba56b33c0b698341601e0f3bc49866e2a2c418f2d376e66c120ef0b2f180f4d032e4ee52a92f5c190692a5315e09fe40bea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b3a3d6fa6516e42bfec7891ed8a6b2e69d0ca0e20e29f9b3a33b54834e587bfdc52d798e3d9eab150ec0ea264728812b268;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce80e233b1b5b8c2602edee40594ebd74f24f29cd97ca30f69f27cafc5286f7317fc5279c0704d37bf738f0d9386d0604a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdae4c8b98593513ed5455135e5a0bd2d383d8ec244a87f818a9dde942f946345db59e2abe5b00b2e0cfbb224409acec1f2b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68171948189095308eea95eba94805bc75b39e7d78797fdb45c572a1ba3d116235103a61eac7935fc78f67a9e07e4011511f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5044f8dd8650b9c2bc29d46df35e72b6339d76cd9c0179c83cbc74066b90c80cb561530bf2ebee323ad12625fd1a8a1fedc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb315a43613496287e388e15c81d51c4f47b1c4179bb6188e0c2ddb902b08534ad053883fe721f4417fc55476857baf2dd5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45980e89f3c929c694e8bc3470307f4e33b08d473fb5e6a9e99c552aa1e678a674728231a5e582e4a56afb701a8aefc1ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbda6c445b67649caba9e4ef0aa77068afe8c056e2fab8f3fbabc39ee0fb7c33114392be478f381090c2ccab6ddb5d5e11f34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc539d3dcdef38138ad61b13ee7f1a0e85220782cab26dbfcb936c02ac3906449ca3908ff2962022d73d9345d39700c3b7646;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35b9c85a6c2d4b376bb30389c02210bd8a79a58f06b473e58001a5a2a9d2e753ecd7de2a3bf8b9fb5d106fdeac82867f27f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7426f4b07f1a74b332789253963c5012db89622e59a7b9e87c019f62bce3ea3fd9b0408b3880a32f679fd62ba7bbd40e6d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h157b06b3798414acf83a17f0db3ec1b5c8e0d243e71e472c82ab640f44d8ac70b86386055876f39e2189328162dc232cdcc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7afc0c38ffa5dd95c5af8620f487b9197c0ddd4f6fb837adac58ef6c095c09f483037fba3975eea619ed6b98e434c0a856fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h489d90fda3ca1cd951708a900628d662f66e7013944882d41d63389e6d74796e0d59d68d0ba711e2e2768f56f636a0471172;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h563ed666712d023c8fbfd83d2d2ca8853a8abd7e58524c956b38b0312a79f208a8c2f6bba4ebb922828dd981587a16942bc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f333187bdaa29a1786cdf9ed949efdea5ec7bff993de74bfa0225c3afcc58c72f33dc301cc3c3cd818722f08b26f6ff633f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43eacba0837cfda28ebf8acbc00e817e762d9c29ac5c558307033e839e837d4bcc3391d2ddb690e1bab2f25ef0ccd00e5d2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74c7980eab18f3ae5a35952e24be41869c5bc07b2494b46cb899743b6bb2ade85a33ccbc4a7ab3b36228048ee1ae812824b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d4811bd0f08da8593d3f6fd69a88cdfa5e71d028eb1527352f81352767f3334b2b0d541984e85b9b8a9ed22b66462345042;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bbd65c9d63a0b57d8d9fdafa0e2b4a15f5c46e5301ab00bda22cfeb81a17b990ef14f2666ba16f2ae6e269008ff526ee4e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4ccfddf819870ae7caac3014f110ba831f323ad6879d966279b5c516851958ff03eede6180f7d8bebbb51104ff679c5836d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d5a647146769c0c8289f9a901f7026adda4ce48855bfc77472e8b8afcd31a7b3380369f6c00675d5845e929ae368b9e064d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7a96c68bfe62d81ba9d2d36b3e6fb9ea95f7a0785a7d972107749bdd7f65c325b8532747751bddbb6507e924dffa838304;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60888f015d73996868c5b9e530bf5e411bf2f79f13fdaeea1f9afa7a1485d8e29523212ac2afa271945c3a453d2bff2947c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21968283d01b5e1cea8ef82d8097ea6d177e76251981152d75c0d505b78b8e131393049d7cbfaf42366a9a74f435ef18e355;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12574199ce68a891635957fcf7a212208ed73eba50aadadd0cb9961a16f76a9b83e746a00880dd86608b6ef7ab41e61c542c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b7ff5424212fc4b765a49461c6f016dd6fe1510be0ca5a0789ba6ad00526a0b7d506ac46f1ecb4c0a690b9440afb5b5b9c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97aeb2c79d7bf9e33c6a570282c5a92b39194caef8c582b481a545da46cfdeb3f4a7f714ef427207f95121b6e8bfa33537e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5fadefd842a088fa336f764064f90d7057a75ac478b7fdaa06189d288e8f335ae848e19809b6eeec6c5cec329665c4ba58c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26c9c4824ffb4bf3f530dce517c7cb59e288332c3d7b1dcc944c69a0107d5ee993730581e28c0fbc9097101b1649e3d5a764;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0473d88ddcc47109d0c20de4c5121d26b1c0221b2380711202c61b33a36fe12859b46b106c5ca3cb833fa41022df96ee691;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h507beff573cf945ad248ff4bc045215330f7cf4e9c05b4ea33eaec96e2d8b84daeed5ecfef3f1fb3dde39ae8cb8b110ce66d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d41cb26e96dc3514b0b627739e4f24ecd61f98ece4b1ca5952f1a47a2d573df6e2185335578e5b3558555bc5aa783491304;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22a3562674c45ec892e92cdac7df0b512f50cc9f97c1775a797756372aa3f3c5044e0b587e8a735a97ed1827c6c53b52a92f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb055bd07d6fa8850b6e6ef06e9d9473eaaa5f946668b387800aa0283573514fc1742ff21b99d9d8750fd720f16a863ef90ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae525e700d8c2235a6b1534f8c4a2cad758f289cead22a9300047e6d20aefad1c3c39abd4671ba8d63b3de6fcba9284750f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2ebda68fca8c347197dd0e5a00db3bfa4427a53f5b62961cadb61efbf8214b9c961a13848e4ff609ae77439cc2e2486215d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9088ec8818022ed1d20e32bbc0590c0838731d3f01e2d67e876e1455c9b5a5db089c8e0bbdd84ad8cef892bc903248421e86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h110d1abb2a5f9c650a2d87d2d7e141775f6d55cc26c475802c29838f7ac5faaf7c2a8e4cde473ade183d003eb1abca6ebe86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70908f56bbcf06463ec10f11d4d1689264a21be1f39f01b61b9155e46f8b909521bce2f69df7af52ac56a2163d4578caae54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffb9ec323700eb42ef8fa48389a62980d2ba4fdf93f03147520addb0e7d435a9e7ef810ac30ed966d3dd890478486ba8e9b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha867a904a1923effbe44b35a30dd83d2779b4387fe45b35bf72eee3d33c0f841ec2e5fd28e663b0359c80bc0d94a63388e34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ba2b3a2e989777b8dadbfb319e7ae62a184b5a37a91a40175f65a9f48d6890e36150d56ef2581ce615b910e6b09fbc5c70f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4948f335b8f9335ede6da85de2c3c3e4e7312caa18c3bd5117c0bf75aa5d2ee9b82c509e3ac13ca649c6ef40f3103a6957b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3028b7078a2d6c570e3bfbbb2509081d6c5b64c68f79404fb5469e36f4da29dcdbee8db240676d4c1615caee543a31b5a616;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf00940421201ba70d789887f8cf5cb3b2af95a3e3e27ea77519e9ec620e274d1e073f4310605ff6444088728b1d6bf8acdb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ab8ca7c1a91d4605e103d9a901c00969c5ddf7dd5cf9c868015ccd205a1b5fe0f7ae01d9a900712dca4d1276038e6dac4c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ffc35f92cc33e537dcea29626006b4db432598257d4b49fbd46cc4c89437b89afaf772fc977d67114a08d11423413618b8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h867b2de41007da00c784f4d286ba8c535ed8330bd6b007d03396aa7edc7d2948a457bcd99123cab2f4c7e30629d2f8ba4832;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7dcbf9e4c7a822eb105c2b691c4af111b730c09dff4329cdfd31f35d9adc6f472cd07f52ea79d1807787f6995639c54d63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2770b6db48e58f0d21ce1f241b54edf2d4afa5ffc5f23e95f462ecefe1fcb476539ddff8472a7cc14c5133c499e3ee297780;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdff28a265619f383a085fdfb6e18d1a4dbf51499ffa0676bf551641e5e6e7c0a24606200159bca9fbf713b6edf88f2613742;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcae5ba57a8719f72d04e2412ce9b474273dc0b04520a636d4118c57f3dd6fe2a7c6efff3b789bca3f0696d1c4e643bda926b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd316ffa2711adeb37be47fd9cb9997295155dd10eb54959272af9ecc28e0dd6e75a388008536c93a5873abeeaea32d4ed4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha37afc6b3dd008c94b03eb7159d32f60066d7ef8a1d3048ba3102565af17805b2cf536518eeb9856d407b17b2102aac49a4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2346e416340e52ef0352ac61e320b7545e571acc7fafe078801425c6ab9e2b4c24991a7bc01ca982fe5b9aaea1dabdf527ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2686c31c30ef502026c09bf72e5ff2a09e47dc713af258e71055722398bbb357ab690d8682bb7ca8977db9325e25e93181fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cb04d64d880086775b56b9db7d952b2db424a8707e068fa85179fa10606f124dc725c5163f8a7dc8f372c977c24808d6d9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0c1b3209abfa485ad76beead9edfa144310c3edcd6f3d7e4b83fe4fc466730cbef59f5731b3b9fdfc1d5907db5447e24f69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5c1f79d9f17b8cc403073dd1a7d45e09a850d36f8749026021fcea40b5ad8c9d48eb138edb8bc714a858b9c5411bad56bae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a55f955ac60e85890c1e9066c7b8f150952abe53f931ac500b96b4998b4d71964cc954ce69bee9183df5e4af1d889a71d64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fde61dc966a8c53d4e6be745a7ed5885379665e1af828d30c609c96e354166b88b909b6c64b1352d40f2a329977f24b2c77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1f36d82de1c8105c78668b2ce33b11407a8366e57f8ba742d9dbb328b495cd8498b38f9905f9cbd8f9e53cc71b0b2ea61ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d3069a97bc0e6c37b399f1bbc0a6808e07676de17d65c343a55e3681848d8d27d6b71bb2e790b7c600c31b0a888bad86c8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4def73760da02010b291d4c538d1483e395c7eae0da3e3a596d2cad2f5cbfbc37482066e2d6a28df61c0994b7b2a661c5e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddbb9abb83e6d403baa4ac206f7567567f6e8d5cde06bea4c10784b01a818d166dad814a1edea4bcfdbcde48cd6d5e94496;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf72e1054964e6149f2e92cfa56f0f4cfb4d2a6a5fa7faa73f77e713445938f6f3cb2f2098da214997f74e5cbd5dd1eabbd42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79b6f3576ddeb720a8b064bcd31aea249aeef90175315163b2cf9295b6646b3e78cfd596e989def4862b26649e946dd5cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6256cc769f990c9225f870148c878b99bcf3e7b41d6c959dbe2e248bee01e7cc5bf86e8996b1a8cdd66b93ad192d7a20a33f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f2f3095cb52ffe630f211353fef34c56c0537b1eb74a2a10d39540c9d9141d8db759fddd2e14e197540a69ede6ac1e0637c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8383b79e1985d8d2fe3c4e0a10635f8e02a9f2bd7dc84a1af5b476602f5e2aa69032df8900bb8b74e897654f2f1727b758ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6f88a485fcf0f8d41792eff3b603dccb124ebace91ec72ed692b44ed1311489626d70f61842179169f1411693f544e4f63b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4a1a8625d90211687da110a23e811952a23d9c969be5c5c7c782e26bc32f9d1c903b274b02207582e3a117bb33cc3e8c3b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d2e603905db6a67748ebb3bd05af006646e91fa21418e755df01ddd213cc1b1dc8c00e224d1efea42e3ad0ebc947abe809e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91c9964b4a8081c92d52664486da2e311347fce60d9bbe74e3a0613d08d7cff9c0d98f01e880b09105169b11e08d255750b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1358593fac086d355b28862ec155aa8db6a1b6791ae29260f5d450f3a77873735f2a4635e1ed8c170f9fc21d16af57e00c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6a5d4caa57922d247e2e530b1eefabcadf3efdecdf7a44fb70bd5d6ea5e72556079f93f65224781248493f00b1349c1aeb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54cd385b8afd4b7eee6657fcb5b1f0476c3050c83e2aa0b68763865307e351885511d6cdb70309e415e8153efb9b08e873ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3adb193d5d8b5bb08bc0be5872e456e148d1da4e29332675846a3665719ab86a86fd27bae69d576eae09dbc2dabc404db9a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7f6ebc125f1a544fffbad0332ae4f68af88f381f4ca573c41f289602a594fda307ad51d63fe6857a58b64cea4b9168f976a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd54313f06ee1b0555225cc29e04b5a5f8ebd73cfec9e0cc79a7f0cd52ae044e9e43a9bfdb22ac9b818ec5f4c0bcbb0a9f9fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9915a5e8c3ff792b1711d6b0def54d00c02ff8e7e428c87655215ed3d80c932be8bd521f296bc779a7a1f221bf827f00d2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafa30ec7e36dae00bab28f3cb98d1156c3a5f1b9d24da591a3a089ed9aeead0317353d45a1f42f4246ef2f9adc8b58316b4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb65cf42ed0cf89d5a80ee69032b7b81e2ce9ad186bdec4810979533030775d999eb2727ac051b9bcde45564597a02074ff4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1077fb1b72ced25df61c33931572d4a7524d9883fe1e1513730d0a1f9dc21a1a976effefeb7eb6a3e3c7a5d2c11d4eae8b99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb5a1aefb13da2458f1c07cb5456c5593974978365419418561d8efef11b1df3c8d4b32a7d71cab9ea1f83281cf966caa8da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7eb8070462465e3b264e3aef53290bd16f1e8bfd926157789ee72f09172e55f30c1572725abf17e6102f6bae7cfe151affeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h591de9f4deba92738f720f5f15a1675c056727e9316e7b478ab015e1a7ab5fcdaac720c8e547104b452913eafb2f3b769e67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6df502b6fe3d9caaec4485409d321de1a8e7082760ddaec8d0553787a817fba6c169dd9d3732b9eaea3b7d280653f034696;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec9b5e0c0daee728acf45f272614f7977852db1ed93d1e1947198c3fdf017499b52f1835d97746a382272605827af85f35c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9898c339d1ee301505e393419c549135636a273a216deb901725205680a6c9e3ea5aa6ef831a5c4f927912d9987b49e11b1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha33f2cf951e46e199a5d4967a1ca4b691b5b408eb960fe9ad34c19222962aa38745a0c64f80f44b6abee300a64c883996eb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9eb142d1a5daac4bd7c265f049bbafbb28be8c4a299b28c5e016d252cab98e4d13fc9d6fc011645c79067ad31b88bce3539;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h907055d6deefe257cfab34f0bb443b815c30ad4e0224a7eba16073794f1352151c83e69192b35e6029286eb70e8ddcd0c579;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb3bc6c92046e01a706e47b918c0eb5294331f61163bf6ddf3b729b6752b320e2caef663d3cb4e30cafa5eca8a86d7809369;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb299a27d32f2f133c423208de417820304d3e85792645994bd84efa7e62a6d0ef38b239ce5b7c4ecef37ab045c0b91689244;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19b95b0558adeedcd0915594f11ace499c47dfc1fbf0dfc588ebe5b47cd8de0c0a32dc4caa370544174bcd1123bd5330d375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd760862c00915b3ca68e802f59a3018c6d50c0cc9a7fe6044e89f4f9180bfbc2cedf1e27be7c249b1e4522b5a2fe90df667d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he62ac9b4aae4ffa0cc14fa30dba818edcd0d11921d9118486db18a8f012d73e1850a79509e068d5e5eedc89b0e43658526b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb72a12d34709e00a00c8a9676c505b7647c8fa32bbce95486e0147f27744d3a4b0e76f6a603c5153686078a65533143f173d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc68571142d49d31a0b13404ca80752330ddba46fdd14cbb92b8a83c730cbab8dba2aa3db76ac7567b8dcdac696df46c53cbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c6383c02d8eb3593fcedf6ec62757eb47f25e7c77f06d18445639bef16d2eeefd866e98943b4934e956cc3dcf97e3f04627;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98eaef4b7a7af4e6c6365377715ae8a7eeb51d5a5b9a6b53d948087f35eacc185555e7593e48267a647b316a9d3f06f39f39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47f9ead6ae1a5544b1ae414490c8343547741c948cf1e5c62983bf2e6d86a749ef9b198e83cb728f8591704628acfab32d23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7671f64f1302e45da4a458b550876bf2e044802080a9525b143f7afe40e5f777014ed0c35dbb388b63ddc7d2ed7f69cbcd0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccadc92e37cc1c5d225da654166822b5db31a42b1a03b965b25ac22c54f8c18f9df3f46487a878db1d51f748f631989654c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcbca02f170204f79e081bfa2ab8f66f0cf0676539e772a720aa50baba820527ec0f481da3fd411dbb160037cbd97222d3a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12f479fd5773f3b3809a9129db9b85bb40de4955cebcb19cfa6ed83767479efb5d3a8ae450dfa47f9a72a1c5cd06cd3da066;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0240c7993a9213782b7e5e6bc2be980550ebbe895a6d4d4f497f233926feb71f0645761dab4712d7abd7778dc827a29d54a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf9ae0fd5d2cf3d91727bdc10a5185d328294b3f0e5fc6b3bf0154a8d5630d84afea5005429e29e316a6b4aaa619f8145b8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2139bc616294bb001d939ffcac7b785f6de4fd1adc26424eb1995e50325be2c29f0105e26a25de2b02f0123ee50c820245ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8c1c3b0481356cc660ce59e614979ecea6a791619fb45f8a1f6e33e8bd576166657322f0dd442f397ef934b06920813b9f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e8fc4a3cda2c3e74cf31e32c5eb43c34a1003a0b8c4b7c2966f83a28ff37fb51e173602ac126b1e1b5df67adc5355987b73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf30921301b58ccf85b939898bb580dcbfb4b2c452fe0f64ce17443a893acf4333e035cc4bc48b4533beb2639bf1b1664b3f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbafb958057a39eab8b272bef0770664680322f54a7c716989bc778567fb17e4fc040a3c8ba77259e1448de35852cb51f5080;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5d86251940af0d4bf0e22ec967afb846e8f326cbf01092d0aad41ea17501283f45f0feb4d272653e652442450243def39ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57e5ba1f97f6d342973951f18d0c4d47c80946ffac9f33fbd86bdf25dc0957578edbc91f56fbbcd39715ea33ff715587c030;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h610d002d76e7c57842ebe4a33123ede89c753d45a6f35cedce47f27979605ee75f456407621aa1febd155f42f89cddece97b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7014f734305883b55da6b81228b15085adeecb35467791c12b65255debc84ca226237e72024593980dac5c14da8d0846de4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b3efa424183f3493a50b1793031e0db6029d0bf256a4d8d6a0455a0cbf27f540595418da2998419b63316f35de7afad3b94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h646d37f6a2387c04f905473fafaf31ad92005603eaeb64ee76dde4f118d3df653b916143337ae65135d0eafd719c195f96e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c0c347e4aa57a21b2c42fbd58171e00e25016ed2ed0b416896ee935b1c478383d19136d7072f4dc8b110fe3dc906e412b7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5dc0244599c029a119b8539884e7785a281b5440ba27fa0da6bef0056277e319998a46e540d464cdbf01f0946dbf54a85a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb36667320dba5f97ef19de49a09f4be3efd7f8a6709746ba31301b788a48e0d00ac694ee0e3b0c819ced73339c4e5ba75495;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7010956f0f664d132fa1cdc3220c4acb7c3841c0fa3a20ddcada7022d267b8bc2227c8ff081e3704c6578b3bb2ec2c09ff7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0878f616677ab2c810b1bd450edbd69c56294de185712903bc4a79ba453fa2591752d0f2f35c8c4d7e994fd728f5b2412c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h227ab17b8b7cd01b71ba9ef5844c5d7d40f6d8bcdba026f7ce3de73316d718efd53a7afb928083a902b512f34696e5fdc055;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e122d7f689b038aef463afd6c3c061483b343b98435a17deb4cb69fe03e423073c52ddfafd3ca268a1ba1ae460d7a2b5aa8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ad8b4121ab22fc36bc8447954a405850d00ddb339915385c4f1cd91f5937fa4ac2a9dfc87ae2263ff0e4edee1e8315467a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25ce793faf6c9a436530acba4d0da516a6e590f86604dab6915ecdaac8c40acac5a5fbf61f4ab04726b85bec624df1be5ee8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9aeb4e6c8238a56ebd214b98f93e2cfb0cf9c08f44b3dc4592e4fd6b5270bb27dc02560c3d10d8b03a96a0c7545eaa4dba8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc803b8efc34e111c59ad1afa63db1bbcf121a9138cc21f7d0e96e817227b2fe857031cf9f5954db2f32a0d323b09b200ffe3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bcca1253a4225ffbc5266065d38662c35aa847e8cd2ccd8b23f03181530c91adedf02b03511c8ca8dc7678dc80c67c0fd1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha79727cd3a23ac2a7249037ca549701cc98c9d332690eebf075d0bd7faf983b6ab84d062f1045fbd7e9c11bca3806e4d49e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3a5811f4ca1abf0616ff3e7fd0ea016fad6f30e8463138e7c10025a2511599f23b90fe2f2ff4089a5bc902eca147106d8ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c4fa91952be01b5dcbe5d3e1475aaea9b3f020c3f9efb2146f285b723c38738f05d34f39952a9fae52a751522c63c9f60a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd22010db20cde3332a2ac618cc0c9e8328bb52ee13e7c30f79e4707fd410a2b597321260e1df910182427e8e5a856362bcc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c12f0bebc2e93b1c3122f01c5e7362444ee4a7df80e8122b424f4c599d782bd572145ceb97170a387b0a235c0c379bf1992;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53ac9424a721133769cb33dd12a34904686dcc0a81648630ca2665731028013980b265d3b068504a4707b0cf2e172738086a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6762b2f43e272586d6624f61fd4b68b465d2f6d0e1fbe3356a8aec9ef534cc25f9943c8602f90c173ab0b624e547a6ace6e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a5e0755a420bf271c6f9f27d056973fe3721ed06d67c3358abdf39a4aa0328aada27f1c6969097198cace4dffc519e99a4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h595bf8cfbf7423587d8ef3b8cc0afba718aa5ad32ae0ffc4be1b54a17c29f36c80134baf6085bfc3380617d3eadf2e1a09df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54a74db81fb3b6f9653102c95c3a39518375c13053e0295024741e07c5c6d1f20eb34b33b04e1e5a5364ab8281461c361dcb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c3850182b0d8c55ad90840aa02b4950e874ca8365e8464a139aca2d665b234a9006f58d568d40941cb4bee6c3fffbc00368;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc193bb3d0f6fd2e8d9da6fe5e112a50fecfdd0dfe4c84fef888fc6f60bcd097d7c073997e3a2ba261147862e8596daeef9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfcdc67b3394ff04e8b7b57059a3277d02ff6d204aaaa46ab8773d4746b1ccc924d127ae977e39a413a7fa047ba565028ce2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab6a0cad9755162189ec2a0c06c06a5ceb88a2e006fe901fa9588940eb7776e742c7dff29c35a4cc3e59e2a4b6b2016fcc6c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71a796ac08484bb0bab6bfc4024c64fb46d8f1351a935c1501fcba2c1a1e8a9649d98d13dcc480e4d780add4edfd5b66fa99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85b86a4c2d53ad8022c02d10c6eeae826223cb4793d818b1ba73c66c84c34a8ecd84c4215af459602154831d7461af02df69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe5e0d9f120d8c5806da5fe77c872553fa3a27c90fb078f109ad71e1b2b2c0b3aa195349f9354b81cf1a8d12626bc45bdc55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9112a1d58b75cfa383e04c8d45db109d46a4270804ce2b88835afbedf1281b9228a93f8482eaaf30ce12e2513e592456cf1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ac50e9d8188989da10a9fb2b7450e7d2482287dc49dd00d43b9cec906d843c0c17a498ec6391ea99013243fa896b190a784;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58494a7e834782d92f806e4e373b3a5364c7406682eff277a322c8d9f5a1c8cd1a17c22d15ceb5110d71589123925f015909;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fb98efa45ce8262bb9b32238441d8d9224b924406cdb95b9357f7733cbc82983eab25fc023c9f94d89c91b5277d7a5b2aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5266c6a08d084e5dbe2a06ae79e07f432cdd5a73d600d03422b5231587027298f28f93a7eaf4efb77a33e79a21cae0fdc465;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46a5cf3b27ecadd7fc740be082bf0135794bfc6b36a51f9a4ce95bde74cd7ffdb62097a103937d88939e53959877a39e1a12;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71051a363bd71c604dfebcbc19bb55e2ab11cf912c6f829db3bc450549faf7193f8e325bae2190294d589aa27fd73d9cbc70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd67620bf29c494fded5169f98cab51b42d89610460b9578fb6d4e94bb71d6238724b9abba3ebdb69abf847a87ebe47627371;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54b89c2d9aa06376a2e2fba89cc6a96ad3cea70452b71ab50ad0e044dd1ddeb20e186a38b49fd14591bebb7afc2c05a6306c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7238eff192956ce6fd80fb0760f0f83ecde9f61642fa25efe39eeb82596534916052ffbfc6e7453cba6526971a16f0160152;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f375e31c6dee8b70c552b11ce4f6ff55905e4cb15041666030287267e1aff4eeba938571b33add8e75a1487970fd388f6fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57d0c8679c5279db6da695da6589ba5f10e7f10eeab8f064f137a8262c848fdeb156ca17faee32e39f72ce95c73922ebad2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7a0345eebe7bbc06b3627727dbab57cd069fca58bb8a0c69eeb24dd5f89dd08c56d6871c4e683b82926a74c8ffa21c537c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h298948d25367c95936bfa4559e974d12a260e84207522a857cea5dd3f6b76edcb33114c887ed23400615fbd38641ecd04102;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc96cad69ccc989dbdee6525f6d1be8d5c3ab97ddc3486495deb0f3877c47c0e58d2b4500999d4fb535a92b0241ea40170529;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb74e975c92575c6f5f044cc4ce1750f3a68499f763897b68af13a849680721cce68a43b581ee17d0660c1f3b4e904a52ae64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he20fabc4444460beacf55d046a97cffd53fc86c6158a2a9998a22fce6a4afb6e7d70ca56e9095585641f2b4a0ec43f64bc39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b907e40eebd49fd7153ba1f48b6e730d01efdf3d1a9f8a885af5dd7aa65bb7dd1792b4d73bbace4629c108af5e0800030ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdecdd78c19ec2f7794d8140783be79b3b5aaaaa880f30e3bdb0367c77e7256274b7c260f9502b9861c28b09095a5d8dfd1f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a376d9be4815838a165a6e3f0dceee42bb9c89b36bb11b59608b9abf26b481c73909c1746cba8be3424e32283bc14e09b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2484cf9bf693e0b6c467d03780e99012d8375c6f623e48b7ed23aa03e16a50e016cd17f264770c6addd584bba0b5c7f78697;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb343027ab9f0be978a3e8e1752490b3fa1e0ad34e8afbe8842559498c6d72b52f24d839061833b54e899ec242042153fa0b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a5a3514d7fbd4eff995b80b04ee2c47367b43963b49f4e7c40683379d20b549dbaf63e3f19628011791fca03f8d516733ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h817353323f007628d5f9f719b359c2ae8137274c6961bdfdaef08b869ccad8ca5346546c8b5dd535cc19430e68bfb128afbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc226a4ff47b3d53d1f3c13bb5d26b939c69dff041223db2e37390fcc8b3f9f628ca49e4d1f2cd9b3b5a170e90b68f7931cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9af3fab867b62f3093f032ebf0eccc6ff0025e76282e24e454ed1e0cc04cf54904c84d10b42e7afe0eb48f0e2b5386451c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19e6b2a9ba5a4c3a90afacee8f174dd13f8954acb330ab50a26d2b44c9ac52634fc1cb209d7337755647208e0ecf4a9efcbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcec99350d00b60a20e934684263ba59e83cafaad2b6ac5907321ce429c5ef2751097dc5a4aea7b4d7f8012e7b9c3bd1849c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc27aabcc39e94b631cf89286d23bb17e51a377ce9c210c85c640f9c3a655d2441828e1c6a019b2810cfaddf29a280cabc6d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3646b44528f5b5bd0966b1f3e755e3ba5484e588e89f2559bc7409383d2cbe39ab372005e503473d7f16c6457a9dfb1498;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5654fe4471747c417dcb63112e010d25d11db77b3b8355349970be7122454f8a59f103a6960f940836653c7dda2aff90fa4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdabb66c975fe8bed12574095acf5bb3ac3e134cd738a6293bd23f739f569e6420f3246668a5fa2d7ccb80e3f953b581df781;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h468e63fd6690704f71a848db3cebc2c6996112a88c5d7478139100155b7193f6ef605d0726d0c8b6e2e49de3a16906dd5a6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb84505b99ec6816bd5f4783f0fecc5f83b961e6d6cca2df8cad284a249c355bbab7838e79fdd1619eee3cb022b1324992cfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89d38595a84ada64c135e99755da78f1bc3e0086019af0f205d8fddcf7351f2f942bc3363c2984a87b11d6025be6c40dd8f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4825b2cb6c9e86ffcd5e615061414e583c6c7a39dd1c9b32a71e8099649aed432584c7552464e4361fbcc735d48dc011faef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf15e8ea1a1210ccd7b9fc20d770f9a25535547e5eefdba7bcf2d76a4354f7449c69b4be8ee7116ac72db23f2e870b66b34e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3588c36f823dea08376d7eb3fc2d92448cbf8a32375ebe50a1009af1f6e8f3f6bd4aa7089ff37f3aa9b27d1da3c848cbd6e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57b855bc187913e3b6e05bfa894bd37f193934f1b666f94a8bd25891befea30ff3c527ddcfed5c0b227f3c7cb4d86afdff87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a169a86c1bc364e86f2c15d09bfbb51b4f1f42201071ea7fc0961b8d38f9295f46a724df7cb5a8c81e0eb27d819c930bffb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca084c636eeb63c43618c49e47d6bf2c95325538e81f9272f10cdf980e2988fe45639fa6e1c5047ad273850b57b4b2f96e9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22c49a1ced2da5e53fa36912321ab4a60481f88ca8c7237f84b50048a1b91ba9d836613e266adf2d76e5fcf824e012fdaf12;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h886b0036408bb16ee722ea8007eb3b16d1a195fbf23ff2b59a0234688180a4c4b6602deb346ebdc605e1737bb8115777ff15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h735471c86bf1959ec6af69d4cde12177d64cb717d45161f0f1dfd220de4890afc0812bc035be008136214eac3dc81d0beb08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76c3e0bed07acb352c30340889567a7d0800a0ebb73800df5a2c4c7929478e3451c02fb0f70ef195253460c422498d59f456;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8321aebe9e1e6fc1ac66c10447cf1fc379f13e4e9d286b344fc060d4efbd2614ce354bb1656913403576e80712848a75641c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64b799d6ae3e18a18335360d1b59bea6985f6decf5faf1a599b982467d6d4e946d69c2990d0b963237defe9f8ead185040d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf808150e26c250d1ca05c65261830336291f6b8dcc3aa9b8036ea29520a0932e1bd704644d9eeafef0029237ad688725127f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h480709ca1bf82d7b9bfed3f79c2ba5f3a1210bb46f102f57e6afc4df12859f3b7827a6c5a8dec8f800bcccc60116d888846a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha90008d01550bb7b6c49237972c0fd08371ce7a39c941f28112812dbd417da35fcbe376d00fb7278bda103b2e7ed1182c07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9822629553aa9b31a2d2d13841b23546b1c7c5019ae51d21c74f646e716dc7edd603a0c8013ae27aa895748215d7700a34cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38b89f7861f3d6c448d014dc25886be5bb13e54b8da248645ed60839e9b4cffa667961fa4bc3abfa00dc0cc5892c1fd63076;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64309d42b7696bdaf14c9ba934fb4eaf5d5ef052af287f525ee2a148f4a341b1c082948e03b35dbcb4d70e11675ae16fa9a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89bde74d462e12f13799b8bfd672bbb5bf64419dab782437282b07561e3b381b1dc94e295eb7d9cf7213ce770096171232d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3639c2fc6b0ef571f69d93c1ec8cd66b9d89583c8da5525f5688982d8595e5b5c0a258c8a6c11b90e0ddaab2ac4390665d85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ae9e4ef6086447e6c49280c7a1bb6e9b6181ddca6adce03afa19da9cf38510840612d561fe6955b92da6456cd56b849c220;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2fc18412e3757f8fdcadabaac055006eca90faf7ea7460f7077eea214dc2503f7ca9ff05d29c3cf2c03581ecd3872cb9c29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5372194c604e2ffe6d83b6a0cf62229f2d7bfa2901e5fdbe725ab75ba0ba4d1858cff974bb43919407677a29a8908805e8da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heab45bd48563510120bea3f44010eda91c4f9491b0c9d008cfa34a62272d6979f412fc9ca5c4b95aaec34706f6eb554415e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bdd809140d6625180ae0ba3ff391ea2277db341ba62047581b79a358c3aed2c90db8e20b4f27612f4b796f1e21771353561;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83a858c6a98af57f4a656ffaae39da4b451bda40ba73f0c0b96a1df3575261e9e1b346fe805382c1326f54481ed89d4cce86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h744686ad121899aa98f2db1a692dfe6c54ad10f833fde3b543e1d5458aaaa9deceefe54ab651a481044358bd590776177543;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6673b6b78e64f670c6ff509548b1857144ba0aa82ad3e624fb5f6f5e69f4743f6149e401e97e8a5718e505bf48f41e480f14;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a4b598ca7978350b5f30a8c560fece39b3b73f6d21935885fd25a67b39cc655cbb6a21da212333acd6fc0802c90cb068fc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd88cf98b0d95c36d2ea2ac08dba9900689714e57953d75b936d517dc0ae35b3d671162dfbdb3cd2be143c8d1efa880868b35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc2cd6bbfb565fefdb0c78ee434166b9c51d2785b10118a2b5c11296cf498c86f86eefbe87893c3b2a627c664eca55cd560d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e561b94d15bb916f38e57be98b4dde616e1cdf2bf5ca61b6a70b2f2416eb704ca9cba0731df82a0c8791bab79fb0c29db45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7690894c770dd3759caa9b8be818def23238fb7a767dfeeb11db57baa21e2d9bc7bbd3dbd23c97795b79cc6dac1217824a22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec19952302a63bd6756d17e8a31e8564a747c9ec903c23aa9c5b128bd59ffc85444e1612c8dd3fe4c6b85708dccf5c1992ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h470d9c816ced43b365f183ec4e76bd0a30c6a68d95ad6aaf4056c7b22ecba697902233f5a73432cc9e64d1778c0e58069e9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13e78e9f4f6981fecdb44dca7a2d8b19b638181e8ccb0a7afb9f05bf41365a9e1f67c2c34d652c1837737363deecfb6f6ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e9e95fa3dfdc649356402ec7f34c6748219f2a5c244fb7a8c4f357feeeb0057877eea62ab71fd009aed8289e14b67c230bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h247bb43acabd0f3056766e05ee1cd1b191a993d4afe8d255780d5011b69a08368e0e5b9d170f05e45d61b1c0f367c2d2d9b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a4072b79ce3c5d5672ba230eb1462fe498146ab5e1766a9b2e25d82fa8a02f6e869331ee424c370a60815782cf57fc47c2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ce3837b8e4a41a1d0c34173c493730c482d03a0f9de9008edbdff836be10676d8a1a9c118e09346fd5237b5b9c757def727;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he734917ddae3578eb3b725eee33f4b774a0cae7676db586c767598c7c7bcd62f3b996b541a3306695ac0b00a0b06ce76274f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6867eda89109e2964565b900420681ea201afd9c29b63b1acf825262bc00a1cb26272a24feed398efc03a5a9c7b154d57b80;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f41e946d442ab1cd80dcdd38b102c5d5406e49ca171fd871c191acfcde7f6d3ef24aa28e1dd7833c156f1353e58cd4fba5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b1a7b7531100b0fcb2ad5db3a545ee98edf99044c3ca87d79faef93d0f1938a914c818ea1a54de80332c5c2da887b680b86;
        #1
        $finish();
    end
endmodule
