module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h386cc500c6b10e3cbe594485;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38c31bc1170eee762ed25974;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc973e5609abe0f36c60252317;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67ed87a0bca1866f8a8b0520a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7517662cdf1aabcbde06446b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8de5a514442e1a0e5bf1f46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc98c20196d714dd25752ab03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcd58bccf01dcc75501a3000d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5641358e91a961e152157d22f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f0975c77a8a6af939e379e68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28ea96e8d05813b9a66518bb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7d7d88710ac0c01a64a14101;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5b362769fe80937bffb96dd0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83876f59f22cc73b14b867407;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc46958e636ae5a3cef06404cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46b3aff612e0f6b032b994326;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a11614a947e42c950fa0fd29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50c08fdc708b75ec19ff8ce0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdce4d19ceeffbecc059130fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fe1c4f9c3ebdc0290f5761b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12c3a50165ebf093062710b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87b115dce052f686ba33197a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7309e1520f56e64898ca1996f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70f121d23e43d5386ac11332a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99a508905d751241e99b998a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d0e1965ea9cca0b133b5dc98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdbe28d1f44ecab2d491e61cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffdc0e9199119f38833da472c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1b8da8fd490a99919b214b43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12339b6ecc827f8ee78732c3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbf54c1122c49d9a96068ee97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b0dd96d058d5587fe807e336;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d7d83f858597abf00094ad4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda08c4d93c181337f93d0b909;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7587c54fdd02e4fe5a33bbc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b0232e6db82ee50f40c01e4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba88e5c224f374375559e709;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6a62be2760e7b6b64b319a88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9032050d80ea77d5ffe02a5fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f52b04c1e0b9c5789ff8e8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h266dd245ac402496fee976713;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7c109b0dfb64260204fd8946;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc98065c70b4b4170a10765c37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90d696325e97b95c705e99a87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcacd73716a494f924a2179d27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc86ab1a1055eedb66c75a7476;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e99eab58a30aa42bf10ca23c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93a4ce86f97764750b9b97f8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4a4e324bf59a6f856c6ce56d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h142c87fdb62719e09ea50e792;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37963c6803502bc99d47f0bb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d76f6f08e92f573dd3c59dc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf99a4b8606461cb8d33cafd58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dd7d3463246bedebe57807c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd490c10f990a812b33736b4b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd050a5dbf8e69d86fb2b40cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb9432d742830ed60afc9e4e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88e4abd8e6190e236ebf4863a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h231b11693ca9a88a81b251bd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30abd71b3f17c6d47b48afec8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf49e5a8c7716e392f57fc0c13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h658026edd9bdc0c14b8eac7b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hade551b53a37b2a2fb8a5e1df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf074ac7b74437204d127499d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc8129a599bcf50fb79350947;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb25064409bfee179cc0f373ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd1ea305ed6732fdf94f1cc10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef7ddddcc46dd30505bdcad14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h239a9010d2596b0199b677859;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bc73b02fb0a4ba35d4562526;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d0a8dfb7e575dc6eecb9b44c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefc9e8024c76bcdedf4eb7a14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb552ba83c9083c57e2f95a7c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h562de5d312fc2311de788f207;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dad941e579e7aa6e07917c29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4d0744b029e95b9a37f428ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9062fdccfa0e51be6f7bccc95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd5b6dcc95f71f3af0e8acb0e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf17fb9d2c00b93268463e4fbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb2ca3b444f00ec6a9440ff2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h792dc5d013dacd76df0b35011;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b787afa7a378f0a1252d600d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb413103e23c06b4ccfcc684b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a005685226dccc9b1694fa4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h692346bee2804b0645eab6ae6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6481600f0635931317f4ada2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e6ffbf5b15f698853fee30bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h174b318de09631fe24e56a4da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f9977171c5714a2b5468b2a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h366ff72a0d0c562b4cca66762;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2d9ec25055fa5bab22abfe4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd865af7361607fab188df2389;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32a299e756fdd4da59e2b3a06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44c773f288535bc4a0d41d0ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf91d1eb34ce2882d8214263fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h705a621fc136f3efe1e74db96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb488caad96ef6d3762d8ebee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62d3d163bee26315bdb11e32a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80c3188caa95f81d6b08e8a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha047a34bf20fee9efd152c043;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd89bb74b4781e4daf431bfe0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf7fee6776af5617a7bc4c0f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd70f6fe7a3d1ce951aaa008c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7119c98257ba43d0fd4fc1f22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc59d4a33a05759fdc1a92b56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4185a59d4774b75ed086facf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd90474f0d88bfa5143a63f62a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h642eac727ccfce6b7df6b86ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd6316c2ce652887a57a0efeb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccadb4234a1503922e851a823;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0cd4f8a705f113da9f8ad364;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd45e8b8e4c1198d4cd3c3e8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he844e658059895b204d1707f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1eb73171ee70234b568f4b6c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc61cd9cf1dce9ef0ea5c8c228;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8244fc87cec271cd0bc1e2a8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43f38d95aae3dfa32bdc524d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff833125004ce5efde6741a25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd807700a2875a9dfa2d6b20df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a076d3026094415c7c4baa61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1f1ef7520c14ba3665c802c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9af11fb13fc26f68944253b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43959e652c7deee5c84eda771;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62aff08ac79b4b97188ebfece;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2e1fd0a85b503a99839f0108;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd6c256397baa198351afff06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17215ad1be8d2fafade9f8bfe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc4f2c7b5296f88cffe9a22f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16a329e79b87079d6eb6461b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98a539282a349d95c5c4ec469;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ca9d960cd66dca7fdec87dc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4f811a3c6c0e83e164f30dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a7505ad793103b3fb9658890;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h195f8ac4cdb3540bc4f526e90;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87a77c3fe542fdd9eeba6b9de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79242293a2b79e82d65fb58f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h980c52369f70b30df35840c4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31b4b6e5c121d6ef101f0ffeb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3000668baac85e1c1e4271841;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha93e46cf9c4c61d22f0c788e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0f3bb09adbf2e13419fa3539;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1ab41b44df590d5a3a79a308;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c1b74b9b53934769f872f429;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc06f54910c4d7d4ef8f22fe26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h853fb40ffe4774ead6299dd73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7506b7cc1b7e5bfb06da71ebe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fed9393efedcae5c9211ad24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed2f016a8884562ef3c27f49b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e3eaa4f3ceb239e516adc86c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7247e2b9c6eff8209b18e751;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbb0a5e6c4dec95a4e003e0e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3fb623e43ebe8caa16588358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59be766ad63c8ed5913607334;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc02a6543ea7d17d02be35651;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf7e1dde7843c92abcb78e197;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h324663d70944e09ab286772d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h154a024847645b1dd83062ef6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb04a36e2a6466be2b14495d98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4de9f06fbde8facad22e677d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f27b865eae5c8b31ad9ebf48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69ffb75ede1f879ada6adb66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2156759a4d961e2c00f4f8098;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c8ef3779a67e811c25eac552;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f2101e16e84d9076689d884e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdc65549bfa23c7a22cf1e194;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd87a168ca90d166c70f765c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86ee83152ae03166a1ad8a155;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32d01763f875edf21453a6ed2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h456a281f9d1b0f4a7ffc9b8f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e80a562d0409ad5af47c118;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ed09fc6f0600d8be1c5f772a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0e66f2827e2a791fadee8774;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb606afdb1d3583f2bcbf5b1f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h208dce1b31bc65eb245e40bf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb179cd2781c5433a1b6ba5bcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6137b7dc052977a881c4fe630;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4ba668c386dc20be1cb37a91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h936dd854e169e0920020707e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cdbf6872d75dab7fb6b59f3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8d9c5a92b649d549ef02c3b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5aa49b5b883a0b98e91ae19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0303774983a1af66aa7f58dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcfa8b49caebee348ce8b231f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63d0079ac7fffe1cf951a9166;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h520c9c558b95fa819f5462371;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e80c6eb6e5bacb031cca22da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h377ee9dc13314cde7ea79ecc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0021c1ab280eed3d9071ba09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ff587063dafd0d733787fb69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8050cc95ba7515005f707a01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff19ee254f9375a4d6df5e8da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd01c2a29ae146e72bc24b506d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8e764b362588d6420a3ad07e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h799588ab1dcfd7d9c2d852579;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a2808df0547a20fe8a6d12f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4def9425aee033efd996895e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h103fddda725abffe8cb77b936;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e68a2c56dd972a817698df76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d6afdbf19b9d39520c729c3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h596de88ff99b6120229c7b897;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7349d02270db0f5e965e8733;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a219831959dad3950ac93af9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6027cb692a7290167dc146c04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4d3103b6c82bd038f7d68e12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he531a7212052854f82f08ed42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63f6bfce325d1ae3167e90b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb2322073684541592f7b2db2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd820d089bd631392211b2fac4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h778b84ed1d769972eea957ff1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8f203089983be1f240ed073e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67474d5315940477dc46047a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1553b90c4406bd78185dab9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d896c9efd53539856ddaf153;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7ead1ffd745c52de91f967a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa8156c5927829849beb53cc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d4e4870934070d43a6978d05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55b4592787e862ed46402bc38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f6d2c128d7dd7948d14e3dcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38d0e8b5292892b993b3b48f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0e5b05cbef70772de4e7158b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38085d6379e66ee429e84389e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habc4c5577583299121240010e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59b609c8328672cb4c9726eb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67341250d0bc994a92269eca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1fe1646cf3799c0e129cc616;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5d7b552af2c774d6061b32c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha76b7cd26b690c58b19f04fd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb11487dda9c9c0a2a4ee1baa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0fefea7545c18c9439e82a36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61c888d621e7cfcb825ccda6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32f87b24df17ac5895c834088;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5aa0636c9c9a51cd2e5ab79e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc138ac23ee5dca51126cfbda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf37e5659ceab9c26479ebc709;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3322432b118548d20116af82a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e4b35abd607b22a52e34a54e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h626a401d2107aff4aec31530;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h284c6a94994715f53b74f0e32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h779c633af154ef13379687b88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he42c0c5650e3432842d7b06f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he811868acfdbe3aed6d7b133d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h686f4171dc799409f68ccbc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba3a3fdf6015a8d2f4e13b7dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfd3746a1635ec0591019eae0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd373cc61376b8bc34f347fcd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b53fbaf18fb4246afae6f369;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4842a14045e81074cdbbfd60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5453e29c0fe6dbc5a67737c28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he72b69138cf3ae3e7c75aba57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d96c0b09266b58182c27fab8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90bd305c707313f0f1f9ce9b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f57a45314e600554ce0d32d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h983052330b25090011bdbf6a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cc3bef288d5c2d7c3d9d20c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h951fdae9c9a0672835b5c4fe4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e10d926fea2444e6ff9d3536;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6db29b279aa0987aaf54c2d8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5cb8bfba98df16d9303e3e0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93c5536a89712b0eb4bfd00f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb65aa9a966b0f06f25d98c81f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce07691dbb518e8f7df5f9ff5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74805c5de078ea59a58a84bfd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fa0c1edd026cd9fd70233efc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf83616491127a6ad9d2bf534d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1233a728acce28624e964844e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42e2d8234bbf41a8425f343b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6179e1cbdc05796b33ef7481e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56ad12634ee4a8f98fbb4e29c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8373d4c22cb996ff026a5d24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60151b55f1aa839dc2dca28cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd15a0ca29ea421916c84299fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf932d22a9f555103fa86c5182;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h372a51e2c8f8ab5256459266f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa20ab75a7e060f987c0bf4b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd215028dafcd8e73bb5b88778;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd26ac0e20e64a000564a5aa7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf78be646b543bf816c6de4b3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd03452d6866407c90200e3e71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd181d00742ff689de1eef8af2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2717cf6fe30bb1a83a88aaa57;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4d686eb9bab48b2d9549ec63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c8fcb077b54c63d84d16125a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0b3b6db33bc00ba580cd6a18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f88d3cc03d1af6e12926f0ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc785d489946ca83da68b8e42c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf802cfad6a136ec7f4261d36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9c444666d412e219a5e6655e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb760711ec86e01dd53d2329c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a367eb67422eee7e1b21e3bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28a1402d44f58d3d7e4ee3a02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82a4a2cb2fdde94e2a07464a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9204792fb0c4cbc048bcbef3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95b029d55a3d94e9483e7edb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e6ecbe77b3f5d3ce7e3274a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f137d87e173dc376d664867f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha71e0b0cd04bdf0c405be2eac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf9572be115f982e98b10fe7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec0b3903b11e750883d1527f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7545948b430d5d8b8bcdba43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a947ac36a04ea3d6b16ef97d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf40fddcd832f4ecc0661ded6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a2d1d2fcdb9989efc550f98f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2fe9be02fbc6072c2f92a4ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcb0560e028055ce9115b08c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d2baf58fb2c38326bfa091d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha40e83d4e1b10371db7f4c58f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8dda2b65865e4430db260b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51caf41f0beaa20af9051b725;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddc5ce51860681e9ec85175e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7016bc25f5499693d57764b95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h899dd44bf9205c7d909a0b92b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d2e09fce98141cc56d3821d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4104a376c70c45583318c080a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h175423053f2a0efda8dd1fd56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2873f8c0ac46a285317c2ba5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h739ea49843cad0fea3f088f8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9a059213c7ef4fe61f0af03d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7026a0c115f9cccefe3b67ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafe9b962918e4e721a8aac439;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9e8fedfbaa16ddf8a6df02b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69a0527d55317aef04e2c2b1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h580216c6c13fba0cb252f1ae6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha989c9a54d26a5d08086b7207;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7c8a7825cd6b1a3260c27c40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd474ba49c9acf533c7240f13f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7d42ebac97ecad66876334;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55e7b10ac772b3f809ab29b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd46bf7a7cf0598447764d7545;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d1360a48b39fee3d18b463ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc86ce7b0a734d517dd14d5367;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d78691c5ee85b10ce476d5e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cc9c83a17e410e835fce89e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59ba2b3d9c8c1754b4fdb66f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec25f13aed34f5c932fe9692d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58a66473ec6863d3aa47f9a29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67c8d0cdfa7f5880b5847d313;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89f33869fa97a14e993ae637d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha13da905900ba87fe7446004;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb3e1991fca6adadb6b67b6eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb4cbb6de1e5d706aea4652c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb21da42041ea6be6350dd998;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcc13dadaf404782e86f276c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dfd84e31f6853e0d31a99214;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2c12107d8774a547f427b7b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf98e854cac6d55322263b5c75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a9da8bca1a42a7c1fa4c4622;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec1c1d8fae2a9ee42b49c2832;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cab5c18fe7c70f0a6b2f1896;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce3ba242433d35770ca2be6fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31da0b463984201d21b82a147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd51d628d54f9f23bd6674652;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b55fed6650a9cc8ce3f04068;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0875492abcbbe6a3f603e144;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51049ec92973d5237c0003678;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1063853f9ff673cc9bd875c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h542c3f35dd7e26b7fc2ce4ac2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce035665defab25cfc086fca9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75dd2493b00430d050b1439cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd59366b3ae8ca1d56b9f0ded2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49c5f35e00ca128e6d69b5e27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1f27665d6b238ab413d79c14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88b3bec442292345997173ec4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93a24ab291c28ce561dd4212b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2884b2f209be9d59738798957;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadf756523c0a038022b4edee9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf900408d1653464b7c6c0baf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa4a116b79c5baa074c82bb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22881930b5024c53eaf1a1093;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d0bf15ec6ef63275b89d6750;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29583768234e0fcd67625f9c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94d6d24e324c177f07a0d10e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf257c5f1e9bedcd2d4bf109f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91a5b2da5e3d313793094cb29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dcc8de8891c36f0994af4ed3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6f8e6f91d225a031069b486e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8ab1e61d5fb4dbf4bc53c78b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heca3d91faea94fe8b44649145;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1140de3bf50f51868905c381;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf8dffef61b2f2885ad07c880;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59e5bad0fa9d32f69eb1c3f0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f23ac20dc0173dda8740ea55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6aeb4b69fc4b8e0669349c9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h834d1d59b85b453f66179dbc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3b68fa61dd9fa2e688f313f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf625f57b932ec67047e69cf36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a3a1a014c0577859d179045d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h536d36a22d686b09fd9ce7622;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3cb7db394487a1af8568643a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeef993e70d353faa04278897;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf000793830a603d9ac46e6fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58cdebeabaa9e5222bc5b811c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cb7344818dc1580e310466bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68e0d521b05ec5ce5871061fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b3749437a166fdad5697d13b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc37efdf32f45f739ba9b4551;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a332c8675b2a27a249f92035;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b1592389ca8195c9fbb0ef7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d48456ed357887ed5c6133d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf1721f106cef5b5cb29c5b25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8a71c64a589fd20ee9ed9bc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4624727ae45e8c79588eead96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcfc8e7c9f50936ed3b12bc49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf3129f7f05e33b595423084d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7dc7375c64383f423b9fc14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h900ca9e69bf75e967f5408218;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61d24e71cb25dc99129136b26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0693c4da8dcb54b869033c02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ccd5b7b509b0f6e817f54f56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81bcefafa8cd96a3ab0ef5e2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2024ce6bef06425d09056704;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7a12196a6ed27a44ecba435a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d2688da116bb7e42ee4adff1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e6e9d933e4b0ca14913b80b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7272b8014f6d3c3ce0388c091;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e1ac820178c03c3d81087662;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79324bdac4d5b23cf1d2e0b4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6d5370f27ea92cd77c1cd222;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf17800c0cbd93e171ffb3071e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a484e8828d6faa5e0f72f3f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd91f6544952caadd6d34bc1b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70fd5f282986e058744aad0e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h117dd7e0489f26e37540746d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h914eb2762621d837e8b8e8e84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53388317ebe6423a8fcf218fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6433574ee7dd50d127e21cb82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h827d2d37b672256b51539415b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6599c8c974934bca906be2da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14c59e22c7e39337df035c8b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9a4915e81d675830ea389a69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf0997b1451525cf6835d397d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb905b3288913f01d8b73ebdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85435a571de15e1489db587a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h291c47907310d0e00a126c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee91da8e3e7b0d7dcf0960bee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4b293bb09093dde0dac68257;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ca1ddca697ef70e645dc60a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c01491e0b3c16428ffacb972;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf6e8fe7a5e6d58105766b508;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51cb3ad36714381faca5ff912;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd59fc315d1ec5a6f7f942fc9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13069d6a40aed58e922977468;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haee8df92dcb6e8d11bf76f612;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h201eeece5ec1ea22daf8cd73c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a3a970db07429da68225eaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h120aadd50998899c31eb6e2ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d1724354b11ef772b810e148;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1122072f0e47c77044baa3ae7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f84610756ab9838b8fc4f932;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55d4d2cc519ae7c11a5e0488d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec6d62bd3f6fb8cbe34f9c78b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8e7a2979f4d846be7c446857;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9ec623f19578a85bde1ed64a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0f4e880a64a823e6c72c99a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dbe054ea0e75381553b3bee9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eead66d5214f7fb9697ffe89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h398f95ab395dc7fcf795f3cbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d4c69a3a2690849f41d41097;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h986d8510a84c661c4ea37e8bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7631136bd8829222d58396aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1f4da3b4280f19b55599aae6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16878793282bf9553d62a9c8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd79488a1f2e8480153147c489;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44ff0a056478cea8a7d17bc17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf68822786b89b16972f2d7303;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba4aed719ee42ec13ffa8200c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5832e493aab7a42005baeed9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb920e436f862c0f05052f433;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he38685c02bf4a7e1be6c1078d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3418d40957917d9edd4ad436b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ba9e9ff1197520ecaf97a179;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a1dc2d74710294c509de026c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h795f6bf77312d2ab4ec0a9cd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17a2762e9b696c737b98dac1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba2881c6f96806a2d7fedbfdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h894e019075bcdbcf0140b1c9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b6f0cac6051790b345202c52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h106c8f89404ed5d143adb29d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9a93715da9b6918bf965fa00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22127158e5d996a8125d1a3f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h512c12a8b1d66e128d6b13d30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec7cde8ec80b9adf52543c2ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5aea4e0f99d2ba4252e7fd55d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a326f078c0187d718213bc29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9ee1c59fd3f8496049c50811;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2005f2bcdc635b4eef5ede06a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41ffef1a8cdb5778b3463d914;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h739a1cd710c9ba6daf09f88cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b96c0e2592a548cefe111d1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2bd4e96dbca3df2495f78b4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heab9fcd4ea8ea1bb257b19fa9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha728bba4872b4122ef75c19e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha838ca1ec46e3664b46ff290f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98c09d1bde269e3f6ebd25fe9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdb9dece74b76fae1a85b8f99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0b4aa626ca45c4461bba34b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7058ba745879c54a68b671754;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f906e7e1df12879c0b04dd03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0fc49bc1064927715c6dc19b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86668814006f11fd45ab07ce5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4683ac482617119fc175edc4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e394ee2248a2d7910d23e18c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h385c556753c7804a611827308;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd9de50fa1164648701661e0c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he103b3955bd9b55ad7aef00b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80001c6b1f6295b41999d0ba6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc5db48dfefe1400ad8cce554;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9b2561fdd321d42672c6cc59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4809af0606c7b73c462416d5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a6712df796a32b3ac0dc4cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c11e5cf9dce71196a6dfec7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e79ceaa77ddc7a42046a841e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0203fee2e6abb0d0b226e5a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaa3dec6b5bb0c83dfbc75db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb51f54a36d4cfa086e458cf81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35a618e91cc59bde583801261;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d501de08a0173765cda68b45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50d0a483f37f604e2314e99eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a94ee3fa1dd5b01994cf0c16;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10154b0a42e37ef649722c378;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbedefb5b53ca0e0780f2438c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h630ba841f0ba38e1ded103e7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda1bd64d95e4a21b5a763d7a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h444d58a5becad347cc67f1206;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h545e7e99a4148fd640b8e35b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd70b339eed71f4cac05e6182;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h514d1307ed9d6fae6664c2d1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3d30821510aced9abf227760;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6787d9d99bc5cee6c05a520be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e53ffbccdbbdb4348d35bb4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4da4b956b737674620703c4cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23a976d6d6e7d0bc69a05a8be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbf28e76bfba1ecea0b6b29d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde2ee4e2a6d8f678fd835e1e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a7ae0e65081ecf32aa2d2c47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h351a207d8661bdea9fe72e1fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7565025960422023e91b266b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha40f4e25ba87c7d68a9a61b91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86582d1cc4679d3c48a08760b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92f2d0bb6f18076a8baa8cb70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52378171b9e330f5feecc6318;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h222fe178d0e9a32ea0eea4cd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h359b9fe02584afd2e47ea70f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5a475b12db06d048f3af4cfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he545c43019715e6d76a4fff5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8b2d4f199f36acc5d2e63d8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8020f983848eb689e986f1fc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75a584127f30aba67582f53de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7ac3663747d819cd33f8e39f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9e496b306dc9b65473d799db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca0d41539d706288b32ef027d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcddc1228eef797d60723391d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd80622fa7acbd9817eb7c9e2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33b051b85be72a687fd41d6a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fc69f7b7134d873607a9a4eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haddea3b96cf8a1e50b81244e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7c4d66aa3e232ced91f0f643;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7d656d515bcc053649943838;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had94286aa79bbfea4e072d702;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b4d8329e0a9c7f3f6f815fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he238e4d3e367d775e3af69010;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97a9903d537e7d8ce3676b42e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c54fdad5abdd06cff3d18a51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30307f348be27625badf78c4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4514b78953fce784b01380550;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc66bfeac06dd52bef835b4419;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fe9efffd198de8d00d15421b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2a10dd1a903c7c22ad8b160;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88e893c412efcffd252f4061f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b63aceb0f8b312e1037cb239;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h520537c76d0974e0e56bc24ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefaac8bc15510ad7932ce1523;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde4ccdc164361a7effc0b0724;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h986da46c7bb9c4bee083f16de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a821588fc873299be866d131;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he38d01a56c2bc4ddb77e563f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b169d88daa097741dd519804;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cf2ec749f50b73f82089ce1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46090c28e09408f69ae43f09e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10628e8cdf45a9366bfc8f4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb12e4833472059602598dd19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4c2fa619b0aa425cb43374fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h523fa476149e2655dd55902e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6882893043ae234be4e5cc469;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h202738a6c1a1674c1d3d08188;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2363ffa056604fe377e914c33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7a55ba897a807056cad918dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c8e06356266cba492b37d24c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h365dcea1b715141c8a6889212;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h243fb4092df5a9d344f4453df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d24cc24552d726a36f87313c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'headd0455bf0827dddf62bb2fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc03f81e04e3ea6a1bb4f0b56e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h210075ae07a2d0677bdfb02b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47d6cbe5fe7eb0a9b4023afe0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c0319d8c66c77614b7f0225;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h391484bd7fb52de818e96abe5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4360c199f5d3204361cdf5570;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10ebd4844913aa123c4b4d793;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7738c13c2739d9a170a0eb227;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3b41e17d35419c871cd81c2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h294784c7e8d2a807708aee34c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fd600adc74c0e338ac3425eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6a31051f2552a6fdaf070089;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3c87a4b59ee63bf9b6fe9bdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a5bf1bab7545cc1210967f11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6fbf20d542a81fb9b9ccbdc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h342dd54b03b108c143f8d301a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28b41ad50658a6e824f705c67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e20ad2d55f94271dbf17ffe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82062d604e1d3343cdaf27403;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda8dd29d9000bf7a3d6088f64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fff4bc9f7d300289a556b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4052ceca3f98f9797213ce61a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h589157038512ebd8f47841891;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf80cee3ccb9fcb969585c01bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c2e4cce4219bdba5dac6c50a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h773b3ebc5fe288c7de01d6d00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f321d01936f1178c53a26763;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9180b2d3936be6bf2a20f73e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9b524416093435d2da4046e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a6c072dcf6ca24e374a35ba4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeb42f117a4d47534c027b621;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e4947d5ba902348e02260e94;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bb76733a88c27ca92fb23e59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21409a7d6e50c4509770f9be2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca3b6142e310bfd4fa20648e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ecd28b818bc4674eb805e271;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6d6ddd8db915615c209b8459;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dbb9de344dc93c6f336b15e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3383688fe58001c1c2a740e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h818bae50622b9ef079c98bd2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ee714985f864d311b3a5d0c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8a8cf1eab92f350926a7aba5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6332692583f0879de3681628f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab873d007987f44f92e83e98f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f6a53a61976c7310402f89d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b18bd6ab160d0d5321133005;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60e001e9423732d59e0a70438;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87c74522e4a854b756ab9d221;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h529ac54c0c3d792cd2ebe78ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2eb771d3b20edd526f0865eae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37495b75a9af4c1dc0275a09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb25f00e9525fea52e118aed6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4462d069a86b76bbef12d08c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0bdd544d3b8f2997f2dd7af0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h607fa8a613ab10cbd71abeeb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76e6bb40334481cba55eead0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb30f05d8535ffe5599602cf33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2b566f6355581896abfea437;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcee7ba083890703bf7156a725;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h658942b3aa08225be45dc16a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb1bffba5a9cf1b316740852;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h640f44dd063414ca077e0f227;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc93e55b4a769bad49325a2b65;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3ea5724505a6babf0f2f8e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91b80e1b64da7e4403da3d05e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeecdd3463728e72289faff8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ee9450f57f562e3649edda2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37c743292e525e396b44d5239;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a4f2c2b54c4daa94ad90bbd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bf24f7e7988954c87356c74d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fb9b5d3c2b49edc4c0b403ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fbd2492fb8630170d44bf910;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c02f2859388c1d238ad12a19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f64deea3d9f64f19c7747f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3945a8584b63bc648696015f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91f830921bff7a6a10023ea75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4ff81c5dd847c5d93409cd02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c9e0713302fe59dffd82ab41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5e1b9af2e87e96a380d7793e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a0b76287ca860df560e4817;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bdbc36359ae96d2d4e1f8167;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf74e7e7cac3c6ac8d796f8306;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcc3d0b2ec6823374c372351d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf55ec94c0babb90729d818adf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ff3da8b0cf868894760dc6c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f48c055c39975e4255293819;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd94f315eb5bc4c11fda55b35a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f2272e8f87969b66fd9e056;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0d87090d6b7030665557948d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he977de1c81db7eb27a89157b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b7a940892ff58c40282ceb04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9599c829fddb9a50c713428bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a21a8c4d1ebba33faefb616c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d298f2527a8f3d27c64e462c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3ff6a4a695e07db60cc52f0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb90d41744cd94d10bb71aaa0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecd3fe6f580d90498bd2a3c3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbba462df2012747c7af28b0ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc49ad048d9acfb71e84538ace;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h685e17d913d47cd0c57a149fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5db3e93ac90350d41349f9bc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h115b1fb4686ff92bf6dd42d0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h667874aa2f654a0c55bb292f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h608b79882b64b62e53becaf6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9147cb4c17dc1b1f823c2b24a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h482ec2a2589da493e8a94ca35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc372105da351ad85384a47497;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0db632473b1c6fcfd139dd6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h312c83cd6aaad2f623f12e215;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9091980d572082a8179d1d518;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha828fb8a3e5ff9c5b2adf2c68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb38bf3f57bf0b23331971a8d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb01341107c9aa029f3357d447;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee6fef75415b97a6c6f9add76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdb17927528a2c4e2faf743f34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c36e4c53a58fc707805452ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cb1c0dd553a525c654e86ce9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h625b6a24f3c786dddccf05713;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22b121a187c66a4ab150e2750;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ddaa87d4ac5f65281f42b1c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1548450a7fe8205a8dd349517;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b23d47590f6fbef8a83c790f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64a4f8a81fdb73f2d22311623;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadf860b4cd1e0dd99d7d33221;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1664b97a8a4125ccd2b840547;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d963983d1beffa6e1709cae8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9928b143d864c043a7f684b42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa826997dab24ee62936a1613;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e79ef2cf8c2c960436b8bdaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h534c3c3f1c885b3db99405e59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee95e8431c7181ca53441d557;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb83dbc4f00e3e31e05464f765;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ed15551e655bbaa89809c43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9482db7c2656014aca808907;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5fd0619c7f9402f6b6c12dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655aa0585a6a6d24bb6507dbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3711a9f7b3020199bf86a0fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e2b3b5c302512d8ea49c8337;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb0dfc91a214cc32e4221d4f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e9d8b0beb227b1a6948a5c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a5f54283ae3e653560443cb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4636674465f713ebd9c09a5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd83ec7b66477f57bb59fb948c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d5a0340f8fdaab2c4cc810b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaade2c999f6487db89ddcd79;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcc51d67f94e36a6dfe7a6a1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2efc79995b0f8284d00f1fca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6b1a1f3124524acb8caac969;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87532a29bdac90e3a0d23bb5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e414fbe174e50c2ea7a3c978;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe7798bb92c37d5aeaaafac8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac43ad497ad44280f9c19b2c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97fb326d4ed597b980cdd6cb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0939a603c1fe0d608bef84d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f40afdccf488116e0263f128;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89c140fa511a78956008d8d00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77545b103f7ce6b6a1b1b17ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26fcea68233e8cc9b50103e10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d5a248e45e1f6ea4d2fb6eae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbe57ffac38d67dec23d2d3ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d4f646d8db9b85cf900f9515;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebe7c38298808a7ce049f78e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe4618306226ba7d86b6c1390;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda45bd6a756092ef7603e9a09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5de28ad064e420da4a1dcba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89ff861abd9f6a8cea11a532f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h605d4c2d90727d963f00e2333;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h590a474304f4b66c1153cd736;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58742c44cbba21d05d8d7ae2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc857ce1336f44a9f2845b2bb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h251c5150e1f5379c9caba69b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fa49321ed938e4d498ffd7a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c7525a7e2d64592a82cf13be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2021ca5e0e6afad69c7fe1c98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h457f98e88295c64446dc627d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he83a6d8c57df34d7f2b1284d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h993879a49624acecdefe833c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71e786468ad4b8d166662ef9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b77b28b397d031a3a5344b8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15715fdb560ee2fcdc3b0eb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56115391ef3a76d222381505b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h480c0bb31e333c36274b6e8a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf35e3889a8ab9a6ecff026c80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63d5c0f07a1c3fb7508ee5d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf60e40a18705637297e4e2c49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4989d6d724ac82a012b08552e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dbdfa17b46c2af6b6e23c431;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h533506c4fb7a2e72688a9607a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dff5ab3250fabbb275c744e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha23edeeb83a41b9f352a6b8d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6610188a6fcfee384b0e3928f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda13ce5fd160540b5caf85e44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf802e457429fd087d55f9c99a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88b72fb2dc778e05cf0958b53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13e7885152aab73295ec25abc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24812dd534ad80a61470d6141;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb081cb343063372e57466079;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdf7ff68e8d88e7676a6b5820;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28532e0630badab1e328e7260;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e11d9776b86b2df91fce8999;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72643306807819fbcf5cf52bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5407276d504294df4f4546dbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98b421aeef59c9aa3a0fb5e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafa70e8d4429d2c075de15c21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f148ea53013c56085786ff65;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2ac469ec4111972358c9143e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77a8b50c2f1288d15b487d5a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7259524aadbbbd1d67f915af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he93e86b8a099f7523ebadf09c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57e802d54fb3d81784a573694;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc5d6c9ee74f477802b1eb818;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1125c4abd6b7c203ba9f4c4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1884af84bbb422bc3b96ef66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d58046e8cd449b242b6853e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8d98d915f4544653108092e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he568c64cc59ddbde39d1672df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h239e1e46ba686e626ba4faefe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h820c1c44e988185624bb8bf04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd866d003c2e73bb5bb8dd319a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5920c82494027e8e08ccee9e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h729352a750017c8833f0750dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f29646ce3f0320f76a4ab3cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dc46132662bf7e29e636c905;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5bdbce33d9a84c3e03aeb17e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a6f229f3e8a0964cb4abfabb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98105a5ba5baf99755a573c28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h557e02111692a8ff51c772869;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3abbebc866a20407334b58e89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10946832c4b290a4fa38335f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6d7c72092e83faecf43b97aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ea755cf5671316b335b66f11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he365a4130d2d94f839488f201;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h293801978d89d24795cc92e5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6efe16764d00d60f556a7d9b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44b90e3f38d7d14d0fdc7bf8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h687b3e57f9212ee891fb3277b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8691fd21e5c02222fc7b08221;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc49a24b5076b7b66d4a70943;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fbe2897aa8b92cca1e7d203e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a9d18fca6f76122f8f94d1fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c6458ec820873a0372d521d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3001a27af68227ebfaaf7313;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd48574f5536b5f726b1753f84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3899d0062bf7237b174686d95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf661eac5215bf0d760fad83a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3c97c8e82f0a0f430c7e4b01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefd78effb522bba80d6e4d401;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0dfefe6655ffb2e47731fc58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75e2243895ce5cc8934f1eec8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33dc1755f27db14784a9e03c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h468e55091140591c6de4c6f6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e48ad833ef57c5cf67a88c9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49a49bed4984ebfb7671ad586;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ef2de6b19f8afd1c859a0d5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5e87646d5e4ff9b3390dad9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ed6ab6d074f94112b0b15713;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3363716a7d3241eda5d880f7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89940e0c915445b143d53158;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h625da6978ab99cac337aca5e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf939678556a311cdb4976ae74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd13ac289c2b6c6b69080b571b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3761ec4f854e8d1c736d48ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9af566fccb4b382ce4857ba08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd74624bd82a7954cf02f09a87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5fb31cfcccb3b7c26eda4ada;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5f8f2d974c4d46cb16f69bc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb2a649b80c424cae259047c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7d959ea550d4c66313af6de4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21b6c967d81d09847465b5d33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha08faeedf53721fa0d45fa33e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1a7611832b426005713ab215;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2d4e30e0215b28021b9bc7d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde9e6d9acc847b223aae85d78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d1499dbe20e864b41c0d9a48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd34b026113499d82d75d86b50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfadf0fa1b75622a86dec6ccf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6150defbe6994c5f45257958;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14a307f3cea043fb7fa38b3c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c6ae15b7790c7ff6990ead75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc5cdb71bb3f1080efbed7ccf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6de90a86458f0ebf9c9266b6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b541adb75d76ba9bae1f0cf5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa836390686fc5a3d74ece08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fc11e0011b99cbdacd7da6fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ef87ae85fb4b8a6adc64c7a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2be387cb605c12bbf3d17a5e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha11d6be2ab72c9b493fdb1f32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84b7c94c201c1421151bc5b5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h117cff85fbefb473965321792;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f45d7ee967a8b50efa211880;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc853244f6a2f173ba621e0100;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3478dfe977176050b4dbebad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7753fc7edcf53aa0ead9dcd8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h394f4fb1f5a3e548ddd947e6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6fadcd4fb4c9a1e207526625;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e23d7f36bced2960a43a94ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had21981738ff27fe6bc994441;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf055b170017c959c62bf539b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0aa0f65a4f2a84c71502078a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45d5cb246aa57a3314e551a84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dff5308710a06825a36a7558;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ab3770cfed336101486c281a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb294af1eb94016adfe76a20bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc73e108b406e88ab82b8aa5f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h899061b81d930f0dd240fd434;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha54520e30976c0c1e9cf97292;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a7e1cb47c217a139b69346a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc81d081a2b3c9300ec9b0d15c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1851cd6c95a10de7807ba7dfa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13ccb33f228365a3013aea230;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64fe5202d77a2c00789f7ddea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5f1c5896d33fb47cfe2fc8c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b5987d4383d8e131c70c8eb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc26b53470db9825cb82ffefd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bc6dfa8e9a54e611383ba70f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6b33c270f3d0ac05074daa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bc50ef0d47330ec365551c2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h272ee5b9e152eba494d13f84b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2d268c82428bf56156763241;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bccb72e7a1bc9346638bbadf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6db4b19f2b27d3c73f80237c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb515dcced5e7ce2f5b413e71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17f31910ad7bfc69f4845277b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59a71e7cffab1743c32740960;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf18af9f74e39660c087a73f6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9325d6d7ed69dec74ef6525a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc54a1d1234dae3890adc1e8ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h864d6518e8bd3553049a3df6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9813a38f0c09bcd2abf1c7dc0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb25e05904b48b2fd608887ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2873e556a3d0d2959442aae4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b73fa45dd70636f9cd3df0df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24f701fe2b8ffa2597e7c95bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c18408aacb9c1be86ad88a22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcedb8611988e9c55f0b218bd3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13b4c5758e36eed179b26da38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aee46c2598c447142cbcc26e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1192823dbac3916addb83664;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55cb4de58a977055c58dc3fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef74d810509e95bd3ccb14fcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb23efff3dd180c7ddc3128284;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb76d198731e34458155579b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c9977f09bd2edd0f35d61a89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd043aff0a5914d60e72ab31f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h897bac43be4a1d140714bcc52;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4470ba9d9e09ece9a0357997e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58ef8ce1d1a2dfc1499524b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22f746f081c4de278f235b43b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41564f57b62c118d04b51f94;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha28455cbc785bdad4be19ae36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hced4326a9359c1062f0044fd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6af87579e7274765017f1de80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdca71ebe0f53b364bb12225fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893d8476788741d823fbf7f38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h678b13067669622a5c0c7edee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd089852d281fac6e24b5b196;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ee871b730db770393899fbf6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b7f032842fc9294dfd1030ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccd6ec27ece6312ddd3e33b60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb73619f7bf0d4d77ea8af178b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f13f12ca98edb8a700b57e8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ebaa39fb665eeaf1b7455214;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8682eefef907166f50bbbed1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h971111a31913015a303d1da07;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac3296678d4a4bbbca89bcb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4714cb029e60de06ecfa736c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf39dda4b4e33f45d70b855c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h545f1c7ea241f0c045c42c3b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fa8b747986b097f200c4160f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf20efd66f604cf2ca8d47f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1ace46e97f1309608abcb9bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa8645da7d8a0dfa88028c3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ed6c3febb3bc7fb3a8d98337;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ed92f5abc1c156e28bb9061c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd8023ff98732b7c0f6cb259a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8de9c52d481c444f448fd95b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he83723557f26ee6fb015881c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6271588254dfcdc67ea3aed70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff9a82263ea23f6b85dbaf17a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c563d63a95930b0150494cb6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha24091ab2f3e10ee8c66a5e56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha96eba5a0a5c50dee646c9365;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98fde9c864bb81f7451ec7b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6ca3580023639fa029133ca1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1792e3e6327a8d99c4ec66870;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha08b2a3989d131aa453219835;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha19dc2aebc022a327d7af8e9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed56391d1cdc44b6b63c28de6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ed3b74e22472948ed5c41145;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57379672a5742dc9f0486666e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba51af1026b98077f12dfdd6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f9d3fe3127c8a4616ef70e92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d7b21da8c86e53945d674c29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10730b79758e46b756da38072;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfeba4ca7f5ee361e22e1fb5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff8a53d844f48054100d2e070;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cc80006bf6e86443efa31014;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd189f81b31ad534e756aa2e66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h790a4f7eb6d43e9b6107cd688;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3af83ab84c8d835cc03e6d0bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa0183b5510edcbf5a35904e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea753d17f1a5f3a43355895c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd35372cfb384863d402d94439;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c4697ad5994850988bcdec4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc349bd4ef45223d82c45a103;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he24e68218bd34f351608479f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h559db2017fb25b1985aeaee92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc8a6ada6b0d27aaf3c67a27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f6a5d8e4bb88ac906b2f4deb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dafd8cad3a0e14d42d0f5f0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a6e47680893e88928147cbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4824fd68332c85e2a38f9d89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd08b161d11ca12692a2ee715;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h173f76dd423f3aae7b4790d66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3564badb83ab2e4cd122695;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c9e4ebaeab16a9e34fd28146;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b96dcb5997907e451ad8af6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c47da29b54e3ccd20e3ea330;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he662d118786a3e10338f7def0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f95db8c156fc80a64e1504ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc95c3985ddd949f83813db370;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h294f1409e89fb2127b9a8b2c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c607136d8a7e6ca0e22f47cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h471a6f7c62ab61e4635d89044;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h763a9c40394d800ac04f8033;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53a722f532cc29096061ade9b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d79b45d0a66955c87d271a4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3724026a91ddf88837cb2f119;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb662323cfcc0e1e5edd0f7380;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb589372ba5d9b8f21c730084;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c4b6bb23ef3d05737adb08fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h519bb45f3033b7595f326c851;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2ddcb5473e5fa82c24c3bd36;
        #1
        $finish();
    end
endmodule
