module testbench();
    reg [10:0] src0;
    reg [10:0] src1;
    reg [10:0] src2;
    reg [10:0] src3;
    reg [10:0] src4;
    reg [10:0] src5;
    reg [10:0] src6;
    reg [10:0] src7;
    reg [10:0] src8;
    reg [10:0] src9;
    reg [10:0] src10;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [14:0] srcsum;
    wire [14:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h793035f77273b264d3acfbeb1fc0ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f29c9ab656da177577d031d805ebf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbca597e9448b215bfe1195f70661c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd08d9f818d184ebe8bb7862048be89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e51ea52aa29f7cbbee975015bde314;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbfd7b7c3028939084ffa7e198b507;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec57116492dee823444315fac09fd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34deedaf12b5361e8a1c1ae643aba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1afab14218071d3ed0fdd93713cbda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ffa9f682adc2b9f733a083a4c716;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21f7ffabb8c1fb5e8e67afa218b7e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51ee170e3531c9df01819ca3aa320a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha141b9ae30c6cc9fcba01a2a5875e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ed736294a751c93911a58fbdfb529;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80f70b3ee65a586eef10d2df1f7cf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed4c0934147a5c7c3adafdb8ecf9e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf142c1a19ebfd8ec8cc6ccc12859be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a442a07d5a5361c255dfcd6df5a854;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1adf06a9b0a2096fa856f556558155b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c7c2854d8d4ed734132f728cc209b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d5a533829f07b45884cca8f55ad2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a1e438b7ef0915455b653c26b8a4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153704bff9001edf7dc054e7aa6d0ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92e519247e655868326c62bb160a85;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dde90cf90086302acca8cb0fa2c354;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155a46294d1f6e25cddf33dfd825d5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d5f744815a2509f4d148b5d777314;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0372e53d6e72721baa1e3322bd1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h62d01c5edae3347e90b89c3b27e98f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc305e4076b36f976934a8f4bfe1ecd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1e46c3bb392d7cb4fbdb12f276974;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8690f0cbda2732f2cd1d601c761c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ee8c73682cf2529d3c42cd0db8536;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160c993e9c5327e737135831371dbaf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1721963d241a9983552c526172f8fed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b6dbc471d12709ad42b2c4db59006;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb05391af9441663b50b359fb4488ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1489c40bff02c7d08b671dcff495f57;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b87143ad4884ecd5c6b4ab591e821;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192706581acdfddd2ddb9b29e9fa1e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192fd4004d04c6111fea4cb7f5cb06e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ca35325b04e25fb7a1b84bd046d14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he38df28fa2210a0bd70f5b8a049809;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h100f72034a0ae52edac970395028f20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7ab7752c35e8f77b63e893f12781f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he62213e1b04f315dcbc72adfcd730a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d4e09e9b2d697324ae6ff7fcbf35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc03ee8d06e069d004929ae67dced16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12738339cdc4a739b918eb00571dd87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb73d36afc383321b349fb4856711b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4b66c300c1082e02c9febab7d4773;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b1dcaa3586c6c7cc05979eb7a46c4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fc6af74d44f2c4175e267597c9e96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ece8f73a3155688d2eb1555d2aaf8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1539719eeaaf69b92b55063804cd0ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb59b6617f1c76b441bbb39dfc80a29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143360982a2912da9d59f5d83341226;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbbcc7094119c7547c86767a7add36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13553de2b6985c4b677865be6b9984b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb33d3de8eb7383be267de040cd9a77;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4a609807668d5a1f6f8412d54122f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c11f3e1a0b65ebfa1a151d321f6566;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf3edb98e5906d8cae3541d2b1ec8fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h946a2f34da21e08022e0aa9a6689ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8f554b11d8ff0eb79b188a829bacd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b2cd883b776fe5d47f8e3915fa8e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1384cd9dbb066a88617f6e199d4e62d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h29ab23be83ea160b118d07bdc74dad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h360eabc636582fd7b73afa5ef68050;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcbf02e1bc8cd95ff86dd86753fc7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e478076ab140f2adf2fb80de1434c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16db8a53c7c82bebe168a2bce8fc432;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0e2845c062df2a5e51f3e62f48c80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136886e778735ddff5a38509bb0a5fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d22931bd01750d853da760de687787;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19089998074fe7e33bd363b9667fa4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e8914fd5666d774f2fb7310c84b52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152a0c387b72ae771988dea57f7e49c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf6c22408f70abc586763c03c2b935;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0175f2c88d2eef2e12b6d292a8a74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h408fc950d50e75343e38e0ef8034a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191ba4acb180e5858bc9fba1cb2af0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hccce4429deaa7fe3c7344bfd3b11f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18acc11809610b71f5f5ab0493b3c9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe283cdba9cdcaa4b9f34f90889a8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13aaab271ec4ce25a84e91d3d2bd4d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea2822967b373ecf8faa554838967;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac15d238ace2a64dc11b827b5379c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5e5426c5719d7065fc5074a6011be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h666412da1b46659141661cd6a13769;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112a7e0b48c7bb41a9baf31f55ace69;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102d16d6f3fd448a58c1071bbb09b83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14aab484c82a2cfd4efc3c6137934ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ccb9db8334ce312b9982208bd34679;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he558b9691906c539c0f55d8c18d324;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1860e1752c7d73b5a7fa7a1d5365ff3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19362c1d6810df062552824fa2c0914;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a33c415de62c7d15e6a0825d61013;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68fc2ab370c41a16175a8e5fd690ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dfd50bb2b154b4dd3798cf9838883c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18682e764fea12608cda237807dc61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ecf50154281471bb630044846e7468;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee753609400dc1055a4b4328f4c677;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h274404bcf7477d70124dcf23fc86ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149f90ad05a5dee53a5cac45329747b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8515c72d1a7823fc6621da70e3c5f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b641598e263ee99f52b45e0c3c5c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he770c625a6f7f295ed0fe6c6f73074;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8bafdafbcaed21329887e662b5987;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadb0029d2b03b56963a3685805d7da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa53e64b230f63be601d325f8c82b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1591f7bd792bece10b6d91dbe92706f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d820c413c2638d00634a023b4dac8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd89c181cb74cc380694b2c70d711d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c3945f8a0bff8974dd6cbe4a67966;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123fba83343fe0f8c89789252ec9037;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcb64d8e03ecae39bb5c0d3c266fc8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee2ef8fb12c1fda3243f9186673771;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ea1462bee592a36c25254c840aa35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d5e37d69669f18a029738e342f823e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32c5f25e835a2f7d109b2b70b14bd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14087db8d52fb8b8fb8784457f02716;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0f0f0ce09888b07eb5c7b8d566913;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16768ac5edad5fe5fb3fb950cb5bd62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112587b4f2dd54e19f262924cab480e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182400d1ebaf368a211b3e9c66fd79a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd2ded624097eb296e75cb4f452276;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b65fcc6c89c3ec4f0587e0adb41b55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1813c9c72c92b2bc4029251a6ae7890;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1e147da55230d7d622effad2051c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha172d111a71b66f0d9ab71893f25e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc7f32970c16f20154be7c5394d2a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48648dd06e80f7064e00ff44789555;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he586767b03ac101ad62e4845d73970;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4e780287327db8a20602f9094c239;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95db030ca60f788469178a85eb3a13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h342b4eb74a3bd60e6704ab565ee809;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2acb72fe1edd15190ad5004f155b06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e1bb753f27e419e4ebc8dbc6774b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ff07dab83215187260b032f7a8f3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3ce0fbec80f732f91b10a5925356c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8e1708b531ee5f630a139b9645d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142d7de4831e866e62408d9d1cf1670;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b24f07ebad078b0b9ddd699f0b452a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1794f574cee8a972e5824368dbbb86a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec2b7f96c6903190b437e45b35d420;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c04ea7f1ffe5bf6e39ed0ae20de9b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb171f21d0318c4503ae69c774d5fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6ddbddf9e2adf8cf92a9dda370bb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f071f593430bf75f395bab270033c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a6d1d961a662498d90335713869f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h285e7657f09c883312a17f6d9956fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d2866c180ad4224dafc46e02c6a8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bde93e4bff77c5005b0552a1e6cb0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1edcd618b3095d80f065f539ae86a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a298bd066563601d803814bf14007;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a691b8f56189feaa6f6d61527a8d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4d7877e849561cbae6808a5827210;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c460185706420897aaa04739fc1d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa67150fbde1b9c5316c230abc7c44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1117f6cca0d29dd1d4a38c725d323bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c48a35f432be904c5f1867edfa6eff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8136a5817c20c886185eafc88340;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11279679e96adf2f20c63a444d3520d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h70daae201a30aff60837cb70b514e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3c11ac72df656b83ebbb502956678d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ee8eefbe7f8d8e70c8ecac13abb22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16433aafc2605728e0a0fa74f2963ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5754ade5e1e735e570500172a51d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cc2daa7e8f4fa0bd335691054537c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11712d054c03cc7d61011386502f88e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b158cf7edd5441aef3b850166ff3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a931bf6576413b03035520f82f7875;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83386342f4e84a391c5a6d0344d6e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49d8522200f14ed7984349e3705e78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h721d11a166bf262c6a17f01c501ed6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h874c9aa6780857a7666950dd74a7d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2af4f63fd35305a3458e6e2042a1c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcd98b0b51563e1b6e9e402a2d165c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23be45a7b23b03fc3a7825d5e9fa2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117c750f913590dc39242a21fa80ade;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59776cede75a72989786bf3373c988;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b4d7b31d093cece8e5b2881bc1e72;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1620b73d20716f02a3418c085f356c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13db0b84aee7fce847b0d75d1d98cbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d7b1eb2eabd53b915c622152c031fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea5869fe941eee02897b6103f90c97;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h477c67c697dabdd48c7da3155845f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he9025d9ab746106ea90d8d388e1af2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h132184866451ec695ca8d3317e071fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a12efb187291f9ff79e751d819b89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b600200affbe9001bfb824b5fa8a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5856555cfe13a91ea54ba6c8faf5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac230ce7909c05f11639ca175ff461;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1696735bc0b9fe4d00be17f314c8a8f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117cd88105dff1e299e5e82fdbfbc05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef64d97b4d58812b459dd85aa4a592;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c581e6d3cf191c222b189bf572d838;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e31fa738604deb2579de27a55bb08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1231e83e5c9a360ee1b18be7b810fb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a23096eeded2e467d7d1ceb2bb037d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h232190682b0067d421489d83beb7b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b0a188b10dd220649ee541eec1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d051b66cc6fb6979c1800db362223;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145c2325c8c6bd02946965c1521ab41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f4334a19af753e640835928388e21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac13a3e715a95ecdc954ae43746e65;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eae380245122949513d5c3a0197ae1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf152c80c55e9d344bd9be98579c4d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191e641bc16aa9005282685f8c1e73f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11fb6188c5cc75a8a4477cdc7ba0428;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h150bbf0e21df12a0095a75dbc40c94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df8633eb80d679ec348cb7e761ee5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h62e447a7d8285c0714bb6b5fb752b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c57677897dbaa2cb42ae568cc3b2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156c5a76f8903940d9ba2ad0ba320f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96cfdb654161323d0fc3756a29b2a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c771643ba46364ed35d06f5ce3310a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b4f7cf876da62db6d2ee3291094e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1abe5e19bb07f3b551dc67e5c4856ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26be6237ad54b358acb12f10a48d6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c247b27c138de07c131d99824cf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167e8373eb69c976fc43e90416b2cf4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0d06a1da9a44748779d6eea1e73ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7446418d2585b0663d973fd971a565;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb52968453760d4d5d7e65675aabf67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44608c64cedcbb2c7017d8ba21baf7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd69b76918182553ca620c2228733b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7879d6f3ca2f8455a50ca5a75e4b75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4955639133b994f5a112aef38f228a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120e5a6c85ab9cc41be4a85226729f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b51b4b82eab73dbec6d4cf6fb9e081;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8df4695fb4fff9b240c0d8bad9fc03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53aae0890f9bc0161ae456f482ccd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7f9a49e8f33c0ba6ea3fc0d8772c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1372a7fcfaeca65f29e6d40a4662390;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c69411ceb97010a1a2b817863052be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d9c3ac6bf21ffbb6797fc28f02afa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14457d5a31e46cb85e7a935ddd7d9db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc38b902bb0169a543873abb9af8513;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h204195995b5fcdb44ab0d2d28f24b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc072341ff137899924cc0d8ee83da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heecb0c64eddb9dec1a092789ea18d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8897ca583f086a00804e174fa6548;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba0e35993a01bcb9239b2ce3f15f67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3982c70a6e211df1284f6982604b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14fa19f0e3ee4f128db5b0f2353dc09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1748c45ab2839d42990084c294bcbc9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c44c21354c604bcb3d2b5409a36c0d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129ad23abe0cdf3c64293baec355640;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab47c3dca873a9170ca5042c1c7f1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0149a333888520f806bcfe50173eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14733c80b42be55f1239a32af09aafe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1ef2f434ad5762fab8b281d305bb1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac9465b11445260d7a179f05458437;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2e9f3bcf2009a5c26471f7195ad0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf72e9cec1666e517ba52b09e53badf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c2fb0ed618203f5f0b9aad04e3b0e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f129e0ed43d65ee16934d69a56df2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda0820ff40b41f9b4c14a6ca85a363;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc366cbfde53c77e74cd9888b2be2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f0fe61435073cf347529f373fb0ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h616b26a26ed8a36d1919880d76a699;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha79735acee1622640c4f0b5a845f74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be438ac42a57c368e5bd9da4145b53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4d17b7791ad802cc14f773af0b15c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e8c082d672989abeeb14be9dbaa62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1269def5623f506441090176e1b453b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc025d3d878dd0354bcf9b0930d20d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc880673ad58fbef898a39235ea1c62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa4d6c58a1a308cf3cfc002393e3f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h491022239a269f016077d2f2b336e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e76fdec241dcd495a0897d900e442e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164c648aae52ab12df424f087c0bc3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124afe8686b94233d56f15444e1a3d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b9c098cf98e96b375c14b617ea55b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7760928212649dc6edfb39b02ddd8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hafe6d213a50c963a8fab6afe96ee47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41484e5e35c6f08db85e71ad4e5387;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a2df06191262670b347bff2ee0da1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b0de04fe1cace3e410c56b54c1fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5c69b9b470a8c0bd70ae61f5dd1d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15349f0b12cf771aefa396a1349a1ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f805085d693fc702245faa803dfcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac8308ed64398f6927b8847081d0d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd26421dd98982262190d252258447;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e6090551daaf9ec55fa80b2aad8664;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff56f5ffd438f88201ddd8ef5a43d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1351640bd95b75412ce88f6eab14afe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f71fb633382a3689bde82ee9200d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd69efcd1929ecddbfe3187fb1f43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1074751811d501dad51e90cf3665175;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1adde809412d5ecf74f6575c877144b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h428684886f91aeaaa9fcfa07b757db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9127be01148710f96ab91abb9363f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cbd20a9e605698f6ebcd7ac558686;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc30c97aa679e9603d174347502b70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h229e6c202b13405ea4def0113ea995;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157a7235e3008a3db4c5755b9d0d9e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78a3924439b44cbf1f6979de2b2538;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83263a1629aeb61cf643b4755fa5f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcac73c15a650299ae5bc8b4dbde4c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1653a26f73c2bb6001af481f0f1bd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6d8d7b16ec258a2c75470ef0dc42f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1074da5cfdd63a91292e3eca91c2f94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167a19262d84d248badfcf3c528be3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e27bd93a04a91aef278a4e0341305;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17706de518e0bfd9931c61ff0b5dcc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28609d06b9427a926ff4a4ce0a4f49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120c49269330a04c304cb00e534b11e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4184e9f6a3fac346920654c2b099b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d22bef4d2f117e0a53fd57d5d90ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171ebcb4688a0683abe4bd4a6f59859;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1116bd46f87df4fca2c7d71edfe4a96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b241f97980f4d9bdce708e02cff41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4771b620d9a74ef92902d5b33b48c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f46c5a07fcebf08f85cc6eb1999e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1e9fa576ab099ecc2b81888155f52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bc74287c7f2e0f9011258be8a7d46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1215b13066747e8c810c0a000ceaf38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ea6a4598b258fd916e2cf121d9c84;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1b028edc0cc2cb94ea152fa969c6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbed279797d862a14ec4fe30b7fd9cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbdaa2eb8951f0ea444755171b57c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e81435c34f0f1cb5d2c4b2a6f9116;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bda411340d042d91cf19720fb0154;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1269982df9b20649c0c262c7e874471;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b633833ae34714f4c090760099cdd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba098960f60aba16fa52fb0964c214;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1529d56311dda973980ea1b23dc0ad3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9398fc94d99476e36f497cbf4ab65;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33d090f7edff426ab1a2d59ea8efff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9ba7a4e2c7010735319812358f415;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d85dcfff6fd46e0fed4ab7a9625ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfd1a6161e00bc057c678d55fcad7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1f0c6e82cc283dd7523e2bde86629;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa49234226bd07954c6115898c57cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44d477207788461bd86f19046719a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6e0616e2b6c478711d7effad9fdc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b79e9748cef590891081b3fe59dee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbaf8f1f268de65466d1a22818ae44b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86aa542cdf341f63a47b4f02b32c54;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac2e66605f0c8027259b2721d5f7dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha38b29ee7e0e2751999e8d1ff813c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10908653831d14d9afb0599d166cc67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d6d5f744dba21b6e5e4cd7d53d931;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10accfdb5b76d2a9f1689b873c39f7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b91292eca0f79dd1feedebdeb7ce3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c06d2e3f179de064781f4eaf120f1b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c431fc1f5b0ba590ce5893d045e7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161de2dbb1b8561ae873e1ddef14769;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab268d2ce71fe1d5d7432461ad66a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac951b0e858c66fe814ddd0662a2f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39e38586b8e3610c8fa7e99c3b0738;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a381f2874c3e73bbe9b79fb156a835;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106882fb8f4014cea67ff52e5a391dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba6d235835ce1dbc633e8c1e95054a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59e4793f59853196c8e70035b24fa2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf04b4a993cd680e6705f69f06517df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h821982ed3b236dce43fb9cb1a50861;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h498d354ea66dbeae9c2900ab2e8359;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1523523139b618fe3a5208e970741af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1479d0f19a6946b54d1dd3cd9bcce17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27a6f2d80148fd71dd9d84b42f3417;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1519b4fdda11864467245a854353481;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1401853c0f0eb453cdcb87f450d84a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a6549b16a792ff4eab63cf16e5c38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6a60c5fd31aabdb60965d024adae3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc167cb24aebb618b55759348569aea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cfb299ef6da426c8691e05b91e5d09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89d186516aaf98c3ceb6bf076e26e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h545c2690f12a6d42d3bd6f065ba8b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfccd41b8be8702212f0f49ed78b58f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3f0b6c8faa6fbdf3af3ff863ab063;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd36f56d53e603f8051ef48f5bceb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb5832cad7e44c29261c484fb67f52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82fe610ceb4f1bf275765d56d1124f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8319c59650ebf9ffee5e56e44eff1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc04237722b4f8ffdcdfcfb2c1de84d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a626e00c3eb4889d08b9665251d715;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1637655554486e6fae4b49ae372014;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3db913d47619c2baef295d7be8b951;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd76cd7fc5a91d3026cf4002944bac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3bdd9707bc2ba0157666bb97533a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58f87957062f2ac2fdfe31f17bf1d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd47517834af2ef9414d0d4b06e0ad6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7e25022499a247c0c52e3476e39a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9b8e2fc1992cc175ec6bbc15d5142;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab2cfa04bb3c6ba8a8baeba3d7a4d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h623e59aab1749d1fadf393b4f7ad86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3daa421e3e2cf7be8aa131c9fe95b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13dab934be8afe070b63911a16fb2fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b1f17c0778082b0ccb84ad8b0afe3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h993f9243b982b6e665b0c712cb3968;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d2ac4e7cd51f54604ea31ec8facd0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef4fcaefc549a965370be210257161;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c835215f7655ecf6076f7e5bb9e3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb126d8f45cde7af37710a91fa4b1f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c99c95a17f1f97e6ccffc168072f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4979d6715fc544216802cda61188e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71134567e4ba4d3c150047175ef30a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d32583e006e4dac5b4c9366cc6882e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ecd1bebfbccc414c4514c2785fb3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1774ec0567fcff4010c8c019b9dcdbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a163c72f2b9bc1ecda0675245a62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab1c12c28827ba3484107507fa077d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bd84db4eb0c5b6bf2cfc7e1485d00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f73cfb13df50209f878b7128542e58;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d20438aedd218ddaff8c3ae9cb41a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd2b789ba4356a9566c385b94cd2b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a6e3aba5c3e384ca4345c24dc98bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he83e0c3adcb367352ae6890b40ce22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9f0e4d9da69c609946819d0ce827b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e21643ef6f9fc5b3ca5362cc0803aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e77b927ffdea4dd94578f9a87f0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed3faf31b121c40a0640f494f3bd58;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7e06ad6e8d4b1145ef4d7e12dd72;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6f537eb19e91cda269006c36e055b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a974d9b234baba5fb7bba8f57fd2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1543c0fbed644b52afdef5239964ec5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129a1f48851521f26ba4c0bc086b7c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h327cb8d0d0a84e08063f229fcc1e00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86516f5643770b42bdf77785ea21f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h93189c02deeaa7384610cbc815c149;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2082ff311dc0db08d645910b52a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ca8231b2d362fa10ad91c46c6dcae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f17906a5eaea73b8bb7de11283f6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7766e87d81363f4ac41bf8843d356;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb987ff18df3d80185b98e3ecb996f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b95939051314d618c0a9f175533447;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbb3f91b0a55879cd9d26570b5cf28;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd2ef0476933c52da19bc0f708550;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c3deff70f4e986667419e5a1a2d7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e6956d03a813e5df1cb6e07e486e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4aec1886c84788dba3992d51ff278;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c96d4a388cb339eb2d773dac084d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf2d1b0d48e4864e3f1c6b142366c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170487ec68f52ea495da0a6dc02b080;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134f336c6fb23f2793b817ccb153b7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he803923484a532cbf860d29dc67c62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f83c4acd379ae7c2162f99eec7750c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192feca8035048ef36dc43aab43b2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13606eabb686b12816b8db5be014634;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb4d1fa4fa0b267ac346d0d6ae8c08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188f319049c126f2d5a704c143c0784;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb568c90456343d94b8d08574ec0893;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h753e9dedaef68906d1ec9dd1cc3eb4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7704eeb5928cf37e4dc64e9c060c06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151bf7c6da68a9e5accf646220a1ee1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f43e70539f524d86f9d885b96d633;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7e2b90e9cdf222ef9fa998a6d18e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d34fa56ab9077612cd39c949296fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h150d9f0cddcd8c537d11575d91ede0d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1461c2e1b912df57d59cb5bfff3ec79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0da8ba6270aeee4bf4e87e7d463a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9333886fc5b5102f9e7d43ccee2c03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc4cd5666d0d8b80c5abe137454c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1803cca2cb95f464762285248e8b39b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f825a3b0576a97dd5f694f2057c55b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13af4da22ea2a5fed7ff769e760a349;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3e1bacb109f296f708ff3292f8c3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0285213a2dbb4ea8a2a1c0e47f7f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5f9317e7e7f1ac35444b933462678;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc52210fe7589cef0ef1ab5f977e1e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14dfc9052b8f469b020e6b53575f6a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a5ec0552c86cd30ff247b2f9f6727;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5126e5c7f9b65161d19cd55748346;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33017dc2e09e9938849b4fe27d9223;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad19774f9fcdc8f7f810a2f0638a3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a10b61ae7e06ae96843fe6a762a5b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h467647bee6f0e68637d5812de6064c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eca81826c09b63fcf34024afe35719;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdab35cdf9d0e68fc9c6690bdd6b471;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ae0d3cf91862e990ec9563df782af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc48559f36faad763496778a129def;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e4c6b6bf6fdf916c67f005ee12c72;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9bf1104fd4c11cb36c0919c5a49ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b88938f2d95c243fdb41f08837390;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he28f4efc7cf4a5d39829eae5d5b9f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1d8be030a709dc596128214655a2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6101d09937383bb99a33fd0e01263;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0e4deda3c70f43027eee976e16426;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd261e4eae6a14c16eaa346336b7d62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4dce6403b2d314b438fcd2e53f9963;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176603ca43e274ac135a54ce18085e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc485481d8915d75534e8c5eae53d79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107c33f328a019e7a10130cbdfcfc0a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6f3913101f688032a63867796e076b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h451ec4b70a8e322ccf2343de855968;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b2c29a2ab215b24431b3e3fe02d176;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b5529c15b9b314d1cdf7aea57be37;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103a28b46e85add824d16769fe99913;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b1d161b522394a8ec49fe1f8e0e59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4fb2a69e650c205dbe1514557998e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ef1bde7c702cae59b66e7d0fb45fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135320fd7e1fe460c2d9fdae931ed47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b249bb82d2823b2aa164146e14ad64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7435272ecb6f04fd3d64b80eaaf2fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f67b31bf61cd2adc9b6b84f2a7dbd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1349472c3a80ed784d995d81c132f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1285e341cef2f92399fe910b5dfb433;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4940e000a061911574b8f98df9fa21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ebacb820ab90166420e0a2cf0bdd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3987172bd4167b0d24cd75309e3639;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199beea14531d19b9bc08602420dc6b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2079ace2560263c719eb97639ca9f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11277cbe38029beb274a83a03494c6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee3eb9d0eb85bd6f59a52d2aef7b7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f17e12945f051895019b20970ae1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134253fd701309120c7763f2ff67d5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11158b40031906916d678cedd4dd213;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h469f1076dea5aae12834c687af36b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h185679918c8b67b6da2c2039b5c61e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128378c8d57b6cd32820e3ff89d1f10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a62a4f3e841e2ec8cf4b774b56df23;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8fc97c56e4188f87aa8667e472088;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167c8cef7ad9fcc210bdb1899faf606;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc97b2906800bc0d9da2fe7a52534b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7527927882f1a627bd2ae5c2d3a2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184cafbb31887ed6e4b043796dc9200;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187074875e61f0b6c94f643513735db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1205332cfd5c056f4d1bff8c906b920;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4f4180f8111f5a3c7d172e9627952;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bbc417a57108033b38ea0c0ec3255;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h154586b473e04c72ca619ea7e3e5067;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7100e7585c07eb463e4e9af10b3920;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a70baa6593f9e30205298a8cdc2eef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12920cc57632df73c1bfc1edb6b884f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce54d8c85fe6923b7ad41e395ac268;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd89e7c361ff85ab134f3857efb4581;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c613cf98e8bf39f0884d398ae39a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbdf8d493dbea0891da52b0464c9e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f19a5dbb4b728bf87296b20584d6e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163a38673c482a47aae9934aa3fe452;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd15d0c976f34461cea6b700b00dc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f399cf95e01b506879e4a7e85b4e27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c424024f1e1e8cef26670747d559b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125eec61411caf1f846f0c9b55ca2f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120a1c47eac07a1f1a3cc729ebf12ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7092eb6ca2425ea9e1626fb74e059b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167755a6838a5a8be1fc61271591ea2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9387042cd9fbc18132a97e405cb8aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae5c930a90af036d0ef255041b93c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10600091aca172f173ae9b88e1831bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a9967c5ecfeb97c7bb207c8cd77d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h438629d92dbddcdfbfebad635c4361;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1795021b6baf09665c7a1927315280b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4e8e234286cbbdb8385589f4f95e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h542d907893e5fd3baa46a064d2ec5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181dbaedac35ced39594e5d78faaea7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0131e7c07fe9d9fc3ea2465dff405;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156432fbfd28fba8241ed3d7f5d4065;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f88a5a6dcd9742b4b99df65e6ebd12;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4d1240005750c860a25c27b886b44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h457a86373d3a2c268594497a41f7df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8951539eaac42354ad5e77797df503;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc098d9a9f595255048730689d0d5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f3bbee40706f3a127254a7108a50e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he40085ee424fe273ceb229b4b50841;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he210b529b3b119122710672e6193b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f9ef3a27615aaac38a5e13646e470;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153ec58b7d7dc2a5487fc3d6afd4db2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1852e12588430d784b6adeb285b1849;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d8cc725009fb48933a02b76c917e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18dc31445ed119c309fc13240a14c48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5b0ef432ce8446e81cdbcf5ae2df2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b548142345b968bff9a923fc99a9f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1edddd8c0cec77124b9b7161fda8aa2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c2764a9c06fea54c92e8e5cdca18e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f63da86ec9a3388e9e4444c87c99dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he202c390718840799f5ecdddea89a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c025ba2fcf048bbf535c1bd04169;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b2bf9d21560e26ad7bb444f17dbd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haabf68de41efa9c25268bf21ab1098;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bdbb96b3d92237b314cc7c12304be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56c96f05c65e0fc6a844fb6e957975;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f69ee52033dea3ed53f8985139bc7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176f6f03b449bccc6827405366b84eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f76bef2e6cac81c022241cd83ae31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc14fd826b3a57cb65a1203aa37c252;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184b1761596d008bc559f53f7096ea3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153cc11cc3c3132ad889045325f79a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c868e63ae69acb8c9d4284b2209f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b864206ab8fff1b30e6641c829bfd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7088d037cc4afa8163e5355c7e05e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1c7874c917f2fff625fb58badb049;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa6553105d63c5107400cec5652d07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1526d2d08f6682bebd3128f38d19ec9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1adba6898943933c6efd33701bc37cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d9a18b6f3b5ccfb95619e58262b5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181cf79c79d46f9f2cf15ee572a25ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d9abb2cde1325db2174cab08ca746;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160c3d3a1fed337ad270780105870ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75ce8bc5f5f1afcd331da130cab2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12868f3db72aae608c7a726d5d67f8f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1966cf3aef29f9e9d974cc0bfd556f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190c5790226b3887ea912dd563a42ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd04e4feb59e92bdf37b2129a1087f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1289d127762471adb1808c54cde0424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175e2742c69970b1fa0f6c9e4e2886a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65dd09d54374d0d876a59d18f1a5f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb42d91732e094742335ebfe390761;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c604bd266d9f379eabb30eeaef894;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33ab8e8259e866002618998ce8f19f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c28ae3d1de5b17695a982d65ed0e0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e491edd38daf6078e3579f76fba6ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f66424d04552f9481f2a221e67590;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h281d301d1ae058fe48b5223a3204db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a66d64d68c5271bf674a0d461711ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51a16ffa9e67570c142a0379388e2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6cabe63df44df57a7c03b9dba45b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab9609fb3a576b1fb3dd516db6edb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8abb7e536f2a1a89cd19ae7db4130;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1891568bfc1b28fe800b0ff278c3696;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae0eb2f430aad534e49185f176d80d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50cac431285a56573619fcc3f12918;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h897b9148231e6a348e50e52dae13fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b1db5c2d016756adfcc7d0cb5e0e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7c29993e9cf4d60de915debda6a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18652e1b5ed640aa397beb6fe517107;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135b280f841470eae80254bbb59bf26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14fc08204039f59ceee27e685f0492f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197d272da23514212057863084ed2c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1877aa2224fda3e10045a8208a23c66;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb9d216551c86dc40f7fe1a7b9949f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1633eacaf0b9e5250655298e24e3a64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11214c962acb9759d7b3d1b11e97cda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbd4acb814752a322eaf8ba877e219;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181885b372e87b9f430a498fb7811e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ee2422afbabe40ff295b5893c0d86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1785bb2e4edb2e473ffc8235dfd1a7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8b3eaf20f5b08386aeb9ae00432b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71b977953160a13a15eece3a5e5276;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f7779c94d779c91ff99419b14826f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a81cd8038d20963e7d6a23ff74827;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b5e993579e228d8ef5e487e4de090;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h337a1e4aa768ac55307e4f5418507;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22648b3b53f69fa5ba4b39f8e7c0f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f608a5b2df0b529f8acea9711009b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3925c72456806ae9b3a65f0d8824c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1410b5f6b2da3e2cd3ab974671a7d1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9ed811a7450da4673633399beb1ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he50b23103e26e9192346d09c66f915;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb1a060ed78b787f51d50f0dc2b874;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81c68b30d28233b0bf7930d5d62d6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce8853afcee498affaa1a1a127e386;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ca38e75918b3676d13bd91036b9b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1128ef162fd71dea123a7a1aa2711ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce09a3e3265a1e82324afe5d559db5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1336f2e860d911df1d102debb2b8888;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102d6c9843ef44213928fa8519ad1a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1196dff3d51e20df2aea617424a30fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131fc4d04528a44d40dfd463ff70148;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0c392bda8f03ed250e40673feb8f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a392f390d9811eb0e9b1aa05f2be96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60caaf8b006f821234ee03cf9709c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192fac26edaffa510499d94fb98fbcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131e890b23ccb87535d0144cc8e2626;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha131b541ff45cb54f03592ea39f1f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7647d3c463121efa8176b355f0ba0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2eef55711640a6c3e145bc0e5fc31d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad1ec6f8d71dd0a4d0dfe75986ed55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cce8c5a358cb06dd7ff5ab154afdb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h656385d3d51f8ac0ef12046563047e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7bf8b15e5df057c28353f33a325e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19842ed249544e98a16f76a1c14363f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he06f75c70eb0ad2ad2c0499fbba78e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d1463d3798eafecbe15a06acfad0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1669fb945c4ac7773ed85a9f21a728e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5882e97e67757a33c9de7ba5b604e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1518d0904a5d562389fdbd096773108;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14702fdaee21a6072d06fd97cb77b62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a64efdbed4f51a7f0db082952ff1e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d93bdf800aec0d71f7c09331c376;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8a11f766a25e8ad8dbf952150c0a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6a4bf2e7200c73f8d4c602cdc3db5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106170a9413a252b4ede46bf43b2c07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h895d60de658f62eb55642f560f0c2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h116b36d0fd0aa7a98df80beb5b5dd7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1a4c055466f5da255577cdf3ae2b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12af40f70c0bfdc70064f12526d8458;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d280dcb985fb25fcfac9b12f59bc7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ab93fde391dd18574eaa8a5caea36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1034b1e5c578b8ea33a4d611938c6d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64105c66f31aeb8a9b87c325871648;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9cc56de1b6b1901361576ba8da1b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168c9dc2967a846edcf7efcd2acaadd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ca4b635518e8526bd259884ad6eb7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a57bbe0aa65d9bf3d34b0100abb4ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e09f75d89ed2a50a455a8025cf0a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bdd9b5032acb540289758a3b4bdcab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4af4feee1c577cf782ce406c787090;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1deb150f1adbaf73f1e23373616268e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f1e3bbde3b2da76b2907d0376336c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191ac5e401befe0f9a98b6329bf257e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1047ecf16564d84121b5c65cab25650;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1726350f552bf310f5bcace675f07f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hefbbb66155a9491fa6692bfc158506;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e7d99860ce247987c913c2cbb52a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8941ef6d9770952d15c1e860bd732;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb692868e675caebdae80987c3aa57;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142df65619ea08b4edf7954a6f59d93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h503a71525efa1ef52cc3b6808a42a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac0478c5abaa69ae10b86880743868;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188e7f14362b54d2ceb1ac21196f2ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h688a706d4ff9c01f858e82e249e9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha060e08ec6adc715c02d5318988dc2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175541198fea3c40481abfe0ab72508;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad4496122c01010032378c0894b33c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcd73691c3b99b80dab8e459efcd06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1824988bfdd0b9d725828a4ef64f6fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ae14bd29cacbff52092e21b6c447c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186ca0271b880cb026db49644aa69f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ae0bcf487dfd957bb1bb5223f221c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135f6df910d53fb75bd80ee38fcce42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c5325353d27ec9cec1c681bdf6f2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14479807980f47e2feea8dfa069a0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9b781f4749fa698dbe4ff5241262c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1939c421cd62b60f9a8c4b6083609cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc245d871a508b428b571d25d21eefb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b4fa26560fbdabf72800ca1344b7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1415cddd8aa80161f424c0b6fcce64b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10cc2896e87e7928c51d07357f8e89c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc50a2a5199029dd3325389a6a6e93c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb1bd362283b0c2d02adb05bcd5c4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1313e9f686a7343933a0a78aca253d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110260402bce248f50630dd113dfd20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ae567a726c0eb00c9c362c1dc6e4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5a64be9491af5e3239bc15becb9cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1951a27e2673a7aee57c2f1ff77927e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb51267990606e259884425edc2455;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f3476b7d7a86801fb82cee36caa83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34ca9a2814e73bd06992f8446b725d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb394c4b409d0d8aef7aba88ce7525;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14786461013a340bbada47042390f1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he15827113db057bf7018aee439ce75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a34a2a7ddf8fba56f49521b2158d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1896bc7878fbdd03012c6f7ec925bf7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1760eb3b47404d716a5da672d19b9c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heea2f3227ccba92c6f273d5c08152e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd333ee70bfee557d5591d4a443276f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2236770b8658445cf55c954632a6f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h909131807f33a11981ed813f7edf76;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6727f682a7bce449f13fb07834314b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69ca1863604c1bea5c3bd301b9cbd7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he5812a865a91a0c0bc93af0d7d8324;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5b71ae45be6647a733d650c3a4ee9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1afa3d7ad6a9d423fd284f3dcb86646;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1801c932cb0e3333b9c7ead3509d15d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8951834bc1906720025a35318cb31f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9201e399e7fa55d990b7e8339317dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d8adc79a540964474ed973955df80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a4c9fb5c6747b84c562b9e57ceb83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e33d11913e8324d9bc436b2ab07d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h621e12f3019e0b7528251f0043ec9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f868ebbaae5d616ee2bb96ceee82dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbfdd5f0947f8e9b9e5f83f03612129;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a83c69f50de5805df59a421afb9ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a850d4f90dad609d200eb9d27b505d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc2503eb9064cb6ea088750fe60331;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106bf720cf8602b755dade6561c2209;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba08935e2625d326107a7cf49a64a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7ba5cf3f784e1ab67c290604af2f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199b01c44901882b0ff1e600f09a88c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha99210b52ba4949614aa2cd8b88b2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8183f1c75f07514773e3ad37769a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hebb32c5277b8ad710a6067368f47d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6b7f9fe7006ac4185361ff3ac0a0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72fbe2e89921f3f3a30203f89908d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89c11564193645b7890b8399a8826a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48e3390e7435486fd71f480b6114a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c0a840ab61aac827074f6fdca6304;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2f440660d85f9cf669be0140d0343;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2c5ee50fe0efe0c58120bceeb0b07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d82d0da05da23d081f3208138d0dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a60bf433f636d83619f535539c698;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b3536882ed72f08f84735e6bcdd5c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7afddcba58f0bc9cbaf5b2826182a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haef0ff430ac90f67285c9e26368da3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66ab3e11290de32f1247a788c0c565;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h280a328bb6375537b08370aec93532;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a0c652eac4131c4fa49b94b2658de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0d7015af85729d4f7b00945013110;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f43d6cf104df10043430b8d9c99a87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118a4dfad1114fc36c39be40d3be9fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba1d157fe7cb3915f818cfc5bae66b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b24b9391c7b9e144ddd3fcf278864;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35a70b3d281e0339233865eb3471da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac822f354214e8e7e86bc78dd9e563;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h543fe7447e588f4c1e1c5e9a5a5258;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d1021778a8e291dcc07cf20725742;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5fcd68a66d2126942f8fca6a072925;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cabb7c39a471501e59043d312a6b22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ff67b8c9221aa44329dd910e15a2c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b2dfc23a2f1afc2d7a26ea26361f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb8139372e35e7949234e6ea203090;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1536e530aef0032a1d43cee52dea44b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12fdd836c656f442f38a0a5dc82ea18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd3b6e55172219e8c139d054a0982e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186c3ae700ac36557cf55803b5d190c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e5ea15f232217dd4da27899ebdf21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb0325cb6e335d40cf6dc3659a7800;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15cbcfb33e94de7d83b1e072261926a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde663f0ff2010267556b2dc4359916;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1684990cac660499c28f06786879d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d912c8a34596720414a8f47582bdb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4b9730ebb64d3a4f2676f1bc6ac82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16249af47eb4afa2e296d063ceda56c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1341f6aebe507ebeefd95232aca2ba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd080ca2fb92c566b23aaf950d55e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6c702ca13d21e160c0269da707efd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dcbf066d5c09a988eef2e8eccf592e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1869fa71db8943f1f0d5692147e8b4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a79430fadcb404079313d81224cdf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e320b3659225c574a5d736c0af74a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17935c441401d80936c722c83fc03c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148e6c4142eca5c60c90ae4c09a9f57;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7c5874b63e867556723095fb4472b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2900e4093b39e0b194ca4503f1834e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24a8fb388a773287a75faf3de38ba7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82aaa03dcc3ec59ff5c579af03bd4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1915ae0fb594fe3d0c0b2400cd89eb1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19491d9e308a4b3839f2b32f5881c0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c2d2ee70124d2ba34b986232b7106;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173493a64fdd83fae5ad908fa37459d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe8a54f8b7c0ac1ec13e98113d464c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha87ce4ac48b5eb557c6ff447198aaf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a5f2d700352f9af4b964a58bbee39;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc40f1a1231797971489c037cc624f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb92ee554d95cacfc7cb7a473d09f06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf36271129c02bbd196408821d17011;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139b0edb97f0be03749c214707a7d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130fd115bcaff01504166f41a2d4a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf14b9cb6b03042b64fe704e9b0616a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf8aa739a58f9029cf7887feaba400;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h582196ed054bc3d932d2a662779c7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102bc8e2135c5f431e011461e929037;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149f0348336db625b3f9976294cfaab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cd052b7200c30488987dffeaed9f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde8244c4c8994446613e883cb4c5b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4506bc2b1adc48b94dfae95f5be38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24c7f5dc68692adc3be0757540e4cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd722fbc33edb9752849963d0f4494d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12706340bc7d6ed38672eb53572ade3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h648b419acecfbf26925f876cba60ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb1f8e407a62fd61299de64fdc06d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18531f0cca3637aa5afd42ab50aa8fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d71c4c82c7af257f169ec997c7f0c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e545a97fa3b3cdcb13232b8735137;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd40ff0a6eae6f4bde3c4c74353d75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140667d63c47d97c53aaf161674ed9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b4baf524ca7ba4995de666e4fbcf5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8f977f8730b403e295d222528effa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10558a7faaa2ed171ad87a25ddeaf5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1324ee0f17c9ad28c2b004f06fd2fe4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102bef284a7d6074d443d1bf1703889;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de3ff25f52e3d7ae9de07cc3b6cc07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec551bb6c02fe145a532e8330e0f84;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15277c41087bb19d449beb3344d06da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf63c639f7c82f3591fd857cedb3476;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfff025c99f92f8170eb1f34c3fc6d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa9c29170c74becbe7b0aedefe0826;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aff574dd8a8fdad7a4df56e355be83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124f035488886357dcbdd555383b4a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ce2ffc75a054ae70946979ef7fd84;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7af59c028fbbb606d04c9fb7bdda3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2cfbad68da555e45632a8c22f73b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca94aa63a3b566a0d10dbd65bdcdca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3eb130c127aeb9ab3329db2bb0ee22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb6fd86f4991c72e77d8fb27ac915e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfcf87e7ef5a1f5d87002c6c89afb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0e2721ef82c4e70c62bba6caa122e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bcc104356f1104e945beee1cb941f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1182c7fc399bd1b8a3d0831481d8752;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd9b551ed8b61473907580f9fb27c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1312d30cde4b24d8d81963fd6310291;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8b472996e040ca23f044dc41dd360;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e3d5070a70ea456c9df49695e06f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0a9822d4d6e9377a4e8ade1dde572;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1293612890fc00b28db1f11d86dba9c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56b72a01e6b86a84a8433e1dbcc16c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13100b6c29b6ffd43da660b0f200a74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac3aff474da030a0e75fd71bda4e91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18301dd6edcb3636eacc5e9dea328fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f634c34b90511a27899c356f327128;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db25742da1c26828213ed0b7c8d166;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1998470fc4943b11663bd71af98e729;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa2b7704cdd99a80005328d1ae216;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1659ad228ba64c1225a94bb46c505c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hca0fb817fe3770f77ca5fc49bb502c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcca41ef5b73f7650289fc461df29f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h460ad795bd63940aaf41f21126523d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1847e4af3736897e83bd1354094adcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4c9e03b4b94bb8d126da0759ad17c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fbd7515587550a9b26789046865fc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4113c192747cb9b7ee4973f863a65e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h484578ab4420d4ac5c9b2fe3c24c45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f85645432d0eb52b14575170773ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h225fa74e4df245fdbbaa660e1fb76d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f835b0cf23c2e1fe0aa1269c3e055;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11e31f78ceea7e0cac49ab5577bd0e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d31d02e8e1bb3fb5b0c6c362fbaef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13103d7ca21f4579ebe4e3965a5c119;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ce8269380effa9a5a2346208cb9c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h529e5d3464bf279705bb934e30d191;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f66310d65ef6fafd192010c9088e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2b583dc0720ac370bfa9010bcd73a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9097c01544f89f7cb27464e8a9344;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16004929fb2f48384bfc1c358e1a528;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1226682a56605152635f8a2175cc117;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1642b2c7e45c9542c8445cdfef3a4f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b3be2f8c4d3c221cefd83134a3a79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h225227194ae2c04a0226e82bee50c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9c822893b8efce1a172d562b1181;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efefe22f3f66bdb331a0ce3dc6bfff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2636850d68351ea3d14926e73c50d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17148e6361804cf2d0a92a9f86f295;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9dd2d078000771a30075662b457c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac8501759cd831ed8668502577e56c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbe667c1cb95e8c8d57fe944d4f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78e2b4d1850e3fa5ac9c7e88bd97c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181538c96a544dc6b703900d453ec4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd1f1eceff2ee006629040132f240;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db77f48d91199450c4600846919ef9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac9c59d1046a7a0384ace1bb1b2b48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4302954b291e9ec99ef7684a562b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11fc14678fe3d7ff8ba6bd74627b787;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa65cdf5909c35f61d7002ece1bdca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149caabcf4ed5f921c9f077d2e83b47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a89cf5cba8a4bc766325eaa8b90cca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h874481e4ac2da242b7b6ea421ab77;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e13c9afd4c3e717d72b32ae85d214c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173bedfaffd752049d8b69078aaa46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he26e6cf18762c1fbac4b8b4cf69888;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136f86c0f3a904d15f993d146e5c6de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb79e4bdb9b55e1d740281a7d35070;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f23b9ca0c9f8cbb39cd63737683b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15007e7877bb163c267f83489efb0bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16baa6431d308815062cf60288ee72e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1448af36414ef3631d7b050d0e2ff25;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h177e4067999961abb3b68d63fc3c3f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e59ffef212105ab34084f9c31d2b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb2b4784778e3196945bad45cd235a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15deee62554ce2ca77325a261dfd752;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4e483e9dd1d85c82f3afa9f83da7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec695dcd37636553d3e658df69ad60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5f4b92e3eaa0c65124220a6210cfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b0d216e75fede04269e9a67579b11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b915cddd0027d09d8a2582b74786c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1e5203bd4d15c120cafc54980be24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc2faf186944dc0fc41d3cd44a9dc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14962e0d870f3205d976017d4dfee16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ea47bbfe7ab08e76c58da2ad6b9a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd91d3acbcfe9916cae67e7d91dad59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbed30627f983e48ff628255f36a0da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde497850d94b2785ebd9f83feecf3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h561f7bc8bb6fd59b45bbfb8cc8ea84;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a688dee617a53e02114d213e1c4adc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3344eb6e36eb9f1d23c99d09a84478;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h663186a90ac8923b6856703033dc4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb247fc084f9f7ecd6a431b57dcf643;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb42a487f0eae8f2bcfa08206aaa6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c660203dcf90b268f0c45e5cb2bf80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc1f14eb6844aa334378a1c225df96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb3f7f19567aefe781699f901c88c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1542a0de625a21c492c404fa7538a51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he334a366aee976b30e869e6301fb77;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b3399d601bd45fa600165f2e633b5e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9d393abf13b34e594c52f271ff915;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca718948974fde3b323e4a8e547f29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd073b671561a1dc66d88ca410ece31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h37d0725365a6174919f124c92982e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7548be8f4f765d68fc512b0214411;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba853c46c6f1189d48cd770ee79d86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44704c65e82bf429b749e2d779bf1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50310892fb233b1c6b2871e6103bcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd26f970ea280aaac9ba042053f8947;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0d5a7e9e7fe8b25376e0401f77254;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he87275928b788b289a5df15bcc19e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71f0d1e63509a590d72437e5d65238;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199e5b5d3631db5d8cbda2b6c4b7b8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9c3bbcc0300ab8465dde385afde9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f33a93a09197a2b3d30e23d35f0fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h794a2ca9b8680f63ef3919a9b61306;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7429adeabce8777332b04386ce42d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a89898e111f677372507a2c1b55b4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f7546a6768047c61c1efefaaf3417;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b408870bb8c8c464fabd660187044;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89b92d6fd6dfedcf1071ba138b78bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19eab37e5932e3cb91948972f830b2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a8b8934c9ca2e30071de5a5494253;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a9fa2bd0aeafe0c6ad9d064036646;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16dbf3b5def09e2d673f31ec7b0ac3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7c2baf525c3e3afbb1d5a9d691acf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8fd5fd4389de2610ec117b7dabf7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16dec28e6e0b016d433bfbe187d89e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13072088017d60d469c7eb797d43c10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17afdf4985a04a3fa078e3107f2ebea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1224196dbcec9c022052ea658f083e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd37004218b2f24cdc4c3ef1133ffb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9bec7993eff5aca2a7f95aefac075;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h525bf9171db51887145715d2a84369;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b5f3d2af004188acd7da619a6bd1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130039b28d42f2e1f16b7fa64d244ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141faf9fe414dbac6c5e1f8787a2940;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa59deab38767dc227514241da3558;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba565b7f5df6169a8ccc892944861b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcff17e7d1f567a7e4498874447c1ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc29f4c23a7febaca3d7b1eef435f29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33cfb224a692a94eeabf362810abbe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f1083301e33e759739eeacfb9b50e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0ff446e58ea1bea0a9f2f0e1d8bf2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8e133a9a8c955bcf2a24bb96d88ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4df6d53c8b1b7c62e3d8a41cb2a4fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3a58134d70ac58780ed67032c6020;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d2a6d6256287baf7525200439e2de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1301d1e9af775470b64ac4777360fbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2d094477aff85c11cd22d4aff7464;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1e73a1b8478e4826ab4e343ce3236;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd8e81945c3c1b33b7b7e68f0fadcf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8dc4ff9017bd25db31119bf0be6a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86a4c5cb895313f875cb65938dfd55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1b66763c753235699c5fbe0e0ba4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6832867d13762263b5bc7527652c8b;
        #1
        $finish();
    end
endmodule
