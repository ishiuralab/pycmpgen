module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c255af36b6f44f53446825321490f7ded351cbe79ed9c03df659e7659f7b28c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fa63e61cc6eafd7f6c534022589641dd17dc6eb25e31d95ea868557f765be97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fe0208aefaef1bd974769f0facb36fb9a3f3c8492dcbfe9eec335df49a9a90a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d86337e76d7e8c30976c928681701b75939d14ded968eafb8b2e38346db165f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ee3775e83ed6121753cca0ae5393d3d7115ea71b00cfd72a01081f85404e5e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4495f2a5becb5ee7f1ee50ca1d6430a51b17c75b0803e2a62ecf5a2ceecf05e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff36f59c802a23d35a064fa45e2c9495d1f2a4c6fd38e2e1ac3b4692a9558d29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h312c0de917e9c31ab4d839a43d1544ca273e108b95838858482a17ae3dadbc89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea471122123d0a39f7ee26821d9a6e1d611c5ac656ffbf05c37ed8f34b1ab87c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c01813cf13661b8115c25bc70524ff861585f36b18e8ff125cb0fe34e8e225;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcc42b691b6ed2e11012a65f7b024bd32c2277f4fe70bf58292f09b2b0879669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbac1af8ebf069f414a2548c4ddde22630da6c2f2a6a12087a8dbb392bb6ebc7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha971854388b854e2827dfcd857ed1363ca14db05444a4ca639028c11787f5cd7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d70c1766489409fe614abe14360db0d29a21c87e82b7653717d4e8b85c98297;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1ced06c0b0f84e586eda808a565695de3359122d337a2710a1bfcccccbb2152;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bb2bff76dde45318ae7cce36049e220fec13231c508ab07f9307d03f97c12c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14a1fd785dbd034e9eab061d3a8b5fc3768528dab505772ba4131e1ed34be407;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0765f9a271e0ed49139cedb5b8cd8f8606e25a4892de1b8f6ed876f15ff8a7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3e29c917aae64f5c37af68fb71096ed0d3b27726141906ad141ec7ce3331e92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4707c4b46382b9ecba487fb1980d31d3bbc93e74d3ed8720aabff3cc0bca7935;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h498180890b0692c3a203881fe2517644037435ce431285604f5e41744b3ea062;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ad6b3b73e1f879b2b13936e3349147cf5a574c07e20853d78729d7433c5a356;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf750720a1e7ba795a4de0a13dd628f0d1ba0250f5ba950bcdf9cfe6de6a77de7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ca05d3badc5ccf34acf1d4475d22793e2d71e9b03fd4cefb32556b171166335;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h402bac8fa00b348e62f6452d53c0168ee4dab6e91c7ee190f41f46a102e7ad3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9c2e9b29c3dd18f197a8948686182efc5dad107d4bc48abce2f30ddfa5b17dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4502243d39d670782ff8352fec5aa397894f6932f3491bf3f16cad3a1691b6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf4f29c31225d9f68553b33791faf0bd9dba04c3dc01e7193dfbd24e9e38c196;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf4f64fdebcfc98fcad47a570e27665cd4bf48fd2d2eef8f321b9f115e7cb2d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h554e39956b03fd1bd56880bcd17763fa619771e46e74ee6173b42d5a87b82d62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e3059518ea6ab809156cc8e8fe7dbd87ecc7e2a7a9700e531d16dc133e4acbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h470e41b4c3e95d8d23e93fd57bcd7852e226e5363463e1817997c1791d67cc3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ac20bee5013041f827c6ca2e42edecee7dc54a5f6d87a40f2fb8887565bbae5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb15fa8e5e8e8dd5431dfaf8b6595e5b20f692f5f0da4dcb42b97493ab42e2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c2d3165b9f43155dffb3c40daeec7fb37a54bfa5ee02d6fdc8e85ba8a793d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80c2978e87a4856e848adb08db5fab064bafdd5fd8d69fe9d9f8d2b7d4077c0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fd2e4c9f9e94d50ea1bcd3b7a6e1eb29808cdf31be307d869ec8a11fb036d57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1317a00f71219192812d1c9052af5f515e7400d5b73646787532c948b3101d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f6872d66f54b264a1965c608cf9d1a09b9eab40448ab10152d0ae0221451bb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h816b06d84e65d78a43caf54654518c4341c91a82d77c4aa3ff41c47019427cfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8bf9605bea9c4309a5b19f156e389926ca32cb848a010536eeeaebe4e3081637;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fd763b3f892c01c5b2b0866f08967e19b01ca2834fcab31b8b952b6860d73f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cb2eca6814f36196840ec115bbfa70dbffb21a6a20da9682fd19e8f0a9a403f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7928f469443a0fe29bcf9eeca3011a52ad5d6cfa1053c17c68989211488be7fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8124a1a1cc8c076ae32552b8762159c84855ba6f2ac4699bd816e4a7a5043d27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7c5ed3deca845211e1545354c36a077db14689eb23925017a5ae12b72488373;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h224a023443facf073d2f04eed5b0bdc95afac3976c0e9ee035d8765ff3cfbd3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc859767b3cf2e229f8a3d1d6f9964654bfd8b7afe272fce914ace8054bcaf495;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heaf4bf47d8c39e47cfd179bd4e2ddcd2c37ac9aa3c1ac6fd6569723b24b27651;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42f5786f85182e364a715f020419f9b81ef5cd3881ba6632eefa8dd9af60acae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heea90e511df2d73ee88ce95a49e7d40fcf426d5852788003be68b3538e1b1dbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91c070b59260be0060efca14b558f71bc8f6d562b8b715ccd804ab7fcdb67ab4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h520b532966d777c9f5e85c032a7895720a3a7f559116660ff1232c7139e527af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3de1bafe4afebb428cf13b7bbfe7c2e958d271fe4138371b98b56b5def3821c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6306c1b52e7f075982b5f948e7f68d188bdc63f0793abe63e30d416723496d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1793b460bb79dc999fe2979c022e4186e3c344b98279b690f27e5fbc9e2676ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fe06b296cba90f94213eec070d75b3b55dfa1735071f1822f6b737ca4e7ab2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae20fbf28976ca8185f85f6de2a754e2dc2dfff178d909f54715bde4cd44d7f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb30212543f0fc4052a8c715dc258ac5b4477a986df6d90ef703356b7d06e359;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb2d649e6ff95dd33b141a6ea0ce7c34a53544abfed3e72e4cad86ea3bae921d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h714d6ddb0f1d90a91530d0cbc139fbf5807268246460fed0af9e07a5787bd6a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8451b1663527c6a35647a33b7df2748f117a1b4a9430ec80ada68a243cbb97ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h753bcf51ca2303c0c057e8bfabcbcb60be164db1b85eca693310f43e3c7f5a65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55d6c407f6982a6b6f0b09321405ce5e30ba44cc7f7b10cf51d15dfe41f472e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea810626330239e8be370b8db275ea279d5d1065d104e9cc36cfd3ae7ae28195;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ccf4ba5c72da8934d0e514242618b1a03ee020b558b747487c2d3ff89ebc2f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9db4974baad18650800c0e7a6812262dd5f862ef91f5794f3895507c21217a16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27ef49127bb300366523220c8e31ecf2b05228de9fc2d45e6bebaddc19d174bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20fe21aee77a613dad26868b1ae09ef2f44e1711f13316bf7a0bda06622b5669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0847093f9eb01fe7cd0266bc37b7a5ac45ab7256048740ac92c76a9eafd2a77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc804ea6ad8d26c3b14e7838912aa9a4f6acf11cc5ac24b56ac9070fcefae14a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e267aab701e27d9fe57cef0b7cada7ff0553318c11307c5d18184bbacbf7793;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h283192b5c2dd5ebb471d347a4f401a2e15c345332dc730e3c99488f48a1460cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5693634b026a0f831186a8c1eb798a09aae37b03406f544fd44ee08cfcc18b7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d6ba72e599edc7f5c6bce309592bdb1be4709361fbbd278806097938655a834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc359ffb6a178df567531edd982417964f5045e4b1a6ae6487db78d1fd07719a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d27ba39143202dd843752281a91ad96919bc5b2966e7c8564fd6ac582ea2eb4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h284e243affc7f1f6036bcf49ae2f33b90a55b564133335bd9aaa5351fe849388;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c5c6d4a4294e5a6e9fbc2fc453d4ac0b4681859e18363f25d20ff0bf1b9a74b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc829dfe672d8c41e4f74c68344a42d6b5a773321716b5968cd948c07d4c2ae57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c70fc45a78b24da0c5e6aa3ef28a526cf44c5013b8e968e6cef30922424ccb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf281cdaab8449af674346922f16496e80ccd5a033bc090c28225bf5e77e94875;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ec470566ae83d7a990ba6599873e0b71b151319cff7f93e93f48cfe7c4062e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h205ed6b6d655ae4d1e0317128f2a6e62ed22520efd80079b99dd1fb62e81ed79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66c962a81187e3b4cf1091ecbc8f47d81c335d89c9bb2421d06414397a8f45c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5660700811709e4ed5c9548b238bde0420bdaa076ec21b07a336c4950303fa94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h384eb4b561327944b58a98dbdd2f4531f5ca8a1eed8b445f1dfe4d5a3517ab81;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee96223a860b92a5b1dbd0dc0b154d14d756dc7ac9cf098c6e73d2e81b10258b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11c5c3aff43c85bfc9c6622ea7c0bb043e2190d9cefdd88156e0b78bcf53719d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6598e87e1aa102bcfe8b2a1c09d6928e68439b86c740e15f74d7c9bc5f7fcc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h634e618e0b7924cd9ac59e041feef7b494948a72402b082430fd94fa8ff909d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha090cb8c9d0277b372959937faef0d67f181d8de0c398287817406c647bbe867;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c344ff4083ccd0fb994400b8b41668c09d7b367b1f4234257aaff0e7085326c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a93bd9113f18ccae8ae90e0b56cb3f689dffc0340f50115e855c33267931332;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67cec7928d96e05d6cb26a9d0bfeada6b14069d784c29951ab68b15e737cdbce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h900868d026b680f46d585dcf610d5b57d526a318b95629649b3640a99619311b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7d9b0dd04d2159bdc9445bc0a83170bfbf6cd355025a67417dced33a0dcafb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbafc8a9ab006ca32335487a3c9cef7b886302b54b96babea232f8a6ef4bb594e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60758486ba70f12246e1e4e6f9733322c86eea639b49e5d81841da63efa198c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6b494baeb6c42448221d11177a9d1fbe94ffb6be72684cb774ad2d8a45cf99a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc205be10a0d57c6ac153c8bc817fb3d87e9f3c7b4ddebd75fbd6291ed6962185;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcaefbe116676db956932d1b91315491d2946e57d25e3695621ff5e5600e394e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha02c811d086bef749586a07890d1298b86c9d17f8329e4abbb8e6b1c643bbb27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96f6d12f53296e68fb384f743057e2a552538730cad155b388639c565e948db7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d69796db6d54fe234535e6277c678a4c4844fa42e08d443d50557980149d440;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6344694192d08d4d57f5df794a82de116c017ba35e170d2254915a4f5818674;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb9b4887993402ced8fbf51eddba2778e799493d90e36fbefebdec5435a2afa7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5530d6318cf829c9779f2b1c96ff648a6de11019a16eaee0c8c38b351afb4e4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff6f0b320316d988912157a631222df1dbba8dff429ca44ae42f2cc83a517328;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf208849955de9ec3f57b2ea6a9251b13c56396732c005033dc06f2fa168c5797;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b2f0cbfc05780ddf05ee397ff362fd7e90d212593eb0e8b9100aaa1e05ca028;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84327135d2a225df63746ca7ecb6495619b13d14867937cff7aef450372cd466;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf67c5d5a859eb988be6519eba9542c73c7b2247eef15b3438b374ee43513c414;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaf7735cf508b52f624461e12ac51c410dd116b68791e5c307cb68fc4f19603a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69f585d53303eac3e11d7eaf61930b99dc09d3921de5a78913277b78e35b6b2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h273f7d14cb7ce7cac50aacaae46ffda919cd271a2ce21e200a3d1eec71cb969;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e07ea982b14be2a02b4b0b3c417e677b0b82ad169038c80418061f52982c798;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h642791194508529cdc22c55991a62f920e795a2f4700ca1a3afee2bece6aa3bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b7e65740ee76e7bd3471317a3b2331eb3ccab077a65fd4e8cd4fe83c2dcfb2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52c75ff3ad52a1ee571e94a88940813eea27281046fd2bd4cbcc76947aebdfc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dc207d1f9360d583ad37c30228a0b201387489c045d9e5980f2a6015f5bafed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44478e440fce4751a9cbed9afeb1724584b3c2c96d8c2999df8aa87a4feacfd0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8c87cd7cfd2afb119030243c5babfeee25632ae79e4f394f78b23611139dd51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbaa123402013e851df9f946feedd4ea9cdfba3fb138b70d64cbc50dc2adb1ca4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7eeac1abaa560dfc0e6f95fdfd2c305b5271f3657fbac1d45fc10ce29d2de093;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc718e6256de3d1c44ab5685e49a16c3c3f803332fc072c1c45a756f87538f419;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21673c6b285ffbf8bf1f3f50a920e726b6c04667be32867c322b93f32e995a14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5ed6710b22ae8ceda22117408e5d06bd4fe630bd76e41ccd064e0d3c516641d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8108a0395e0ef5847e4b0d702786e99af2f6d4c736e72c50720312f85080480d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha638cae15c23ac932514fe8c9d9a790063a4e9fa3e3c88784c7728148f90061f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb04a70452cd4880949016f6beef0e9172a03af721536c8b9ed868c24c1572c79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f8ae40fc4ca6f681273d3e85ba0a433929bb6ec6ccb2ccafad08767bbf25a3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he24e3434a570f21ceca954c83fa675d45ad3adb06be99b6a9434048d01445866;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab9bad0908c020a213ab51f0aa76386530d60627c1917f2b1fd415784f9c275b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac33aa0d0e85cb3cff6d4fc9a376b8aaf7c8c4f05a6182be366f13ef7b737d49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dd06362cf4643541b3f4e658084a775bec25e784a1648edb88f28d0553ea51b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e8344df686b818b30e87fde9d2a3f816459fbcae5bdb328a5ab0018c11a9c3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd0a24a46013a4ebe287a789a8933b90a16dff73889896693e65e91b0a80e769;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8711d5300470973f31da594013fe0be3630224352a947f0cdf8ef633d6c2b46a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h261aaa0d90127aed08992f9e3655b11eeac2180be95a1d83325159b114f4a4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c1c0586730749190967a894790c44344bd8d3b002ab6d503148a3ce55b2f076;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e89f936e9ed4c9eb3bbda1b0bc14a9a2242ea9d37ac7dd78bacc062786f6f8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h282b6699d5678ecc494e3bbf31ece11778a624f52ca5cef2b5c62a50b664d4d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha44924ef24ffb769f6c9ae828c3768c497cd1659e03cf85e676fe90b07382554;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e482a8086d2845333610cdc0c30675f0a2dbd5f5eec2a6d5fd2ec201bdc1dd7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63d3a79748b2715d488fc9fd73500516a538d7551deb2b546191a57534def5fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8d20985f6af08aff3fcd5c721333722e4707f550af7dcf80b9d38bf8b347c65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h324da983a6c171428116ac62ed4e37023e8b04a85653661f45e3e267de7fb3cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5b3fe1ee883eb893576388828228c0ffce7b15528660a7a044d8f7fc7949082;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h195ba0c8069de394a66244bd4ec8ade04319a63c029db1c2e6a3beb99c76f961;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h413d58e157233ec6b923d1f4b65b310ebbfa5770bf441f4cfbd5535b941d1e69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf498cad438e2c51713c979d204d807711d77c21990abc8bc0b089581b7c49b2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha52b2c29f423045fcf26dd15cdc95d2056fcc31f28012d4c0aabcfbb1253d32d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e8e920decce625768eabb9853e04f046402707f7ba0c231f4e3a73a8b7100af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a2793dadb8d91b38f99022c0329c8480a7fa34442d193b3fc622ca09ef58477;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47578723609a373695b79761486a614383dad67f23c0d0e0127810cffa0bd9f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85af56e779771d4ed44f7653110d16230b62a3c4a127ba264e5471f9d5080b9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0905bca12fba44443b2e7d4921de1bf75279b4ea368349f4f7818248cca6f6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b282a521f239e4c66d7d39681d6c36f9097eaebddf5aba43201343f56ee7da3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f967b56b547f841c867147b6478efa3be3ea62bc68b7e1a64be891818582a74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2eb86998ddb3fd4cc0b53977fbfd26b73eee992041cadfe8f26a70b8be81fdbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26e4facc7f5aaaa68667cf8812a06f6dc531630d12af734bd601722d318a62b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2237a82bf18f38e6a74889eae2e2f482d216dc1dd4335cc5f4c6e7acfddd0b83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f790108f254cf6a47bc7eb0114452c87e8d909b29e92aeca4fdf8e80df5bb20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4ff836e84843738cbb56b2b0143480ec2b502678bbe40a0eb27d13ea76afc67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h669fd1c5ddae196cf69c68d97c66d51af75b35eef2e23f083d79104c892fbd1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9dca19ab67057c32af1395a9e5ce011e15d38e9c93398e90b0f702f03e85a20e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38c6d369aa6bd36040104ab4b34e662d08c1589e1e1a96c0eb45bd3df8e09145;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7add6f3e4fd99bf11bac3e209a0ef6708f90a0659ddf078ce5baad3210e71eed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9abb6140d1b5f005a5525c68a9826582f0c55421b9df899c8740b06a1af80ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69c4bf940e76f6367d36ef9758cab4d90902da7bec9a55df43b8a033f9a29f1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85467762d60e99d08f7d12ff71892422bde4b7a8ff78868e46d5bb49281b17f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h559cfc76fa9ac2bd495320a4b458b985155bbf3599ddbc913b8a4c97cb3bd82d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ec0b7801808b231628f4774bbf113d09862778e5ce50f3623e7c06f86e0b503;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd65323621399655e7f997e45a2d2c48bb712275600f5695b26c445a008c76a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h961ed126b7dfd073f891e4ed49f9be8dc20b3772ad7baecd0c75897f28f6155d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b673765d33a9eef75356ad9c0d2bdaad9427c9dc234085a48b3fcd7d6784f31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6241dc7f4ffbf201984e8a317657ed8a83de11d895251b169d39556ffbfa1497;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c2bbf1e7c923b6ce545068b85876086fde563405617332260ae37aa46ff0fce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7545e282b5f01c924e9f9d2849364b3aad668e375351664c5d5e6c74ffee9d23;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he966175395431fe9600b30874ff5133effa70db2e37a38db256c794a62906115;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72632316007a766adf1b49abbe448e2684c63c8ea98271b903cb7ae7425b4689;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h256032a5af65c9b944b2826110c552f0feb4a04b5f5662327ae0c4f04772c4b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h789b13ab2f88901c75bc854ffc28e3678bd614a1588e860ec746c6460b9679a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16c2c54f9c1c964c30a64ca868346c8249f73634b227ad7c8b7ebf74fa36101;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d2c7e3481f9c652a68183d3599c3a250edb94a61b86fcf37fd970e013cf6c44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc964320e94c3e6bd34a89dcf689831f69dedef421457189550496b3dfe5a99a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6f63cf77a37bb6930b942a3bdb0c9ae85addd2b7e1a75959ca3e3bb0ab5ec82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf667f0b42218cbfd1a1b2ff8eb4e3694d6f63eea029313594418fef4cc026969;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a30c2a9232aa3a1b6407d814e361becdf56b1a838d3b8a0e1d4321dcf099912;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha06c50a5480b7cd8170639efcb3cf77725043abba7ae1c4256201b9d1f80e523;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70b4f15aeaa500bd78928adf09d7025357b625206c5c9d82a3da7e82e1b087b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c0c6e9ef6d8f4c055dfee2e28d08fa0ff932120232111bd486c2d4d1170e60c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5353b9d0a6831742e26cecacbb07c0215cb832b111250b466242c04f40ebd452;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59c8ef4fbbc228332bacea801060aa53fe760d8583175f7fbc317bb1e9d61bb6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d2112509f45ec9b577b70d7d8836cc0e72f35ec82f3de0d75b79d331a15cff0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80aba2f90fea9af6b37e38f7e6c56eb9882a3eef9aed2b3d5628d8d7fea1ca16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9c4e06cfd26b7ce3269e971d1b4e2319974e9e0673cb14f6bdfdd0fb6f2243d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76f76ebe58b4fca8a160ba7d5cfe9692659e4a4e751905e549be646403689f12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b349606b4c4dfa47aaa1836a7a6634149a2b23539ef921e9738ebe38dfc768;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf18001a190606fa99f60f5349c97b0fc6afc75c143ff4fb3f2657a44fb764f64;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec39acf30362510567ba886831f574cbb152b883447fe9bc7a6c08ed87f22fda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85e961cd5f5558f7f39df9d3e10f1421ee7dae4c91e12edbc801af0336cb06f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc34689e74ed16c651d6c474abfa883541fd050c03c2ad17ddec8ef667a86ece9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c92e83378646f4007746482e7a13e84c4b9b83813aec6ecc24b502ea80b3e57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68bb8100dc4e7a669dee19c537c76f08b8a49dffb1b0a546f477059f93fb0ece;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf51e68c3e6b7fa430a0f2e43fa8fd3e067985f83cf8837964d98d83d2a556608;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30556844e054af43cdb36ed56117ffd7ee040129accd1df1565aa5079322898f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9760522bea0ee82ab2221a005f90923f49092f1983509a2f42a7baee8f43589;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae82904a56539f3824801303d8740739376387ce0990ffac55286885b6682c89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h657a272b43394845bac4e377b772aa4bf964b1307d20ae5f486785dde2d803f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb115261c01153faa42c5b26fafb758c7444730361acf3af2d94e04e3a0ad13a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b3cd360a5e52a8a479b083cda71dc9d35bf68e2eb38eb7e7e7105e4a4d8469;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h646adf7d3758693abe5c3bbc3ac27c22ee3dae58186e7a9c9c5e7556c8902496;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75a0c2858aa1dfca7d13ede8a1084f4910e2f5d88a495f3350cb3e1f92afaf94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha71f78d88b1fdcf713b98bde7f687c7a61f4180449e43349d73815f9146c2adc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29f31ec6c31eb98a40efda864eee8b5e3de2af97b59aa662cee977318821273c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bfcb776cd5ca116b2b2ac12f64414060cffeb39940803bf51a70fe7c9c94bd2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f774187408b799747dfa3374a3306aa0cd2468e096572b5f2fc71e20698092a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97e722f457048072902cab3362ade8e7acdf20412237e46c1c94927056910f30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2a33d6bb84d24b3bed99d0c09609b5e85ba014c8830bcbf75bd954cca31cb95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a8c901d0d03ef3e2562a45cd8a552369c6e9d5424d17a478819a09be5304e4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0f3b756b310d650926d29560e23d83d5ee730065eeea046edb1990fa6bf993e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc91aa3258507811cd916074e07af41065e1eca6852c39f97d84feccc88ee2996;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99cc59c3ac1421aa513e8754d3c9c53d8ae00de82f2e975f6174642238dc9485;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dec2019896ae3dcdd67de3bb4aac236c063a5b6cf319d268e5c6c48a62152c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc64e80af2cb14eee37951521534008bbd851e17d6bc268152a8c2738cf49fd1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he681ddbbbddfc5040fc50958050888d70d1601e54d56ff3b38bc6ad99f093160;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2feac364720aac1064dd80c69a293c503a67aa9c5b3e1d0d8ee4da013ea6223b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4a921803d7ab9b5358ef0eb1ffc71d947097abe080af90d9f09bac29f77635d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3026449a54c6c1ce71f2ffe4c8a8d2c9b457eeba5426e708c3fd5519887966ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h690d2e95bf494fb06d0dc7f3f8b71eff3bf519b20c8ae4d5dadfc977e9a10025;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46ce597efe8a7a6d8060803880b6b3f54d80b244d35c55ed21cd71b08e25eed4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf68b3c2feda44437270f94ea3894c748ae9cb74df2e2ac93d4d293d100a0a0d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40a8ad62ce46bf6173f99749be4ed0a4a51c4a0ce1f1e7dcc0698fac168f0971;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37d3f086ae6ad0294a47c2e168b597f8d181d59a1ca8d1fe3afa163e3a529323;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4ddbfd89ddfc1b673b8c72a2162c024c83d4d9a26d241b505ce1e370ff116ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ef603f68213367076a09c9cf7ed14d367a192b05db1d67cdbcb8d4add09e91b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c22aa621d08cdf1ead1b7d47dd9ec2c8f9a527a8ae4533bf10e0e4d384ff573;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd26a6b31cf91f539e1f5bb560f63e4b7d40485c4ab468e3c0ec135541a7b3231;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8fbc1208b03d814792a92e8b9a71946cb63809728c122da66d6e6f327574a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed3aaa6ebb2c02902e2c47b1dcdbb7111d6e606905065252fca468e8b4cc63c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7cffceef399aee4bb62996defa3e94335fc4860e86b2251884a32fca6894ef8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74ffddb7ee1c27b075dab6ea1c1d27e3d33d5e8ed3ab0f47350eabcfa0b77ca0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3f7a7e15a7277e7a069f6124d63184df527377ee21f5f807d0a65e87b0b24e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8c6db59b042ace67d317a8ac96f00715323afde2de66bbf128fcbac7ec4704c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24d3bfc50a8ae2a29ce82d78c515a40ff023658b14a58fe13136052a05fd6505;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb564a50db6e0c21a73f2f3fce0b5bdb2584275e98ff6f751fd04626191d4c3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50872b0a0a613bf191cfa2b505b83246e0dd122b63d5f0e3fe798ebbc8400906;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc69b391ccf84a599fd2794741383b6f402db661df07315b86568e0fee7411a53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74d2713784de35286e5a4271859bc4e07bf9fc5a72584eba3c081211ef69f15c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd50c07aecc34c4d153757dd38e5cc0e7586639c245d6b576e0d74df9ac7e8501;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44025de994bce13adae8ff6d77d140feb2358d20864e24bb97ba52f47d225729;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6eafc2cdc78663b9f56cd2b9d970d5377d8b6ef7ffd38d99e008f53575e39db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc384440a974d8f38016414cf3b054559b83fe86399dc662d25e085a5598a0f0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc40bf6e988d45d771b2e8ca061c82c219cce83c8ec6b2750a00f41d3c2ab8e67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h853a74efd033cf46ee332d7d195e600d642e4f6e5b352dcf1b493d4c46d131a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he488b47c87bd81c7ba7f7deade69da6da59a5bd0848527c833e7d8e03de6ea38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h954abb723046994dada5348096c37e0d7edc9f824ae01dbe3be106c8a4ce5dfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59863c9659c5c29e253d8004561f12640020c302d395379f7bbb6ae5f509cf56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69d5d934007a26b62cf77aa4afb594cc5ccf57f5acf727ebc372019e786f18c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a356c94fe282c823024bebc3c5d91cd310f858de225978c89df8c5e6c02d266;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfafa1967617d7633e9bec270ac06c7b55d8ff8f5df1c0b20e9c398fb4e48d99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86ca80dd17183a8fe9372c25d4c2cfea29bead3ef24131dde27587755be6c40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdee88fe0bc78283c6978e49fedb9099ebf9cf22535324c9c6126b1d5008b116;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd974be20f82414d411bc9376a670e2f0b311fe401ca4d91e5fac9839c0b53284;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4b95163b1c53f0503e9cf3d20a05633657996c0c79c79253c4ecc5805813ca8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8c3e9cd82d859854b1122b27b01d27609254f883379006e9e3ecd5f493148ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3c7c4f74137f70cd449d5d87ba3633acb5b959d43c0555603563fc1161959c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4af6333d00ff41a98e2e20a8044c3d25984204163c58f9429bf07ed0adddfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h374c2bce5eb86081f34d164c1c071c88027deef5aa55d777d7f2811a2c6c47c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5d9cdf23ddfc384e05af9122c717564b60f279a50d547177678207977439abe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h580ee6277e34be593b8dc3d2905b09d1345c8417f41ffc60fe403f1e257476d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9825fb3df23e9c8a35f4407430d2708dfdbc4d26d2679794db2b979eda0a22e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha09e93a32f76dbc867ce7c595b7a0148711401cd1b511bdf397d80d725a8744;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a0caa85b9b97f103097eee1631adc6fb11eb8cf980ebaa2c2dffc1398ddd8a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5596d5ccbec64534ad425770d84bd333b5ec459607026d82d48e08b57768d1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90abf1e360120a3b1b6d6e5085a767139bf27c4ef997af49f19436aa07cb1b17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7a3598c161adc5364ec91e0c9507e41307b41d380f582688f6d87e941a27e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1276ac7c78ec59ad590f5156c6cd18b8a0aee0da8754f3fc262495fe7770d926;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5691454c51628ef4d1b5696aa7021ed7367d42d358d9f2f86fe78e42e0935276;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c772919bf3480d6a4de2d6bcc2671fd89c2d08a66a6398fbb496de0f13049cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha204c194092b17ab36c2075a7c109aa3121fad24936742cb9700e8b0fcb36794;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf9d603cc5f555fd2ec21a18a2653fa221b5a0f7d50498cd4c9f7f4ee3e2ab9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6d354a8a3ab09a9f19d1628857060251a94047bdd7255455ff4fbaf847f5238;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda8361da87b72a7d4a21aff7f440941cc5c770501ff3733da48fd08096d14ef7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f842f90bc9647c6b27e214ab7c44872434248c27ed7663ae58b81b8d2e1f216;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he493aac09ca51ab8a38ec46a0f35c2170bc09c5731d5bdb19d34dc528f1efa94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h236c3b3c01a52f851b669cce6b40b879777d91eaaa2cf5eefb0fd299b4ca7e71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a916eaad368435ea60f2bfabd71a864d4a98546aded8bbaf7a751efa0403bc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21d774572d6099e49ea7cc769b571a056b2ac4933f1107d4a5f6e26129262a33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h506c6b69df89be99cc5b431be026abf2e0066145e8f9d3ada2b6d29748702f54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h142f78d51e83b72575f9f0026d59e89d890b884a6762ca59ca8303f35fb4aca0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbcc05003ef0061d004c10a814ca4e12afe232bcc373ab00963e860611d74a02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b0a9c9bcca66b79d892636d37effdd8a625c67613f41aedaa9a14b511da38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h762ba4f2aa2500a1a133036416f8cd3e385f34bc5b530f5cbb6aa0191a505751;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31e6a65d8ee0958a1b3a41779e3d438a6e240efd1e04f40e22fc991e47a10fed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9ddb49d821a4f9b6458c388382e2fda91964f3242d3c22a2eece6112440c5f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2aa7c3641a5ca2c975cf8ee42a69438880c76c27d4c152d6cc8defef89a5bd77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d42546c87dd551885bfe9689282d783fa532720bee12e537878f2fc790a2234;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ced0ec3f64b873fd914b4e108d448d3530038bd61fd20b37f447985166530c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadcc06ac4bd8d5f383c729a61d234ff33be5de5c4ede7fe3de02bcb88be8c293;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h460bb46201582fca7c3a2b24bf64d2f9599ba774152ba7510b480c5374f39342;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bf7b93795337806393169ed2ba9b2cb447ddb193696832d0628686ebd414f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha60fa4959f6f0e05857bc30b8a73ee42ea03dff8e81444109fb59b7fa1dfc662;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33d75b22d0b90c26995afade3e5d17fe41c610886b0bfd1a50e05885ee2b796b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98a4c2adbec42a2e2c6da7495469e10b40c371ee35f43a5e786986b19a9de8f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35ac4592d903d1607ae88891aa1bed79d186ecdaff5ad76953cb96af62bf562c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b4436c6cbc98fad8352ccf775d84227017cd078fb1debf56c559b9d0c5ca111;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa490453d5472ae7de9d27d0a6de93019cc24ec600cb1b12f3841c3701da5c9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98d510ea1861c03f8b1b1cf9c6d032030563826f934c99dd7c6de6d9acad537c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h593c0c34a411c2bc43cbd8c0d552ac9917c8b2d24c80b52851451e15129a1bfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc6d1921f65524546614ba4805c085ebc917b169f1421cdd6c83e34da1589e76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h243f26a09e95ea986f52aa18f3379b54a226d54ef11381595e666edbfb3308ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd58d7f317b35d8f7174fd2f49e8a6ce18d42fa320e18848a36574137a68b27f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9439e5ef6f4245cc030a109ce28eaee0d71f7c758e24e28923cee1dea6499ac9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b0e44909b1d4bc94d0f365a8e71d8d162b9c7e9f6138a09069435147009176c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf53a6fb2d2a99ceca0b2f38ddd3ad0f3f932220b20d3495dedd627ece109f764;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6f687b6aab6e42e480396d79d6bd93390f628b51e64d6a0a77f172f8080816f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he540814bdbbf5ea3530d0818f0610008cb94857f9c4d2b5548da5391ca681222;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6486ae663b67e27c3f0acb051e8ff54b2e0097730effa97b55ec452104f122af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbea9377d0e664835e0438d5e6996acd0635f419252d34ed77168b6f1740c362a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h750cb0658aee79a53693ac85690a6e9035fbc521f7d53386ee5b6f92792031e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h750b040ecee5bfef65fa17cd2844c0eab79479c84a95013d7caf06eef1f04a8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8888c7ec497aa3f1a71e2f1331c3b69a9d468f01274cfe1dace9e2bb55735613;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc5643c0faeefb8afe60691eadbd982b3cc167dd3f6cc0d2b5d6952dfb8c8fe2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11b646521ea9f23ad8775918df1a1e54509850a34309a44ef916cb9bcc7ee781;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60d9b5eae2b922b0840156a12119dfb47528c38310e4ee031d3e9710209f1828;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88c32a39fa4ea85dd4da5785619c5e2e38543512143739d874530f242c0a0d69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6a1836faab0b230520953a946c20598d8920a337156dfce2cc0c66eb027e5ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78a19bb53eb626803b9b119795679916bce0ca4b18526808b69e902e174916e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h863bfec6dce3ce6a8dbfbe1c459eab11e346b8079e0c7e940a4e7a2b2928d168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf283d4e1aca20585bc00a06085df4eca6a74cb3475846a13d9f58d10d17309d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3bcc33c37bf95782e6b7938d56f9ffdf721252692ee09d1d5158db52ce57ea8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcbaf993038a323ba9e4b59cd28e02d7a6b2a871ddebb696b6e59da64f14bb30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb722eedffef5414fb94fb29029cbf0c0bf007df952ae811606b9d2d9375c7474;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b1876082088f20e40673a23d8af58a4ada600f7608a1401977084d092bea9ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h288cf736a6582a4ac4fc7b222f7b9cb68a8b5e822ff840831140a619007b2632;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfec06f3401378a1a922632d1eecea8e771fb68f6023e5fb7adddcf5df46b694;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77b2259c7d48dd8c2a24a56290f8bca913cb022df5bc4746bcecacf8dcc9bfc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed0a16b9364b6156f595b42fe070dc152d2b0b813aa65c3106b6a40708c1711c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7662e4265b3f31bb6a84e8d37aa170d84c1c2a2957afaab07bd89bc149df2211;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a4594bce6ff74484cf32909056fc1b172de58040c35c476f3a3da4a365ebc4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f478738fa1a0c687f37bb6d10a8cc2fc4ac6ce674998bd8dbd1fb2fe5d011f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50e32643d339b4c36adfff7e5bff03da84813da0e549f3d9f2f2eaad3dd99745;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b05f327ebfef0195fbf478077f74257563797ba49ef286d841012502b7ed16a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea3d8f30bbad6aebdff94004af6b6b7894c3969dcfb3dd612778603239ee8b96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bd73b684c7b2357fa6ad7831167c21e980c1be8f20183d7ab3ef660d837f009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4be04156b14b5e390f609bb2d2695a2460ef8b4cb0d13ddb7490ec9040720f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72f6e762d3a8e797c1247cc0036d8032a43e33c96a4065c0890cc6352a229fd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h322bfb8a29af404411c04a45e54dd4ab544f21f86438bc1f979f9d49c7a85916;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d7fae7aaadc4789325fa4c4c2981ed54b50ad82ca05c893a9354d9098aa3b0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha73efa85b44e34c6b524a2d5924921c06337f26d6a81d8c2f7d72a9ee249f0db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc029988d45a9a20ae4da04df3dae50d6f101266fd2846c3286f7365cdcfe0ddb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13206af46f071754b329ef27c81508be7baae988ffe81593c75e1ba103dcbfa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2eb773d9cd9353eed02b240c71bcec82b065fd2731371526f5ec9cb40de22fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha653c99b35ce0fecb0cac0e9a5d1c4fe16ef3a2236c1b91dda4784be3ba4aa9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fd08e25c9f14831bacd906d28d48445a1e544aa9b5416f371f45593df959384;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ae3fdbad0bcdd2bef23ab23e8b7b233f31d9c8cabf43c30ee6a9e407c43468c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fc4e9a1128b683af1d5f6ea8aa8d0a40a91dc5e6982702274aac4fe20dc0067;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf1a988a11536b428a3ae091ee080bf3a57ebe8b6c0e10d12ccc08adb87a148a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb81a4644debe1ba5ce80f5a196a8505c0662100d952a57c360c15e7b0b5b5545;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a54e7839fb925fde3a37846a3b1c654b14c0f5990c9e2cd773a954832ea2746;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c754d57f092346f6c65ace9ec4b96cf0641adca404b68c00500e4a6cf86e5ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf03bfd7c43a4415094acbf06883f64dd10ef90e52bb9328ce644d973c7807c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd2714749c4cdb85674447b99bcb52f8d16c4e7ce69e684dec6a567bcf1960d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c8cf1ad48362caf82cfb621be732072162bf2e51f652b2c744cca83d28871d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20f1ecd81870efe9ee261ffaf3513542f799a0fb7e8a7a0e5b2ab56ae9065dc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5589f607b938be58a3d9b33976cdee44b8a0de4ab02ce051ddd47b22db4ef31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2d1b8951e23f994fd6cb2a6c646abda75ab0ef21523c1e6a61e931fcd8ed9a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc3420c7ff4721bb999edbaa631dcdf7bd9d75e9cd44119adb008d581c2946fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h715798afd54e9d4918b7122a9759afe76542f2b8b93eccdca41a0fd55bbab38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6359755514a18d8cfb287144a0251d11fb5ae59f9f9d257a38831b2b8f94c70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaa5537e93c3204075885e7ae7b21efbf0a895902168b6add578a70b7aa592f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9968026dfe539819280ce746c7304a3a17372f8b8df1ddb67d76e83d626139f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93237b7c7b297c9cd49f24f61214ce76c05f448a66ffb3bfa74e0b82a231d56c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9809fa041ebae3b4c6ee627496162ea1f916598a47bd67ab96f72987c246dfba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4301c4d2ee4bad1f5f9531c5a68118528b32a8f81e6369f7d1384d6f96c40de7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d33e9be6d53304f62fbdcda4bae02d51feab429fee7df3b6cf5dbe05747613;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2e5f5faf6c8b5e521da227c2b1b56e30013f63628aec07572e7d3f63d35d78e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6ccd58cea1ff4808e2ab2bc8b09b248c89c84f0fbcd2bc13544f9c45567958c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf7ed7be3217fb8eb6ff29ad49fedadcf5213564b23851adf35d8c8f7327590f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcebc95a29a549b4b38b00071dfad926a99badbb857c94080094a7582baccd6d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60236a6957ce324639a546ee5a4d74d6b9253819b20e87f0bd0d058bbc3e990a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he637afbbc5f5714c60a46ccd56c1002860bbf20bf9605d3b9ba52cd91759aaba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7a3208f38ac768e16b875fdeb45383706e548c1e0281aa056ff61f426362e19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d41912ceedbb803e2c9c2ba859a40948158e0c6978ee723c0f26f2c6fd3a07e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he280cd58b487447c0d7c2bcf351ac397484fd011954e89a13e5d93edfb1f853e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc610f45be6fb9801e57fd9cca8d4e90770eea3578959419ffb84073897c0d11a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28f3c0d1e6c3dff0aaf3f4874e7d6c5bbbc63c7e9832b3455763e9ea102b52f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d9277adbc9f9ea35ef87b7ec06a9afaa71d4020491475234768ee98ce4e7b2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbdb8632694a4b1bd31e794a65f92a0c4f49a3dd42000c8d6f6b5c80e0f5ec4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75176af679b2f94a549a599a212051839a026d1c69e9eccc71b0c09604c1c0d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba507618502007f72d5087345f9641301b13d35f727ae4ef7ffedbacd78c3834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he99e93c24d0f356cccfc0c445a951e77971c8c2dcffea11de59acd341fb613ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d00df772c76708fed04ae721d40cd2236524e9c2f132a9ee41889a2ee41fb71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb54969f9a855a84664f5908b912168400bfaf25d7bdfa4616c7e4ed13b0ba9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b5cb72bb023f6e6f39fc1241873127577cc2944850a9f81b92c98be6dd37202;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10234082f36aac2fec8e9e4c2ff4034a36b8132bc432129f4e1ffa8d8649546f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaa74a0c43ab6e0c08b170298345f70338dcc016fec0f1a4de978ccdc6069710;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39fcd136a34ebe999c6f88efec3eac21c8b4371472118d816bbf5393f19beb07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76047203d7e7434dbfb04dbef42009a6165247cfd879c0337ff2ae17042e95d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4124c3699152de8791b44da13d3d2d22d5cf4590e624f1f08f23d56f6b306391;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d608aa5eeb6622e98b435b5e907128bf65f7191bb245d69c6769267789c0ae2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74b96702213d9b2120a5cfd5d0ff1c3524e9996f8b9fa22e9797745ad8c37ea7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4b5ed7c23691a9f2820100b1a2c2d5e72ef14dfd755171bf579c0aa38324906;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae6993776539f882d26ea72633fa620e299c66e0871df5d4aae5b20041388a3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd6c6678eca95fc9555deb30cfa16874cd15a58c04da3e37a94e2f2d5903e4fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf2244769f08bbab686d45434adff7ef23f1f983fb84c322003901f0cb76f5f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda9cbcccd55c3d079969d6e6fa591a944b30f947ff31a40fbadc32537e1599d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf97e3cc5fb29303f50ce732dc4de0a10f502fea185cd3c0e19363e721fb832e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb54fbad32e966609587593d9e89bcd2b724a6eeae7aa642ef2284e0da1cd304;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36171e1595d214f8debdd860cc6ac427b87c6d271331621bb079bef6af31078d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40eefaafe6ce4294458387dd0fc6b4469592e42614fa0fb430f9121e2f556510;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41ed11f4a60da6d137570e85aef4f17c915d065b16723027f2e6bbd4a091d49a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba005ccc5314b9d8208b9e57b1a43f6ec33154fa0956912f80abfcb9df8918e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4dc0ae49c9e92e3b439df1fb5aa997061bfe3db5935c6d3b76a590c0f46dd815;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc355f232babc3b2953eaca0439a29df16abfe153036a482e273d79522059b4b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b63d233887f24294f4e24556606b319dd24532c6c7b87d801a3c23e502fe8b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53142bdcb6dbfb506c3fcb66c67ca01defb03a23e7f6cec7d8b2283ec956b1c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83daf36accf075d57dfb90958800382e343b6a67355ed05e1ccd3055d8b184ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab25c7ca7c19e5e8bcdcfe53e57557ea8500120240a847024594b2162abe33bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d28d833fa254818476b1ffcb745b45b49172fb808576aa6269807f5553a58e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6c8185547877982dd19f3f2beeb61987f1c56597cc4d9a554e2a74b69e2f9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h674fd8c85ae525073a1fd91798eba95d5fa9805f77cad0308b77eeb322bf198b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1e95a7eb496a1138f5a989b3f0b83852ce452e1d1d161b5449fbea821124d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0ab22f3cebe385f1ad3733506a7d7142878c42f6a30d3c7c184dd21a40594f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5381188c206dcf1158ffc34a06f395ff2f56430043e740785331b27763c7fb4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9705e3494efca2fc175f49711cf54e46c4638799828bdc3af18120e85d84d7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34154b1ca4eb5f2f9d6956ec2fe927297665bc70e04dc873dc91e2e1e2cf250e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab7fc09d9ad40e75b4585692bfedb0ccc433ee98f68bb457c23e60e680cdeeb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b3593701c958f27530e55ce0cae469c01aad55f7a4a9567b0f897d518b74c0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2cc5905047095ae7179d636aa77236af3b0a8533911749c1b2a500b16ee2903;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedd78a6e4995c8e126e6d688f3a9697fa0c5894158061c5975955a3d9aff365b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4b7d70247332782a5110c61c10d97970f8c44626cd83f87132be3a90766a652;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b99f8c76a2a5584be696b5f89adfb2f0e5030f55c144436a037b0ea6b128dfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4fd1a65f6e85a96b5e0c571dc553534a3feeac02638026b473acc260a05d84b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38269836d4a8eb476791bd9cc36349a2f9e98875ad85e1ed0e6cea381c43bd9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe00cab22d3df912f834eb26952321eedd44c9a8c066d1db3ddd7e5ccad90ba9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbd8997aa97034094489cc531c49b9c551230d85d1e31629d23a1a6f9d302e8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a7ae265850d5aabeebffc60b270d8f6c7c078231cf48d3685f630dbd49c570e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd055e25d762f820954107ed1f02f3c8dcd2c2161bf02c1bd29a30b772edfc30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha82ff722e46275a04c665ab6cfa2d1ae46fd8ef8a457b2e1ad17aad983a8ee39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd776740f4516a4e4cf01ccce0a13f315c2d427a3575b6ccf612294f10f209fcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b58f90e672fd8ea407f703836f6b36462ecd5cfa4ef315f87c5c40278f029b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10b1e2724e4d06b0de5896d5d7ecc1a2b1a6df0c8bf7b67238840aa69a4df355;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46540a2adebbe068579a6393936445818d56b588fb4562137aba5c2e2614502c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc36cafc8a8db2461f0db8c54e13a5c8a7c67039a713f2df621be7ee389ad9cc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6d65c961a645c82cee7e36d8e0aa9d722f98db5d0607fa7f7d1cb80981acdcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb919681e108eb8918c148d78953386bac39010a21924523406c1cfc406d29570;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8691c3081496edbbac0f50b17962c5c658a2c40e7a06f19a28e0269dd2cf0443;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8615a1421649043fdf1f64aad25cb951cc0a04f4450a8bbf5a827ad0ebe6bcc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6670b46e224fe57a151db8f584414702762c967a495e0f0872a4f6c5cfd4e31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92fa6e3ee8c9b73cbee1758bdd41c6f675422f1de1f8c233a53f8d276c65a51a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d35eeb6acc646689d0f38f6acb337dfd6ddb72f8271f37662de514b87d18373;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h412a86a3f15191e00d541f433e3d783c334f028592123e22ca7395ee87912ecb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha79f5ad3f73cf01a9b6ef8ac7e2db57323d036f8fc3a3e5d4db0b5969d2b6b97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91d7a4c4b4d43e5cc713dfaf371fc509784e26cc8e788283811ffe087d7bce54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36e397dbda8898bdafa311e9e3c9f5143a7a93337d0505eedfb12ab915f04811;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd91c370250402d77e1f1a016b94059264bd4bb6990b0449eb0a65e8ad65c9462;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e4a297c977d99fe5f8532aa881741b5cb211e176f5ec78b092b54cd11a1db0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8efba9eb8513c02bf9283ddbead8b221fd9936a56acc30ebd8babb0692afa10f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1be6eb9bf90f7469e3be9da464f571ddf8ddb4c7900721bbfc5afa33a02f9f35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc75f5b92406fd123c4b21d7881c3432d4c41ab2d7b387479d67fef33c3e61628;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf08ea3d91ee3d0dcce79189b8b346858c1af66c5b187369e875dcf5b0f63da66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h928ff4af789518c97abd7a3f63bfbae0219ce38a5b0187b270b8e613e822f273;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed89d9e31167c1913840cb179ed77d33a7fb5b22bd8f62f152521c85f7a0308b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9177224a21aa56dbbc6d5c097b61ca48f6f2afd9e41f145379d427097dc1281f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd51c4c64ada367d223edd22af0d43929e780de263ca751a67a9e4ed8282fafe8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd8a4382b95dd2762148d5b80172812fb937d5bedbc9fdb1202417423397a09f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc7f15525f9fd76d974afc677527cd7797ac361b1e8d6a4b34837b850bdff3a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf36631be449a802ad1c8f6fee0ae9c455099e13b170e707705cb6a67945b3176;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5279bb507f8560c08b18281c49bd12edf282da8ef82ceea9c96194d7e07233bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1f3e29296c13ff0e1b2a9800254624382e7c68125e31a535aa2ab937bd5f62c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d7a855e57833d19803d8368166cab7ef9e4a59d2109edd773882ee193e83c89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0bd645ea7e10058835b2703269704f31ed67d0c3467475c6a7366c111642c42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h366c203883d0aa48186ff8f46cccdbe3807baff575d02936505f61ee3d59b310;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19d38676cd521631c3d0dedfe88bf8f1e929316f53fc9f88bd23dc91784b9931;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7a47cef781eb44cc9e7a30f31ee5ff0ef9e316d84092fa2deebcaadd71e4857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6be6069a7c479a261a79c2f5c0513f3b85866402c6664aa00bfa96cd03c2dd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c579cf807d3ea4f82375817557d2cd4ff9394a01e89af0de30800eeddc9a1ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fcbc7fe9041acde7173e24e5ffbe4508f27882de92db24e136d84fcecbaa826;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf222171361479da3bc2789d4ffef55a74e17e442023d52d966aed94de9a2e431;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha29403ef276424883d39118049b2f3440644ca7019763822fdb612d73dc6501;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1293cf0c7cc594e3e20a2880b40a9b6551478d773ebcfe6756dbf86b8e3bfaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6073aad1e1e2b2ac3065a520330d600bff36ce42cfb9708db7dffaf3cd89bcde;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bcffe94f8efaba548f75b98f858611efb9f50b93da3bcae640c5d5f4513a772;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h880821ab930844745beb4baa29dfc4e3fae8d7f93d6f3dc4df8940d1dd05541a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6127479bd64bee7a76ed0c2fbbfad932926f651183adbee2634cb0c10eff683d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed26bf612c163044853f7e670b3a4df7f937fdd0711d5dd9cdf96327d6ed9903;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a20c86e360c104426174bf44b75d06ee33f76e2fa12e33a71e12e270ee03f76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6750e16cc2a96e308fb321b435d74512f452f0a2680183789cc9c0ae86b2c2e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h886757f18e2217e2e821b4efaa6278499a1b31c7025e8e0edca6dfe049bf7598;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5a4b2161fdd96ccc9a14f8177ce61d370c8823b769cd4676396344db65e563b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb9693f61a4ad0b2c06d62002ac9168eb71efdbe0045cbe4006fd4703b40d425;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60c7176d353bfdb2e3419e1aca9b67b221f63938acacfc20e3994fbad2350987;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea19c38c79528542d15f4fff80701a82c869af896e98380e92aa9dde0346d648;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0669587d8f805e88e47583838149e1aa68e1c44b9288e62e68980590e07ec14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc269aa5692ffa11e7ac15272d807e64a43e026a3865959849512f6fa110d05e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a94514955010410488565c098646f75b957f73876ce51c8dae923aafe98426a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h399a676b995ddf6175f20bb6c366bb2d4b2e2ec35c93d543231d43c68c9720cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd211f8e8fe403a22dd2dedb993b22e5ccd43801380457b3db2fd23b7979fe0c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha00b82bccf4ff6b36ff5a29eb7eaa34e09ce57bcb35dc6047f37064964f8d5e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d130b6e48a72c10b37131cffa1156f67a8dc67b90dc0cb1de82e0d74a72af6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdecf6ac1ce0a6aa5a3e2472169aa7f173367c662e427861a411cdbc0811d2c27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfe55c65c24c87a8818f14d97fd357d2e6870c30193a76939626fabaa8015dbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94435a72baea28efde2c1b8614902bd6d3c23fe4a88f2cddf5f5d87e997719b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he759c2fd150fa793b24f7905fd8fd39356ff9ea71b307d591c043852aa4f972b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbba40000db050136bfcfd42f9fc3c936b06bb1661daf1103331b8e62b21fc72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ef2c636583a70179a1e01073a3315c1429099d5ef0847b2e0f1418f87b15d87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1da7ba2442597971947fddd298aa629529e90f0e56f1afe3958d945e7da51c54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86b46e324eb0ca7929859752459e1b78d999401eee1fc70f380d7b3f88921592;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39e3c651d8564f87228ef988428832a87e874873e62c47b2acf7fcb04383009b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb38757a47a75b2207bb8b4cdf7c6428b37e8581fa273311dbbcbce4dd45904a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfaf55976e2541030efc27125f98e168290e95e004a2e42e38e96f0d3111449cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0efb46d7bff60a2daa9e670f58d12369c10c1a9844289a9a0755b61cc521a65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a808d180d7cfe99d32bcfda65744631a963ecc939550bb40ba1c2241f0c7b06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f7e06dd13659f8dcf3859b2ad47562dffbe2b5e322134a69554fd6739b9889f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e8737850dea7d7cc86e0eb5ed3b6d503da5a91a724514eda57faa715a68aee9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96732be129bebde3c978d6b0e2aca94698bc7b173d053d6f86a563cf1767c61d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he297100104707bb9a238bfa12b803c94a5b576b47b4e856d1835d52c86beacc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89d29e04fc6c62ded8edde570e01fd9c17df51232c301724d91747234888530f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8de8aefb2910fc3a1a27e0bbefbecb886708d0b2b67d0919d070a4bc9d218481;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5288f50cc45b8a75424a33c0b14bec89a0f0dd35abc60df6ebe32c6fbf254760;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha52077b237550bf9197d226ecec0b6ff78297a51343796f27e627bd3a061196b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f0d70f0660b63a6e1e48bff6d820e622371ba858a94083b5ddde937f8e1c4c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h328b94c50e33c562a76344df8f69935fe3d027d8c6020202d8777f3106f541fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dc7ef57c88a63405d1eca557686a0398ee02c50338c1a1937e839b6f89a7919;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4740df4fd4d60b8f366194a280e2351e1b3a4d04a5d844ef09a0d4a1bb4541c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h301e01f54e540940909a97457ae53868934edbc391f2b981c318d808121f6b26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4006b2f7665d4c77dd14a54503586cbc72b3ef5307eeff571598d098aff65bd1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd149ac603f6fd731d9f66983044d3090f7587ac28648c6b2a11d513b7f0f940;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcf398f58ceb53364bb2b4f2a3f6fbc39d69c16fc83c2ca1965b113865ca6afe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7be0bb25762656a0ab2e03eaf2eedbb1303448467b6b785ae0ea33e2e643dedb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha815218c1dd116e230b5311b3099ce021fce983bf44f7772054488125a5efb5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73b5fa429d663ab8e4727a65829ea8bcc21d74d4b281352cdabd229b42367e53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cdbc9f093a35cb58056962fba7a518dd27e777c2c2e0461d9eef002be09cb4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0876eab74cdfa14df8a81c2cd06df7620dd0fef0062ebe79d50032546b49245;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h322a8b6f86c0a8f5a5fd36106255d3c680d41d932c2bf586c0800a866812dded;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ef87b79545ca7493ea3c0b73f4123bae8fa9c6ec53983eaa4ed50d130fec76f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8752f4f72ae2e8e80181c20c8a99b962528b12caa342a588559f06010b1b82c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e8bd229b8851b512ccaa668bb19bdeb57e21cd80c08f05efc683f08cb5e1f3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d11aa02dc6e7088a8d5994073cb89e8c202773fb8216d1a4458a0a48ea26b0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h775db3630c05166115ac0096b2540724c44d85edb5d69e5c82b9e9da2ffd4e38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9726a6316344b414061f3582bf887fe14670039bcf029ab0ff4301e3a0504a63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5d93f6567e910abfcb249edccec4cc66c264956bfdc238019947e0d52ef8e54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha23a0732d1a79a7638f11fb2977d93827c762c3adae5fbfd64e6585af39d350a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha18dd049da95e50433f699159e5f7eaa5f39e1428adcaece1dcc603b5a0a8bef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6596e7d5626cbe83e264d45a28bc504734abf6e2edf583755440d2d561b5866;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he81079cab3ee2433874c849560deffa9cbb8d50118607da3f48f74eb3c41cc52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf849f6c00646d739897f25f7a3464176bc784168eb324e46deb197811480de56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2f5cb8829bbff7decd02cf9fab6bc3d585b5bc727d17169b40b84b79507e95b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf09c42a00687a6c0a475063aa92e375fff0d96e12c69cb842f7138811e755455;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb04c390799554678b5b9ca801f84075cd8d82ccd66156a0311a0ece4b6570d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb237eb001e820f381e4e094cb3193daf2419468f330907725552266c4e9db9bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4c085eb57fb66ea7a949f58441005168c5c952057fdf6c439c9ad3a011c8a5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e396aac09f19a7701fd3a08117f922d6363efdcd0ca7f2ca6ecbba4a15bd455;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha428f7bfa1a77968f38a5ea7a87cd6884b51946c35213732ec74b4730ac56fa8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd69ae5c6dc047fde9254f9e38a84e8d0662b3c9734425ecdd4874c34e54e304;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbce1c7f397f4210b94070e959d5347209beb0ebd002fd953735a70e13e29200e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fc03f77c38b97c5b48626eb11c6c6aa8dceeda9e5d55d4ea105280a6012f488;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9619e3dc46640febd20278be730e2ff30c869c3ce6f38b1623d0e32db307d85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c0c7ea666306e71b960613e1412925aea44ff613c5419d45d3f7ed669b4558b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd85d40cd4278031e93b5fdb1c6a639bf79d336fdb7db9eba3f66b6743ac432f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49f8fe27581550dc0caff83ab21f77ffb81c0d10d83931addcdc631ca8c7fa1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20475cc800242c3f812e3425e6fc67b619f5bc7ff8f12fe421e6afc97a9b7b1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a9a6a6d1f4dfa80a5ba3effb06e972bf278b97ccf59495a702049a5405f42d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e9018a5b81598c2a06c4d6d9500739adc01f7cf67dd2457730c4d7e07df8a05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e17f9679ac8d6516b129b7caf4dee68943d9ca1e3b63bb2ef784855c5876d0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a6d3c7372d4c0aae98abc62fbc2a573cd422db93eb2f34a3579e86f34849c35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h173ecd3245ee2bdc52d806beb5164d61e0d7594b64e9777d52ea28fd81bde8bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h588d3be5112e8c2dc701f32a4c158264b315a1da209d00053dc8f2c4b16b8889;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d708d4bef546ee6de98fe2f0b2d839d046648d8472db9a458df0cf33c4be902;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b34a86f222b808afad3e191391db467db7db6578288c93d320a2eb24bc56c77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd98ff73de648c39bf8ed743f1ed50deb1980460e0dca342d9a5e615e4e9e823d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe036493cb44b472e395820db1c1ba27a4ed81aa8a0d2f6a50ed29bdcacf87d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fcd156838cf8fd9f29d373920cc01b9f3cfcbe2d2a91ed6fed5aa40adc7a341;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cd0b8607b24bce5a354c01b3dc4847737e5f163d0489b0baaa8275ca229fe6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1dfd10b04d746555788ebccca3e0c3c5908bab26b5e8716b7f02126be93c3706;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c12ff1025774c4f48108c40f101179def4131dfdcca2e2d5a936d9f3f53bade;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10a0040990b63fb83050f3f06ceaa0c75c72708264df3b5edbd3c8729647d536;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7b561a444590ff75b0dbb8e23603d5e4202f512b67cb9d5a360ae60259663e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76799dd84934281ed4415b63d7d3cd89293074f22688c481e7ba5f98dcaab876;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a7d14aef17f25f047500aceb6178fbcdfe90750c221682ad61322e033fc27a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9344fcb68a6087fbc172792e6ad5c33c5965c43154b9ce9089101ddeb4a5018;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3b5204b77a303edd656408a25ea68d5ed7a30a4beec175b83529e4eb35cbd50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ef9609ad424ca5df6d4ef8e3ee5525a9f8a5a00e8d20ebc320ba15acc264c2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6b5a1c3927f388edd0d5d1a7f8459a34fb380c18251d566712214abe96c15be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h404b251565913f32b57e7766c5d28593cbf043a9292588e9a8a6c2ed67765fc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f586903b666567d2ee91aaadbc6210abeac71cc0192f488e22d344b83c93c72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb24d9afa1d16281c7ccca04c6bb1484a6a8b4ebfa5c8c00cc0e3799bcfd5d4f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he594c30431c7a2ca7d44d1067efa597fc512bc67f696ef81ec48c7391d711e00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90ae60a9546474b7438d0f7bda5a4be663224ca842a362b0aa76a7d23c849c32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b8d785d837080c0b92256245589737341a30b72cd90d18f9f2e1de01c7e5268;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a668ccf832e99c6fde5372c2865487fded8a5ff3197f74a0baab08bd334c083;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24631ae7a85f6ac4c49cc822c92ea7fb136f068796aa44872d36af45ffecc7cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a536b55248a416dac4c29fe5caf51cdb62146f2c9f88f62f87731d72a503165;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa3de47d36e1aed88f26a892d4dca08073288db0e6664723e3faf47dcbbf336d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41b7a87bda07cec9f1e34454fe27e0b12e0a94c166b0308291eace6a782bb0e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf9ced42a1db492d52cd40310a334caa3af2913b3d57992663eb1a06626030d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h388aee69f8a1406b28a98ad88a6683a0b515a01ff4d8171bab3ee6f25707eed5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61860540d995daf653b1986d419c88c4e3294e1e998b7cf406d584bebe99ac82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4aa9eed5759242c34088530bbf5a815b707bcb6534b2e7a1c967106a1e904535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17ec38adf4873b08d0b4f54c90313f228477df4341c4efd072b261e0f27d73a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcebb1516ab79e12f26275e95ec862a0779c0fe204e0c10554396e70ee39d37b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbec1610fa82745d2723ab91fc0542a113942bbe94245ab5ee249f94619900fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcef55adf82f3e9789a9c7b08483b26d3db9aac667b93a2da146f4843e2c67e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda43cbd7b26be5838b3ae2aa544d661293fa11157fb70a7a9723df3e4c16ac02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2310027fc640d4844e49c69ffb5a5fd63fed5175e20936c0d6e3215c4db8651;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f3235e7a69b198728b2fd8e9f8012c6c12af3e099847e3eca0f8d095a434218;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ddbd69cc85b4f6dfc6131054533cc56f198304254aa5b48915bac66d5ad1801;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h236201c74d05e5dc23635ce0355152dbb69cbb440bdb54aab9ecab2ab118ddc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h824241fc6c3de465e12f2439921d57fc2bb8929c877749eea20b62be9003c03b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc605366b35a4802d3a4d09c93baee87b15525102a047e4790dabdd51b9e25083;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda764bfc7f4dd2c824c0ebb2d463fdd3a7bf267b9b276cae433f8730384beab8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb484bec75dad77b7d85e95345c4799a65b1609014afc79697b3e4ccee6f74f97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h640d225352ee7c5fa9f9b55af1489ccf62192cb854d26e8b41cad76adb42a962;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he10a2eaa3c4a13cc38faab17706872e90216c58bd1c6c09d71db1d5caa6c2930;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bb935d91d9c30a557853684a10d568950f29be8514a48a487d66eff85e605ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h669fa63d36a5abe0d663852c4869b7bb7d332b49b73919790697229e6d874258;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a5d244969d7e0d43bdd02614d8b93b97a0bf8880f68dfcc3b938eca92eddb02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h401261eabb14d238e7b14529161a31ef7bb0ecfdccfb50bc6bbe0d582272809b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6ed96b5fe7735886ecbd756ff4040b32e6f62db3f9b6c2bfd05b7ffcd57b423;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dde1a6f534fc7b1217bae7835f64fba0ced693d09c456c8a3b8928c336aba3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbd5dbe2f7b113efb3867c3c57d5e7e9562fd561f744f5149f0c140b8f316fb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65fb5d918cac129a0945fb653f6b3ef88b3260a960facd76934cdd08e956c164;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee047799f0c02841a4a4c6dd6a416a83f1009a6e1d567fb9952930396b728600;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h149f9163c5dc8dd6d6e6e48ac38c029bd7fc525402d43616c1125cfd586da2f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77215b132499a6108bbfac33f89196e8c53ea5289d2869f273630699145ac207;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7750ca475e28c8ac7396c5afc01a8647379ddb4dc7beaae1c5c23a91b4349e55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d474b1f31772b48dc32284ab9ce3e762f107f34cbb1220b8baa45557a16f903;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb706cbd848790dd66d4fbc5f02fc1a5516b3f1726cf9add151a5ab8b302946f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3440aae019165edf95a498e5739da73e4d7754e188ccb73601425cb9fff7b9c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he95c5732b0c802ca6106baabae631a1d6bf0d028d353d1fb92e0f9087826a812;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc0b9d66a05788a5e2c9acbe568005907bdcaccbfa317e847b9786bb27d66904;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e98c65aeadb0b169885b599187da2fd762304a2e0f74ae8c87a013398e6fe2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb5b19418a51cb1388a5b524ce912a43c36cbfcffdfeb5e88d5bd2b5706a0a47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc160486f57f766f0637a905d7f256497562a41952fe6f4142d014be44a53ec79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72cf3adcc21b1d7694a5923dba284e97d7e1b5a76add4923b0b88a9f57d13d2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9e0f42080fc73caf89279b4cb75e0a62c90a6cb576e5fcac4a61be76af3692e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1b72eeebdc33593dbe9a533dc92d6974ed108806095646070edd18324acedda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8de9a16d50e34bef8ea72b9fc768c6580d2e14d85678ac0acc7cab9a7c10fa9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc60ddb5ff59978c0d8fb7be7bcc2f5e5da555fd1fcf2139558b51d9faa98f360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8c2bdb63b915ce5d65b30aa36c8c1ec5d90dbb219387a0de460ae4183f9394c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f981e2a51deb4dff536a4c34bde0a04b89a7f34a6c2dc99f96becdeef4c1f7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h974b0de193d6dfa1dbaca29c1050428f45dae066aead673ba604d52b2413eb42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb06cb96c1cd785df963bd498efdf42618e19b4608601825348bba3e1779f64b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h536aeea63048a7ff2f52c9987d26c7dc78473faf148d8883b5ea11bd93f6d4b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had6b800ced1d520f20475701468eef021b1998ff09585243a7fafd267b475f94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec47016bc43c567c82d5ff03d112edf9a7baaf3d5fcab70b2734c8882196136;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2adf6d2ee966be2154bfeb277aff3cd91288158d90b348287d5c358ff66415e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e2768777636969d20254f583f64722ebfb6712dbcb83881009d1091fef01606;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40a51e383413f61dee63f8187b70912ed6cf87d27abb16532a8bfba2487215f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he78e755112768f1e72cd68db1cafd0c353b6bcf5b8fd1ccd797e3717a36de889;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5936a487f9d6a3d72607ca65d497e8af15a607b3ebb689a376e551ac9479b06e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h703ec259d1cbf6e888ac05554c424464b09e6cb09c96e501c817c9056649438f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cc89f341b787af73eadce335fe8de23ae94714b3b360b3bcb856faf1d89fe10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h509ac9b034222c4a9d6d83c2066ea064cac45b0d4b0f4e172355079cd2c39b93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94f6c674a4a3df10df1c134875a7f262ae3e73ab85d72ecef42229bb6e7358d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc47bc6c99d5a8ded57a2ab95a9464374881e5f44dcadaa98d308044fb67fd3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61ba2c89a472e627727848ea20de501730c40235b011782b14a5fd930f13028d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefb03246ddff57cba8c4d65d4445b87fdf585c2e16f464f9b39cb91437881bbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35ffdfdba98920e17a036fb71a8aa9df3251dded36a62659163a40aa98d69ce0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h272fc134acfbd78c328664c2f5dcdf1a7d0c06dd774b64afa66b7d22724470b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52746b045e73bbdad4b6722adb62120df48f96f71b1ebed66d70614682803a87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba87228faaff9926dee60b05d752ba1c845840d078f2a4032eb6895c640d48fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf19fc58b784dd9f4bac8623649334d0496870d04410d3dcd57ffaf4bc68ebdd1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc812d58cfd7265a3fd489dcfb1728af9e5e8c72d90c865d2f303436ad76acec5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he316d6a376aeb6f47585e5ab200a967ccc31a9115b476e68837816ddc2d1bd66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h554201c119423464fdad4b2871e9eafa8aa2dfe81a6e0eebb9b78a2a73b9fdfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8dd25f9b5528e8455ec4f530e7816c199b11372769d5dfe57b064d3c89cccaf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h348c873a430ac6f62296a7eb6fa7e3123fda730899731c5382b37c92c841b745;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63a9fe6907d4454f68d5f7e317dad7e797d51996a0c66403531092e516fb17ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h244c16484cc3381ac3df19a1a14acb5f9c32790f2ee832129155132f431cabcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36a867b6a3f4d7cb8df107171762a0ccc181e4a4d96907e2b34ac94570ede619;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h116a5cb30b4fa4d65dba9edf8118884bc18b35d3332eefa038d8fd7cc369d03d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30d84a35c0e2dde8a051cbf00ba9268920a0c4978aab5364a0ceed74d71e6045;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96d110e6f24b7650e546ead12a529d999e29a30772698d93688a694413b63294;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1484f92f77b95c6aacf38ffffd3fe6c14a6e640e4a815921ddaa30447c0d5cc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa4014d42183c0f328fa919c21d025b4cff04751b96974667b9c27c37f3f094d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16cf9bb830f5eee7b2b89f1044b89da6e6923c3c579d185e17c2ea83bba657e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h732139c71ab1ddb2bb42f6a4451f2cdd1964d04b42f041930a3d3323c0e87082;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4030064b419f5c5d48f632d6ca9746922050529b8541a95d01516ed44baa621b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h615ebc8fab5e5f18595ff99c8e924d61c553503a0eb271df39ff5ba187814125;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he64c97cc0220aaae0e102f9f19917f8da72cba8fdf912197fa68d7b984e71b0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d8b14640e271ef49cec25f21644cf3b80df245694ba94cc18155c4940449e02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59af51b65bd6eff50745c7eb55bd298961d360cd9b6b480553f069847a63d226;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52c3d080d7ac05b5f4c79fc56ca95e975e95edd2e9bb84eeb499777185925b76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ab18a00b54ae0492d0e8e7ee9d7ea2d3defd6f6ac307ed4354f15e67352e7f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7a3e15f8575d3aa6f0ddf6a1d584e7908295462e6de809fdc75a1d2621a99e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4916a84acb8839e1bf47cb4196712b91f0de3af42dbc2143bfe3e41903452b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h832d0bd24d2ca714a612d0478402fd8f488efaca234d32992532d82751935e17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e307986eb1a663a981996eeee646471a48d244614b1545a72bb1560d4427db9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50e1463373c5bf1a5568b1d020ca4634b3af13a8c1e6be57b32b397ac762fa0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb2bb509e3c6a5a83317a8923f2a108eefa0c7e9926576ba4035f2a79cc84b40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cb47bc32a2f5d8731d09c31a5b0e7fcf04b4d318f552bc90a6c17a82deff057;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1bbbde2df589d1f786d5598c1ab3c7a121ed586ba7e2c75cbc0afd6a02b08780;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd689f5a7bee1147432e7d88663b282c54f8a02b7cd55d10f2f03feb638eaa75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h345e967c93571e65e7ec7b39c2097958d49a3165e63672c87e69960c820474de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1664d7f19538bc7b977593ff3fee448291016447f2b1d49a765fae986ebd2ecd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac082f12179501dae50ae6340aa89e706edfebb46754d624b9d6ab949275235b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa26e7e07bc07d19943cb0616eda0a5a9ee9d14653ca67a5deb4c73c257e9e76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h284fe54fe895a50d1a7c8c056b0a0fc6e0fc346d836450cb080ef40c38137643;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h196096030eff6efced4a087a81839e2d632b86ba6465b3b8456a2c372c838af7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea6a3f9a8ac088a94e9b5b6dfe085759b92fbe8ec2b02c714ce03dfa483cb026;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2636e7b04a83ecb0ad2361a585579301376a3adc75cfa1165084172dc778afef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f16818bb959c5906525aa5d5d2b1fe596f60670257d20959cc5e933a46e6b93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e07d253b31d896293d4935014801501b3030191a3126c314004dab5c0964cce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b1b636dbb3b73186dfbcbf8fa695cb66328b869f9a97620efcf893ef3e9a566;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h726ce64f81be1ee6d23d0be18473db2b84e1a5b90188289b49c520032bfd7e96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3f56cae8ba3efaef861a08481d77f976dc75c9d52d2289e9ea30932bb753c77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h351cd938a1042168d7e9a80745f67cdeb04e2b7717dd3e39779e2a32e3a9dacc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45f210a5f7115cbfd8c186fa9257a009dc41c922bfc54ec294fb40c50f35e916;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9ddc152f1d16b625e787c9de164b78c454cdf187528490b7f8e6f1e4c59f382;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65c5afa938cb8ee7d7581d2194f37efd752a6d8592241793c3c22413851660f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43310156e280372fcfd579ed53227d99c7bdcd6d33a505c200d5e5cf25d75857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fb1bb7821a53da4ded2864159b78155a868013a25875ca5b11f9c5e671bdbc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6da5294f85cc7c80a22bb175c0d160057d11561aa9de90432324f0eb0114053c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea6661343bb35155be285b6a20a81b1559008325e179506b576fdc59a2eb483b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc814267335478f565b9d308c58814aab13b8648fc460402ac091df470b53475;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4c8e0d253c02fb8662c475a576321e78f53f7d4d0bc925e86b07fb820a43f61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe908fe91dd5c84ca11622b5eaf20082519e78bf3e41e35648cce3d7d1c8d234;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50e7f2bc968b3f82a24fde7a5201adcd756e8dee9cc2f18fac7a9ebdaab247a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b48fdbc38d71b46414090184618412b4ea340a3f7a2b65a3734d30a0f6336d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bcad27033f4de15b1d271675d8b34539c6696298e5e20b16e09e674bed88cbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf742b8702cde2f0a9550f7dda74e78c3e092ec41f6cbd823c6e06d6d6f1008b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a50f8f99e03762e7e37b8f1a04f37a52b1b3eae6330aff08feb4d8f7ff79e94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a339ddb9136389ec09a4546edfdef6a65d2a5f1ae21c336ebd3035336d59140;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce493485310ef9e14f13daec9b01e2d0ea2d43749bf047b1c9b617f83be81b4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h653a0f292a056cd1c277b466ba308554847475c1c78041f4a1bfa3f7ffb7b5d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8045a405ea6356246aecd3858a135fd56fce9d678849a14380e22e29ad2f6564;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f2f57247d790831df7f94be3ca1802fed8c120fc6b2f2f82945f3bffeb82351;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90d71ec207ded600d4c9559e2fb6a6143709c8966e2fec29b7d5b4b5357b318e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he838159ac1c1fdefb68be96fe1e6492d7aa08194ca67fd6834d0a4cb808756af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h832dc95c088f6a903056af8cbc2fc5ed4c706164f51213af8babacd96dab491d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2ea6eee6534a63be236ea99cefb0b3fec59d57c439496bd5ae3afce192cecac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12d5d0fb2ea37e72ef9b0d30469100489f8945c662ecf42b5406817dbba714f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12ab93c5da4a2710b2ef901ba8eab650a89a3fed30df419ce717c3f2ee22a7c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4c02f442c746663e2710acfae8c94072004479a6d59e8d3bc094da9b15451eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd3ac11689bb408b4fabf546e328af07ca1d62b72cee117fbcbcaf3c53bbe1f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7de546ac116ca8b850ef5c971abb24f4267d22296ae70f5e71c5650e7cc98a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb04767953317648c4cd2c9c1741c020aea53f80e84eb09216d4ade47783918ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8f1ea07c052e78e84b20acd0d0161f7248f7e208c1c3d90be961ea42cedda31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc86276ddfb535d2a69fb07eed66435418ba2ae297ea6bc6d3e3d2ac26f21ec01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd97acbc82a4c6bf9d93257fe876fb3dc91d278c9c76566075d7e610f63ffa7b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3432c0b23fd433cbfebb52624ef8d21f016c37f737d04b9fd67b1881a634e862;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h450b81bde5ada9295b1cea43921da7e369e79d1d915df0817d34e0491cd22cb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h703f8a32c53810d8319fceb0aeb6c6d85e37f0df484a63607be5ffdb19ca9c6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha86b11a9155ef9891308b9f31d98bdb25fd64c5bfd7dd398dd938d92a1876de4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h780194609adbda168f5c1213c26458652a1f6d46861fba53759aea77ec5e2cf0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d8bc1345ab7be8b8c46b01b90acf509509cd73cf8183f787ef950fcd14b01f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74c7a9f353de7197148520d8268dead45e663cf9dde4a479f249512f2934b33d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78863246c45055e2bd0969c26bfb733792effd6c5cfe0f3433f6715c79a39a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef5fa022343d359921de29ef762db97b7faa91e107f378a618d4fef3e1e246da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52a4614be56fc4068e60aec2ca65258c568848ded56adccbaec221d99e8dc349;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed23f469779c976c8ae8e741ebed85bb65c087fa9bbf5d860eb5b79db3c3059b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd73c67137813470925d2a1e7a13c822181d0711b8247f4927a6579f58f3924;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa4ba802e8aa1263c4aa7c3a32df3229ec769d2b35f23e782b0dafffc2b30fe9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfb4fc8907db89d88517090a2aab2949697f45fe9e6715f9d4a378d9ff473bd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d6b6138654f7541a550299ddfae5ca863c133b0c87f802a7230863aad0bcc2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70ade3fa5f16305d51113361261492f94ce7e30cd9764cb240297070b56975ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eac649328547d159575e87ff10f182c6ea91ac588abc0e0933416872593f02b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f560a761f069e62a94ee5b92fb710094ef8fe962a9948bed8922463eff90a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fdfa1bbaadb47216fbf88ffac5c6ec236b50d4a61786a9d24a42962c5186bd7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42b91ccc2240313f18d4099842fef9716515bdc7b2ccba2214ab243329a9d88d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ad2b301eb25192fcfc32ad2e52958f7fa33936ffbd9c56d0fb4318ea917512f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e52ef4898be0f900713412a63987841708c9b3d35865f887c3f1d8e61a4947;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59993e4162136e7dfc3d0c0d7089d79a06a542b1a332d9907a5064ba68be86f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a2dd6d556095bf0777ba79e27cfb354d668fdc5077500e146164638e60109fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf10cc42c4d2ecb9d8cd6e5fcd3c9e25d849326ff56cd400a88e20ba3d15e997;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7b5e0702061b1b29a62df18ea910c57ccecb597dc75b0213a64fa81ebbf951a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8775d1fdbdf37c57754a4e02553c4085c8e24c526fe7f17157c5685bd8eb0cd8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bbe9a57fd94366618f9b0ce2ca479a1568577141f611dfb1de43614f9b71a52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f067c67a8cfda4b19ab9ea2e9464057b9d74d6fa8256ff2398808c69d24dd1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h639ed6a72b28ddd202056a9d7d99f0e1479e32b6d3099f96fe12036630db506f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9b08c28aba3f5f42cfe19f9c6e6cae307d79979b0fb78cf61300cd75cf6d009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93778585ef4eb80a6c04716fac88f5636a6cba5187e599bbd982bc8346e2ae23;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47251d9728c4aeb9af273f2ad118dd720185587357b7d7d313b96846e7471aa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h508324a258e77e1c191d0f2f4446599fa0a2ee070bfc8054bd31c8d0cdc50fa2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ae28bb5b9ed35ead80a2204c51cbc5ee9eca8f38d17504b788b45a4fc4190d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc39db98db74f23f44c8ddb2ebcd9b03972a5c703c0fbe0edfe5b8d444a29b59b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4889f25e771dc46b1d82232548bcb60ee1f863552f8cdc7f9b768af9d83f371e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63f4c039c73a0d78dc8b43746edd2579d4fb146e8af1376e5316fb7b74c8a0ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d6659ab7a7bfe9d3dc280f77cb6a4869e0533dafbead84b1452ab3c6ba33ad9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b6b786d0532db6d2e1647f8b09f60c3e1f1be50ee1e8a3db61681e6ed97a4d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc73758fbdf041ebe8c6f44aaf6434a7f90385dc6ad4a793f4ef32f28dca42cc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66ec39c138edb69422df8c0db0ed43242523b5421c70df8c9fe085b31059819;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2470d4ab6525cb5fb98a5bfda7573222c70d23bea8a5c74949e8ab073ebed9fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cc718e0a30e8962ac80e6c6da9ca67881cff7f893e5f08c9e106b309afb3988;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h216409e53c7647e3fa7368ce0692c3670c7888274c37451f061c699fe8424ef0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f75102376ea2cf3abd6d75c6fbc26ce14e865e8c54daba2110f6d734bbe45f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h996e8a9ef4a6789c5eb1b897df2ca246d4ed32c70d521aec658bf1093cccd677;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a38c300880d8e56816fbde92a3d3ceb3df6030e043b8841b2a9107cee11e7e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cb01226787cd52e19f77f33a107f6d46741920b7638ee61eee86331b7d75f53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd781248b999f75c0b5b38bc668be5099384cab0867e879dc0000e36cc662a2c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0cbc46b68499724df1ebf4e98d45d3793fbe45ae183e518cd9faaf5a30ce6cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36cb6761249f7d28f4bd418ccb797f038628ac2b46b2e00eb18750702393deed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ea893edf77cfe8fe4b743054d43bf8f6b0b01c42b0e87210aee43609a008d04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e6e02bdc6b5c320f311a35f83424150fd5ff4239d9b666553ae46a64c3fccc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6915f3d73086f4b80b8502929d8fb7a256b459e8485970006e3c00685563af66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6074201707b49b4eaaad39b424453d8ae655c0cb129c0ed2f48a930bfff8101e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88a75836935cdb331630803a728d1920ff1e22bcf88039401cf9561f22a22268;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffde2b1084de383470892e2533c1f52baf6353fb713b781641a2ad5ba42bf096;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63b9f28cf08c04292f5fcf165fbfa29aa57ae58dd6b44f3febc9eadfd18e4d20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2955217fc082d36f282510aa9da68198e1260aac503b7f73b6118772035734e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafc91ea11654bcdd19552d9394d5ac771ab63967fb09921e3824da18f93cec4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a785d735dc0ddafeba956f075fa5c38fd11a83971c64e1f4999a7313a2dfa5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60775a60651d49a6094c4c2b872ce1efd81d6e073bcb8456583628653c50227e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c5ab3bc56ba8e1a2db4404ceb38b9955ae7feada54fe7ce849c182bb03050a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85941cd04db12cfb623b65de3f4239b8ef4ddf5b21dd18fc97f60d71b11ea575;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f9cf22977dc05bf2f3f7bca53b79c76676ca6b84b7893f3f7653a62df74a3ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fed9276641e4b4542552dd48b251f45556f80fc07892daedd77e3e7aa3a007f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf054ec35992e91604143d1ba3584e31c3af3e1f9f7391663a99f4c0af5dae2d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h608b193bb50954b7419de530b0e74acfadbd85b9117774355d6295e02e3f70f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37d2ed753490d1d7bd312e7796b0dd99c54c76a18af560239d293bcd2282dd85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3c42fd64ee2c75ec618ab3eb3e079170a25308890645bd81c2a075aab5d70de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h285f219ed040be2cf14597bbededd1fb819020ebf9645a39faf4c298ec958352;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3d65d1451e4acbb72951088b73f8eea3b70556e2908c949d6fb691e2146224e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb044e12d92e84141dc5d645aed95dd2b20cb9b987702ee2afbacc74cec744727;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde9fb78d710f538c001e908fd7e411c946ba30fca1d7bf5e33a3684f2b9f8d0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h320b3c7e3dd96f0032015295ec62503aae89e2e64b9b817a2ce675d895b060e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f045f2268559cc8a8e6aa43ae50f268ef7bea03d445351105c4d01bb2a024cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf658ee6d4b37912156c746d156ca29e056392f14f17d611d25ba96a1de195211;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d8ba73194d54a087034d41174974c060f2e62b10b441e3a761f71dba7d30e87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9524c1c3a3bad01b7a89e757c84302e4c4d012675a948407e10d40b7d7069a82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7ba422d29509456ad4a50718aeb075d15d5d941ac16c36f0ca44f7e11de9959;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde94590f3a3df2de63628558e0af74130c1bb62294590c04a2ed78a0079c385a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5675e37314eba18ef87928c8142fae180bb96024ab25fb5bbce2350a360441e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4434a5b3a6659727d0271558778066077cca093c1a8bd52e808e97f2464ecb22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8b5c98e801fe55c56f2bc24e2b77e696404abbbb94b44bf3c5f8298198ed90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c52bb37bc8d1f81d878c745769f8b8a7e5c2f5d88ce7111469f18014f46481d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb6a4f89e22be32cd883057882c73f001dfee80337b87c7052ab4ae3a51d0d99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h512eb07cb982cbff5f32c887348f13a5440bda06d2932a73a8933e47f2ab6f11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd16c4aac58d4d3cb80c342418a24629061c47618aaa8c23787c92ca0d61138f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9055e63834f24c6f8f4dd01b419d2ad0b5ab1aec623acf54b2485ef4555bb116;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc790aacd09c4677b45b846c3634b2fae307950922a480e3f1c6f5d828965205;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h135a174e35ca7ab37def6e925bcf00154ecb9a16bc0e258a195bc3e521674ea8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5100e95ef46dd23da0e1abf05e644ce1ed56141dc039a7f4e11eff1295e0b905;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9a3d2ac1e096e909de837cd7d6d9579d096eec736ef64b20d81ce630d3c422a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cfb0f1fcf99bd9ac98ced621ae95c8044b4a72dfe1961ff427ef7f4b607015f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had74c916d8ae6a679009beb21c5ada912c29347faf4e154b0ab6801429cab6ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdbadf86bbb9434ce846b7c7e8a821b60d9464e2d169de82cf510f506d94fc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9fe38921e0e9c3267b3b0ccc08526a1ad65b7434824b28349f9633ff6e3c70b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9e567b2c7cb0c4b6dca17cb915ba25ee851fca3f5ec4a25a834a67fe06c2a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he72470347a7b645bf01fd3b70aad30cf4addf5acea9a4e92bd510258fbf8ec52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h994b3b920f5fca5f97cb754146d2582194541e54de448a7192dcbc511b896c9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h272ee9610031c8f72dad122b7c8a5c39904cd07fb65da37c3d11ed205718d6f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4cc7c2d621933529fbdaf34c62c99cd6859eaf874a4dfedff6de9c197540731;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57111c3015ef546801ca6a28ea2db4d1bbe95d944d19a9c98450d43e48d8d77c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h801754815b16e64715901a5fc4413cc2ec8a1e1ae9e641e42373b2edfab7ebca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc57e57edc2f2b1aa76b807571167a906a6c75b1e44ddbe87f4abbf823216da0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcbc77d20bb04550d701e31deb11b482b83bb177be18bfec438bc312977cec58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb39610366dd954f206635c154aa0967c99cb2cab3eb3e2f8737befae3a26408d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9b4a4f85dcd2ed356582430ea5f8e197d810b3c5ad09ea25ef53e3b8fd4d2cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac6df3f5d25041de5edefa4c1d2a1988838118dc2a4b08c67ff6e91c1541025d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h122e46dd3ae9319a9b9cb8c70f90e940a7ac4b0894a6ab0ca7823e86ffa316b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc9e877130ca52c0c2c2ce006990a5a90dac43c51feb7ae1966f4cb3d469fccf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e68fb1093df4117f2f75a7d7f7490b375092ceaf2dd6d6a1d865abad8c6a04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eb8bb9c05b69fa45bef8b5debba0fba4a02852979771470a8b66529dfe6ede3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82900f28d97f430615255f551fd58f99621117dab5a6865da5a6a7e8b62e51d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he85b1fcc99654fafa12a43319aea5c47817fc0942cd37774343408b4b0b5b84f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44f9b52cb38e30f5dee411ba0e9cf51779149d743616c57a38b58af8178cf2de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4714d31b8c954994a803d8b9dff85f0e62fbf46a8fe03be8bea34bd37a0dbac6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha219cffa4b3d2df3ed007bf7e843f7f57448c14aa0cd80ac0d68eb42780fa2ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3d51ee04b0a7da9b83d2fa9fbab41c038a3128f38c7ec25562ecf513c5873ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h716bb1825d976a6f893e9d586092cc4e42c4811d3fddd9f67490941fd389d476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41b0cae3b95e15536af85a37dfd611bea389f453956566ffdcf11075b7f0583c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e732caffae53cf8c5e398a99cc96693500eebb8dca47cb1c0bbd545b698b8a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc71d183d261f64a013d18b8b9aab1a455087bbc8349a94c807338e50050836c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h897dec0270a9ace89ae650021726e60a6f01354751ec997cde7c2cfde73d98c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c6ffea4b8b3d2b42b016713b60096da32f885b171b41a4c0c8120ad0c5550ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dec500c656975229d3aa016c7cf0a1088bfc14230f3132f521eb40387e6ace6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haee9d6db3aeb5c4461e13f5e53e5375da7a15225ed8354fa126002ec47699dbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c34e86a5b4937c874b97d699c580c8fb952d4be16199c2c4ae27006a91ab82a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91325ddcb376b631652b15baedf2a1f813389bfd7a2e3da1309824b1d0f3c4a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68a1b7ca6302155cb04d109cb6343b71ac57a0c15f01d360899a495e6ed80041;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6465c1180c17232ed2a173ba2d03b36139114b95a95b372a3e57758af1134555;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h211dc5394fa78b0e23e6b0bad2f3d4d018508189adea78b3ea7fe1f962ddbcd1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4066c19c08642d5e459077c5b6158fe1b07f049cf138bb46c6cfa868f3e92799;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he96c942a0c825ca3716f14c8124d5cd6c4fdc550c34e9857a6d785086b64fda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bec62f43185dac9a026a6ab7fe377871839e74c60967b3c55c1e0f2c8dbae1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h387386891152e47d5ba28b93c588ecd029a251bbdad8b2bee8d18ab1f8dbdd1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf6497eac5f5b7c30701c9787e7e32cf0216518d280716d276aae642828b0288;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1528fb860351b0ca5e3f094180d0978c86a5095959dd10ccf5e6a2bdb131731;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f839790478de753da91ffbdd3b85090018f6890ea0f41d26e2a06babc02f565;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd08ff054b22fd661dd3a54586bd3c6417861b98f39e15a9ddbd214350a0e4d4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a8413eac6e9bd9c20e19d21646d8bad3a83b42ae65aab31cc1e51f4e07acdfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0fc6f8594e4b68e7c6b0980531c876ce63a1f785397467f6015439da99f7048;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h202211301bd37bdf929cd540bea82dce2239199ebc0a3154b4a55f3c670627a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa66f9af09b1d5538cdc3b1791718af9d2fecc407f83988cece52df3e34a2c38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he988756905841365d2bd41278ee175a8aabbff78a4e9cbc65a7803cc287991e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3bb16bb3dca6a655cc9558565b8c9c1c291d8f278ca6dcadcb56b78f9a0c194;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2c97e4c676d9cec2363908614ae1ca79dbe0bf2c8a1c5609820a3ef0155598a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd81ab9028a9b0dd8dfbed5f827c6eee0c2588a02cd8f468695898ad867e0e54e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed5f8bb70e3a618eddb8169143f1457ba65be91f154b0500857d4765b43080ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80c49e7a1cc1945ffe341df661d9cf6508009b6f4719c18b08a9ec459fef2ec4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72d740dbd5672f5a7956cd3b19de91f33e26a48bdb5b600ee6983267b3771a52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7c6ef6b36b1d181e84744c93a9968aaf96293735a9ff07352ce1063f2a47862;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd787a8902a752658479126cfa6918d3dac98674f98f580111dc1e7ea36ed9766;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc565758c2c90f1045798ee474fd16c9771ee072296dc97a13b939acd0fc2cc72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87d456e37050e04f77a8bfe81f15b5de99e3927ce229826c4cf6539d21c7e410;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf79b470cbe025e43684f060f8c9856db973ffdf1fbfa3bdb1d69afd4f1fcd81f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c065926e84a150e7fd81c8c974805b707b3e4b9155d03537fd10c2a6ff88ff4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2453f6b3e9df8715c3f44a4c28e335d54c102e9ddadf950915c8fe1d63aef69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6c31fb951e30d28dc069e57b9e6e114312cc485f32eaebc587cd75ec97e355d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6c34819dea0c775f9999f7ba6b474106870c5b9e522b847e24509207713e0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb87915ba798cb7622ea2f95550026b5861d5226b111592cd69e5d18c200d76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc34cc9a8cb03402119bc496f31dfc871e4b612148e15289259e80cc538d2f374;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfec515c31c9b30a6cb9e0f70e7c17b71aa52329ba9883e9f46e520aab1f91835;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h572409d36e4d99b6ce470645ef1ad5b50be20183a65d72d603d903d6602205a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74176ffe3328d0d57049f11fdf602d7b19276e5e467f4ea5255a75b3e7f361f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46d575937469814ef7cd430901cbad7d7f57272915c99acb00d707cbd3b31819;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc27320d12a45a15bed33e0cdf008dbdd97898a221d6fec7fd82028eb466ffb3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haad37045e7582501a678ff91ad3f74901f681ac74062cb04971fbd0225fcc03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdafd119b99082246229251a2db8cfb524c9cf91dd387c4e8bead8b37a8d2419;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4e5b6cf2d05a2c8f9268e220f4c59961b90e21a3863b3884a2d8411c094e335;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ad2a0f46a77465e841b6989dad7fa127ae038980e459b65eccc88012abcfefb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc36a2464e233cb681bf23803646283946892e116305ad51019e2725203593c7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha18134c4b49477965d42c3d7c2ddeba83f2577d9fc6fd929737a9ccca95e9e71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6054e8b312cad8d48d3baf274795ebea9e82934fca818c29cbce3b59d005c246;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98f01448df39d88ef3dee56b33f41d7e6df4d268b4a1099b802f766455293801;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab7fcee0165cac8a092602ad0e58e332fdb3de168758e24347590db7a9166f12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc32f4a42afddfb2bf6f1c7b55e892cf596ac9d55ebe3625eef70a3229fa64564;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68fe969aedc0e1b43f4ea652426f3c5fbd25507499290cc6596fd74b20d4e91e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha07693d58ea9f99f0bd1a8341bfd87873ee70a74c3073859740a7b79e4d1fe18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5570c5e7279f8ecd0f43cde659c9320eac44a63de5687092ce978606b720a77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3333e26d713b7a357c7582bf0650cea22ae434e2b747ebcb615cc08fe99d83e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cec3f628118a393be51206dc8a443e75911787ca534a9183e076107ffd282ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ad6b74477a9fb8ff786db89fc4438899a351556c3718b46d26f13c526c05d57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had26b248a221e3fd8d29992bb19a4aa1437f59c5e8f32a64b383850ce7ea535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h893805143b7a609ab5a86ee6d245da7abdc14b67c5e6564fcda5b0e86fe5cf16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46b1f3beb5ca24c267995e0ff22ccb607a6a336e62ee5c7a282b0b5333c7696b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1883030e59878cd3532729ad54ac5079c988c9c778910fdb77558a8d1d48ffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60186c7c48c21bd6861b3115e93d7f8baaa9f04527e489d4cb527ed1ca0ba804;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4db413a37fbaf52d55ad6238189b989baf9c7e5fbe4c0e00301d99ae86d72eeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc892f0eb7d7e4938e8292ff11d487fd6554e3e028fa5be13f8e8d7865e6828d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5a0b30019d223c07b8da3d54861ea1d2d367782ec960629b22ee3a2729fd047;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5697826370c12eb5425cac067ab702d8ae0b6f61cc2319fa56bb2284bb601926;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h210ccbb8c84cafaea6f525ef89589ac9b5513d675c93f42fb7f59309621e68cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31e62ecd0048a818b1047b2f643f46dc669f83b338d256d47d470eb9e476f269;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c13eef204b9225fd7174ff227e672b8748f836b312bbd1b3fda50ac3ebeb2b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90abc89ba167b9baa7a4bdac7d939d397253315f678b9a982554831974da561f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7dd79569dc5162301f84a79e22463583afc297e59136c034f660acab8314ce7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4afc9a855559612211cba00b806d795783b34169d04c0a8b27cde18c71c79e96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4e0cb35572422ed6c3f8917065769d72d6101a3e64eb226d1f46440132c5a43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb182a043e9560f66bb4935dce24bec27a97626d7caa16f641d13c7db89c59199;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd909e01e54d9840e2440ba292031b95bb5d11b48b2f03d480fbae55932b0740e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc62d8db7e7ffe60e2a648ef1780210d09c3064b654e9afb25ce9e930bf7dfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd63107a6759c310fa7e3450af4771b0f6dc913d72f7a3964e400053ebd254add;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73865b4496b691f87b3ff96e5c5d469a3ecc335d8e3b607d2f4f4ae955d66cf0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7923d4187ed7901ddb4c0a21e446cc7dcd64e6cecca7fc900ecd9767d501b932;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77d76a3ecd8685b951fa26c69e0324cc7296422511c4ecd143da496580652331;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bbf33e6726c4daf3dd4f1c6765979be46f45cf29884e6989a6e76279f775b3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5be44cf4bcc4aabad93b147c119130b1dd476632f43ba043613c189f31b4056c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec45002899f2c6bee1c7800d5a766c711fd521fd6cac80f1ca1f4878e397e10c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc81902e3899e13d26f899085b58dfaaaa42a38e8ef606f2d9e4564e027ddf5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b85a1d568224334efd06c37ec757a7388c26031b1d264d04f13fc629c5e2662;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bc6196213b34846ce7a67e4508ac9c09ad58b6a6a2b1e90dffc7ca4bbbacff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70839c3a985a0cd828753f1f605a6f76865b0520631b72defa8494e04f285092;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h792ca2f3cddc91179e9d4db1d5645140a1bc7bd2bbb05512350fe7465ecb607c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12033bf9576e0ec435ac11fe516cdc01254f5af56c5c2cba0d22ae4781892823;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42121c3ff76d6529b943eeb67472786452ac655ef031265cf16e7c48e9154620;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81b8e728fb08e89b6d7170789cff0fef49d3a705320656bed674e7d1621676cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdee64134e2f2c4cc1d456992ae875edfa51576cce6e526f722e731c7c40f0eda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb56d79b0b1b5e7e7c9458ad3673f10efe859d378f84c7a59db1d46be2e65237c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98600e9b10f416237d39ad9bffc6d4b50ff02db6127d11af91715d30feef3c0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ab9d75c1fb835c41709d3bb0f520549644609f3fbf150eea84f1373aaeb246;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h899cd1288faa20651586462181f1b3a398495d24230b1a880973e9e65ae282bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49d0d8ca6894602375bf2ec0391182f21979b57cfcb88690f859c00e3bd162fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5128dea496209e38d1a36096c62fe41f7108f61fd1431e0ff97760e3684c585;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61d3379a8bebc6ab0551ff50cf94efa82a85f927ae25bcbec878d43d5aebe8b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6a19daba688332781c39c214320681a57fb08bb80b41accad566338376e531f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99398397efb4d4244b293c1127a51a500fbfd283ff8146f5180e48752bca5ecc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64b46fee49a0db8f25a2f803d8357f05b457f8528af82bc2b286f31e1f4d0eb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f143c2f1c67bca724fbaa1b33845cf4b72a48e769222f3b55ee78f082c706aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0fec3e74c659cf7945ee6ecf31e5182d5c91a7878bb12200bd08341fdbad7ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h722899d235dad800a4bb6ddd2b81beda3c6ac1e0efab585913f51fc79267430e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf58121728524ed2784763a7170c059a8ea7cf78025f5a05b8329a1680e966d6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h776747444e04975779f3194c6d269bca1ff8d79e79e36a5eb362ea5c22c7691a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6864a2a2fa0f4ac8293e0c1608f26d27e3848decea9492995542212fdca4587f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24efc0b8e7297cdaff9a9dda654b7472ea52ab092f7533203a75338ab5f45d9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf4f4a52a0f809019662380dcd8eb2b48ff82f8931a4119cc3fbb74f865937af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb3858e68b9432d957f6519c83e1b17e001a60325b43cc0de12ec7be9e7045c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf58b8b626af8da30e47d60f86f34c138c59534d22797c022849406f37b08edb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ead8d0776c26cbff092149790dc21684c8db29aea728fe22512dd5d92efa1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8aca46999350da764cd366edec17ee87b96b4e7a5e67f833b5ac2b9a47b3cf6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b91a47e05b93acfa995b9aa919d77e2496fed4864debfeb85a5a5351f6df92f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49b70f94c7998ab54559dd498568167bbcde9ca020c386ec3e3fb3667e556f04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a318ebd6e0e58e6636dac965f4167f75d00bd6ce91628e9df6e5646b68545a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66839d88e0aae22f5c7ef5a9a63a503e4c04e73b75bc8d29ebfdc06c44bb2d67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea7797e98d69f883a78207a6b8f17284870d79b42b740f92b05b1267069bd008;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7478dac4321381675f365adab5f2e90c25ba544d28517b37f41f0a66e6a9eb8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e7522b014337f008a277f107d6b0f39416c28e621fedc696074b48cf8e17af3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca5d8a64f3b7d84a124fc25f9587ff633aba5c347af97b82d8b49602fe1042ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb84a57f3b85adacc2335a70113ee890eaf335dae74f8c69bc96e21a7562f87ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5841bb88d3e06bc498f2694341b10b26870a3bd6ed8785d8522ca8ac8536f2a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88e3b5045d8dfa462c759624f70bb3b703a2d64185d907de5fceafc5813c1857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5790c745e25dc060d772c86228021a868afae24905e421f6e112ba7e3aa40b56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2f235a75c3e0999d9df32aa6a8cb4fc44b2b027520ddaab195de00807b8cc05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15f26991cf1c5f1b915e015515fd0f8498e207124745835dafe352abef6170ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9916b82c53676d9b5cc57b66294504df981de54c66371352bdfe99f0f0861bcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7bef07802cc71eae0fde6ae9f5b67e90c4231bcfd30c82e873e696f90d86d98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cef6399590f8f677e63f65929b3d6e99c1cf684a83c0977eea6e876c0a140c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a6ea9687e34e1d998367fbd4acbb45a67d6898b9661012fa0e4fd3157e73e21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8df42e3de001da43ddee2fdc32aac3201b9a36ca1fe6ac30e7f4bd51de62790c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9878958e30525dfe08f4cc70338dc171a1c6a537e3ced1388b822f39f64c149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha02dd83fa709de166319479ece04b1ee165b0b6b095e6a8ca4ef7ab96751dd41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb558860cb9356a1d40ef7aefe5b77525031f1e0922f079f048af75a0dc677ba8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74ffb8004dbb892100c0ce497e0aec463caec9f6c18fe426c9bcaf0967675c5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c8dfc5998aaed1381f58019d86970ac823d4e6bee085a4c5c437c202b53a749;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf79e5cb7b633b69d6f140b806414f20690741e8b4252d697de8abad6adec94d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f4be92afea417f225d646f1d0f77642e421f8a8a52253c1498b365cf62db3ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ccd2e1b40a542cf7f3db81f12b1c86b932d438743e24ffda39680dd867ae7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h372ed65026cb98f6d600b77c6059f518384bedd96c3ad0cae15efabf20debc18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haca51b60367afd80b226370532aa874ba60cb10e0193d27696656621ab7f8798;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a6e01040a54c04bda2a892f054a351174ea86fc0db272c1b12a059191a0a82f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c08c17c7de200d049727ac69567f57661edcd76514a9992322f3a9ec7f0d230;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2def483e33f1b43fb420038ad693b3a234ae001563c56d467df481135ee07a26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92fa63cf84398198a4fadd66fc97e3063622c3d4e50498f4a3037535d755f6d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5290e5f75998c9e015a9638d7c973658d847184574cda2570e7870ab49f7dfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2740835317430176c39493c0054f9d11e41ae9b2e40ad51eb3201ae994392c6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55af938901794311d49dd8913450721f9366f97caa66535e6e11363e76f12d7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3fae6d95eeaaa6c8035b55bdf85a5860efe38de42190acd22942a58436240a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ab3deca0663dd6cf9cd3705ac788a6b61492ddbf164c50033ffbaeac3cf217c;
        #1
        $finish();
    end
endmodule
