module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    compressor_CLA64_32 compressor_CLA64_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
        src16 <= 64'h0;
        src17 <= 64'h0;
        src18 <= 64'h0;
        src19 <= 64'h0;
        src20 <= 64'h0;
        src21 <= 64'h0;
        src22 <= 64'h0;
        src23 <= 64'h0;
        src24 <= 64'h0;
        src25 <= 64'h0;
        src26 <= 64'h0;
        src27 <= 64'h0;
        src28 <= 64'h0;
        src29 <= 64'h0;
        src30 <= 64'h0;
        src31 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA64_32(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    input [63:0]src16,
    input [63:0]src17,
    input [63:0]src18,
    input [63:0]src19,
    input [63:0]src20,
    input [63:0]src21,
    input [63:0]src22,
    input [63:0]src23,
    input [63:0]src24,
    input [63:0]src25,
    input [63:0]src26,
    input [63:0]src27,
    input [63:0]src28,
    input [63:0]src29,
    input [63:0]src30,
    input [63:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [0:0] comp_out12;
    wire [0:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [0:0] comp_out36;
    wire [0:0] comp_out37;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], 1'h0, 1'h0, comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [0:0] dst36,
      output wire [0:0] dst37);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [63:0] stage0_16;
   wire [63:0] stage0_17;
   wire [63:0] stage0_18;
   wire [63:0] stage0_19;
   wire [63:0] stage0_20;
   wire [63:0] stage0_21;
   wire [63:0] stage0_22;
   wire [63:0] stage0_23;
   wire [63:0] stage0_24;
   wire [63:0] stage0_25;
   wire [63:0] stage0_26;
   wire [63:0] stage0_27;
   wire [63:0] stage0_28;
   wire [63:0] stage0_29;
   wire [63:0] stage0_30;
   wire [63:0] stage0_31;
   wire [23:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [31:0] stage1_3;
   wire [34:0] stage1_4;
   wire [34:0] stage1_5;
   wire [27:0] stage1_6;
   wire [23:0] stage1_7;
   wire [34:0] stage1_8;
   wire [27:0] stage1_9;
   wire [28:0] stage1_10;
   wire [28:0] stage1_11;
   wire [43:0] stage1_12;
   wire [22:0] stage1_13;
   wire [44:0] stage1_14;
   wire [31:0] stage1_15;
   wire [20:0] stage1_16;
   wire [34:0] stage1_17;
   wire [42:0] stage1_18;
   wire [19:0] stage1_19;
   wire [37:0] stage1_20;
   wire [27:0] stage1_21;
   wire [19:0] stage1_22;
   wire [47:0] stage1_23;
   wire [43:0] stage1_24;
   wire [23:0] stage1_25;
   wire [27:0] stage1_26;
   wire [21:0] stage1_27;
   wire [27:0] stage1_28;
   wire [37:0] stage1_29;
   wire [29:0] stage1_30;
   wire [27:0] stage1_31;
   wire [17:0] stage1_32;
   wire [8:0] stage1_33;
   wire [18:0] stage2_0;
   wire [5:0] stage2_1;
   wire [21:0] stage2_2;
   wire [17:0] stage2_3;
   wire [18:0] stage2_4;
   wire [26:0] stage2_5;
   wire [10:0] stage2_6;
   wire [8:0] stage2_7;
   wire [16:0] stage2_8;
   wire [15:0] stage2_9;
   wire [8:0] stage2_10;
   wire [11:0] stage2_11;
   wire [16:0] stage2_12;
   wire [17:0] stage2_13;
   wire [12:0] stage2_14;
   wire [23:0] stage2_15;
   wire [13:0] stage2_16;
   wire [13:0] stage2_17;
   wire [20:0] stage2_18;
   wire [15:0] stage2_19;
   wire [23:0] stage2_20;
   wire [12:0] stage2_21;
   wire [17:0] stage2_22;
   wire [16:0] stage2_23;
   wire [23:0] stage2_24;
   wire [17:0] stage2_25;
   wire [11:0] stage2_26;
   wire [16:0] stage2_27;
   wire [17:0] stage2_28;
   wire [17:0] stage2_29;
   wire [11:0] stage2_30;
   wire [21:0] stage2_31;
   wire [7:0] stage2_32;
   wire [7:0] stage2_33;
   wire [3:0] stage2_34;
   wire [0:0] stage2_35;
   wire [6:0] stage3_0;
   wire [5:0] stage3_1;
   wire [6:0] stage3_2;
   wire [6:0] stage3_3;
   wire [11:0] stage3_4;
   wire [5:0] stage3_5;
   wire [7:0] stage3_6;
   wire [10:0] stage3_7;
   wire [3:0] stage3_8;
   wire [7:0] stage3_9;
   wire [5:0] stage3_10;
   wire [3:0] stage3_11;
   wire [6:0] stage3_12;
   wire [8:0] stage3_13;
   wire [7:0] stage3_14;
   wire [6:0] stage3_15;
   wire [5:0] stage3_16;
   wire [7:0] stage3_17;
   wire [7:0] stage3_18;
   wire [12:0] stage3_19;
   wire [4:0] stage3_20;
   wire [8:0] stage3_21;
   wire [10:0] stage3_22;
   wire [6:0] stage3_23;
   wire [6:0] stage3_24;
   wire [8:0] stage3_25;
   wire [7:0] stage3_26;
   wire [4:0] stage3_27;
   wire [6:0] stage3_28;
   wire [8:0] stage3_29;
   wire [5:0] stage3_30;
   wire [8:0] stage3_31;
   wire [12:0] stage3_32;
   wire [6:0] stage3_33;
   wire [1:0] stage3_34;
   wire [0:0] stage3_35;
   wire [0:0] stage3_36;
   wire [0:0] stage3_37;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [2:0] stage4_2;
   wire [2:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [2:0] stage4_6;
   wire [5:0] stage4_7;
   wire [4:0] stage4_8;
   wire [2:0] stage4_9;
   wire [1:0] stage4_10;
   wire [2:0] stage4_11;
   wire [1:0] stage4_12;
   wire [5:0] stage4_13;
   wire [3:0] stage4_14;
   wire [2:0] stage4_15;
   wire [1:0] stage4_16;
   wire [4:0] stage4_17;
   wire [5:0] stage4_18;
   wire [2:0] stage4_19;
   wire [3:0] stage4_20;
   wire [4:0] stage4_21;
   wire [2:0] stage4_22;
   wire [3:0] stage4_23;
   wire [5:0] stage4_24;
   wire [3:0] stage4_25;
   wire [4:0] stage4_26;
   wire [2:0] stage4_27;
   wire [1:0] stage4_28;
   wire [4:0] stage4_29;
   wire [3:0] stage4_30;
   wire [3:0] stage4_31;
   wire [3:0] stage4_32;
   wire [3:0] stage4_33;
   wire [4:0] stage4_34;
   wire [1:0] stage4_35;
   wire [0:0] stage4_36;
   wire [0:0] stage4_37;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [0:0] stage5_12;
   wire [0:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [0:0] stage5_36;
   wire [0:0] stage5_37;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[3]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[4]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10]},
      {stage1_5[0],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage1_5[1],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage1_5[2],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28]},
      {stage1_5[3],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[4],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc606_5 gpc17 (
      {stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc606_5 gpc18 (
      {stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[7],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage0_4[18]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[8],stage1_4[19],stage1_3[19]}
   );
   gpc615_5 gpc20 (
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage0_4[19]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[9],stage1_4[20],stage1_3[20]}
   );
   gpc615_5 gpc21 (
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage0_4[20]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[5],stage1_5[10],stage1_4[21],stage1_3[21]}
   );
   gpc615_5 gpc22 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage0_4[21]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[6],stage1_5[11],stage1_4[22],stage1_3[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[4],stage1_6[7],stage1_5[12],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[5],stage1_6[8],stage1_5[13],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[6],stage1_6[9],stage1_5[14],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[7],stage1_6[10],stage1_5[15],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[8],stage1_6[11],stage1_5[16],stage1_4[27]}
   );
   gpc606_5 gpc28 (
      {stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[9],stage1_6[12],stage1_5[17],stage1_4[28]}
   );
   gpc606_5 gpc29 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[6],stage1_7[10],stage1_6[13],stage1_5[18]}
   );
   gpc606_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[7],stage1_7[11],stage1_6[14],stage1_5[19]}
   );
   gpc606_5 gpc31 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[8],stage1_7[12],stage1_6[15],stage1_5[20]}
   );
   gpc615_5 gpc32 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46]},
      {stage0_6[36]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[9],stage1_7[13],stage1_6[16],stage1_5[21]}
   );
   gpc615_5 gpc33 (
      {stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_6[37]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[10],stage1_7[14],stage1_6[17],stage1_5[22]}
   );
   gpc615_5 gpc34 (
      {stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage0_7[30]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[5],stage1_8[11],stage1_7[15],stage1_6[18]}
   );
   gpc615_5 gpc35 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[31]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[6],stage1_8[12],stage1_7[16],stage1_6[19]}
   );
   gpc615_5 gpc36 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[32]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[7],stage1_8[13],stage1_7[17],stage1_6[20]}
   );
   gpc615_5 gpc37 (
      {stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_7[33]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[8],stage1_8[14],stage1_7[18],stage1_6[21]}
   );
   gpc606_5 gpc38 (
      {stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[4],stage1_9[9],stage1_8[15],stage1_7[19]}
   );
   gpc606_5 gpc39 (
      {stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[5],stage1_9[10],stage1_8[16],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[6],stage1_9[11],stage1_8[17],stage1_7[21]}
   );
   gpc606_5 gpc41 (
      {stage0_7[52], stage0_7[53], stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[7],stage1_9[12],stage1_8[18],stage1_7[22]}
   );
   gpc606_5 gpc42 (
      {stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[8],stage1_9[13],stage1_8[19],stage1_7[23]}
   );
   gpc606_5 gpc43 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[5],stage1_10[9],stage1_9[14],stage1_8[20]}
   );
   gpc606_5 gpc44 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[6],stage1_10[10],stage1_9[15],stage1_8[21]}
   );
   gpc606_5 gpc45 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[7],stage1_10[11],stage1_9[16],stage1_8[22]}
   );
   gpc606_5 gpc46 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[8],stage1_10[12],stage1_9[17],stage1_8[23]}
   );
   gpc606_5 gpc47 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[9],stage1_10[13],stage1_9[18],stage1_8[24]}
   );
   gpc606_5 gpc48 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[5],stage1_11[10],stage1_10[14],stage1_9[19]}
   );
   gpc606_5 gpc49 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[6],stage1_11[11],stage1_10[15],stage1_9[20]}
   );
   gpc606_5 gpc50 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[7],stage1_11[12],stage1_10[16],stage1_9[21]}
   );
   gpc606_5 gpc51 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[8],stage1_11[13],stage1_10[17],stage1_9[22]}
   );
   gpc606_5 gpc52 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[9],stage1_11[14],stage1_10[18],stage1_9[23]}
   );
   gpc615_5 gpc53 (
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34]},
      {stage0_11[30]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[10],stage1_11[15],stage1_10[19]}
   );
   gpc615_5 gpc54 (
      {stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage0_11[31]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[6],stage1_12[11],stage1_11[16],stage1_10[20]}
   );
   gpc615_5 gpc55 (
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44]},
      {stage0_11[32]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[7],stage1_12[12],stage1_11[17],stage1_10[21]}
   );
   gpc615_5 gpc56 (
      {stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49]},
      {stage0_11[33]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[8],stage1_12[13],stage1_11[18],stage1_10[22]}
   );
   gpc615_5 gpc57 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[34]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[9],stage1_12[14],stage1_11[19],stage1_10[23]}
   );
   gpc615_5 gpc58 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage0_11[35]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[10],stage1_12[15],stage1_11[20],stage1_10[24]}
   );
   gpc615_5 gpc59 (
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage0_12[36]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[11],stage1_12[16],stage1_11[21]}
   );
   gpc615_5 gpc60 (
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45]},
      {stage0_12[37]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[7],stage1_13[12],stage1_12[17],stage1_11[22]}
   );
   gpc615_5 gpc61 (
      {stage0_11[46], stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50]},
      {stage0_12[38]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[8],stage1_13[13],stage1_12[18],stage1_11[23]}
   );
   gpc615_5 gpc62 (
      {stage0_11[51], stage0_11[52], stage0_11[53], stage0_11[54], stage0_11[55]},
      {stage0_12[39]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[9],stage1_13[14],stage1_12[19],stage1_11[24]}
   );
   gpc615_5 gpc63 (
      {stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_12[40]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[10],stage1_13[15],stage1_12[20],stage1_11[25]}
   );
   gpc615_5 gpc64 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34]},
      {stage0_14[0]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[0],stage1_15[5],stage1_14[11],stage1_13[16]}
   );
   gpc615_5 gpc65 (
      {stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39]},
      {stage0_14[1]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[1],stage1_15[6],stage1_14[12],stage1_13[17]}
   );
   gpc615_5 gpc66 (
      {stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44]},
      {stage0_14[2]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[2],stage1_15[7],stage1_14[13],stage1_13[18]}
   );
   gpc615_5 gpc67 (
      {stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage0_14[3]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[3],stage1_15[8],stage1_14[14],stage1_13[19]}
   );
   gpc615_5 gpc68 (
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54]},
      {stage0_14[4]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[4],stage1_15[9],stage1_14[15],stage1_13[20]}
   );
   gpc615_5 gpc69 (
      {stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_14[5]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[5],stage1_15[10],stage1_14[16],stage1_13[21]}
   );
   gpc615_5 gpc70 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], 1'b0},
      {stage0_14[6]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[6],stage1_15[11],stage1_14[17],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[7],stage1_16[7],stage1_15[12],stage1_14[18]}
   );
   gpc606_5 gpc72 (
      {stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[8],stage1_16[8],stage1_15[13],stage1_14[19]}
   );
   gpc606_5 gpc73 (
      {stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[9],stage1_16[9],stage1_15[14],stage1_14[20]}
   );
   gpc606_5 gpc74 (
      {stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[10],stage1_16[10],stage1_15[15],stage1_14[21]}
   );
   gpc606_5 gpc75 (
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[11],stage1_16[11],stage1_15[16],stage1_14[22]}
   );
   gpc606_5 gpc76 (
      {stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[12],stage1_16[12],stage1_15[17],stage1_14[23]}
   );
   gpc615_5 gpc77 (
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[13],stage1_16[13],stage1_15[18]}
   );
   gpc615_5 gpc78 (
      {stage0_15[47], stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[14],stage1_16[14],stage1_15[19]}
   );
   gpc606_5 gpc79 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[2],stage1_18[8],stage1_17[15],stage1_16[15]}
   );
   gpc606_5 gpc80 (
      {stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[3],stage1_18[9],stage1_17[16],stage1_16[16]}
   );
   gpc606_5 gpc81 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[4],stage1_18[10],stage1_17[17],stage1_16[17]}
   );
   gpc606_5 gpc82 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[5],stage1_18[11],stage1_17[18],stage1_16[18]}
   );
   gpc1163_5 gpc83 (
      {stage0_17[12], stage0_17[13], stage0_17[14]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage0_19[0]},
      {stage0_20[0]},
      {stage1_21[0],stage1_20[4],stage1_19[6],stage1_18[12],stage1_17[19]}
   );
   gpc1163_5 gpc84 (
      {stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage0_19[1]},
      {stage0_20[1]},
      {stage1_21[1],stage1_20[5],stage1_19[7],stage1_18[13],stage1_17[20]}
   );
   gpc1163_5 gpc85 (
      {stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_19[2]},
      {stage0_20[2]},
      {stage1_21[2],stage1_20[6],stage1_19[8],stage1_18[14],stage1_17[21]}
   );
   gpc606_5 gpc86 (
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26]},
      {stage0_19[3], stage0_19[4], stage0_19[5], stage0_19[6], stage0_19[7], stage0_19[8]},
      {stage1_21[3],stage1_20[7],stage1_19[9],stage1_18[15],stage1_17[22]}
   );
   gpc606_5 gpc87 (
      {stage0_17[27], stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32]},
      {stage0_19[9], stage0_19[10], stage0_19[11], stage0_19[12], stage0_19[13], stage0_19[14]},
      {stage1_21[4],stage1_20[8],stage1_19[10],stage1_18[16],stage1_17[23]}
   );
   gpc606_5 gpc88 (
      {stage0_17[33], stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38]},
      {stage0_19[15], stage0_19[16], stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20]},
      {stage1_21[5],stage1_20[9],stage1_19[11],stage1_18[17],stage1_17[24]}
   );
   gpc606_5 gpc89 (
      {stage0_17[39], stage0_17[40], stage0_17[41], stage0_17[42], stage0_17[43], stage0_17[44]},
      {stage0_19[21], stage0_19[22], stage0_19[23], stage0_19[24], stage0_19[25], stage0_19[26]},
      {stage1_21[6],stage1_20[10],stage1_19[12],stage1_18[18],stage1_17[25]}
   );
   gpc606_5 gpc90 (
      {stage0_17[45], stage0_17[46], stage0_17[47], stage0_17[48], stage0_17[49], stage0_17[50]},
      {stage0_19[27], stage0_19[28], stage0_19[29], stage0_19[30], stage0_19[31], stage0_19[32]},
      {stage1_21[7],stage1_20[11],stage1_19[13],stage1_18[19],stage1_17[26]}
   );
   gpc606_5 gpc91 (
      {stage0_17[51], stage0_17[52], stage0_17[53], stage0_17[54], stage0_17[55], stage0_17[56]},
      {stage0_19[33], stage0_19[34], stage0_19[35], stage0_19[36], stage0_19[37], stage0_19[38]},
      {stage1_21[8],stage1_20[12],stage1_19[14],stage1_18[20],stage1_17[27]}
   );
   gpc615_5 gpc92 (
      {stage0_19[39], stage0_19[40], stage0_19[41], stage0_19[42], stage0_19[43]},
      {stage0_20[3]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[9],stage1_20[13],stage1_19[15]}
   );
   gpc615_5 gpc93 (
      {stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48]},
      {stage0_20[4]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[1],stage1_21[10],stage1_20[14],stage1_19[16]}
   );
   gpc615_5 gpc94 (
      {stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage0_20[5]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[2],stage1_21[11],stage1_20[15],stage1_19[17]}
   );
   gpc615_5 gpc95 (
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58]},
      {stage0_20[6]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[3],stage1_21[12],stage1_20[16],stage1_19[18]}
   );
   gpc615_5 gpc96 (
      {stage0_19[59], stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63]},
      {stage0_20[7]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[4],stage1_21[13],stage1_20[17],stage1_19[19]}
   );
   gpc615_5 gpc97 (
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12]},
      {stage0_21[30]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[5],stage1_22[5],stage1_21[14],stage1_20[18]}
   );
   gpc615_5 gpc98 (
      {stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage0_21[31]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[6],stage1_22[6],stage1_21[15],stage1_20[19]}
   );
   gpc615_5 gpc99 (
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22]},
      {stage0_21[32]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[7],stage1_22[7],stage1_21[16],stage1_20[20]}
   );
   gpc615_5 gpc100 (
      {stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_21[33]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[8],stage1_22[8],stage1_21[17],stage1_20[21]}
   );
   gpc615_5 gpc101 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32]},
      {stage0_21[34]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[9],stage1_22[9],stage1_21[18],stage1_20[22]}
   );
   gpc615_5 gpc102 (
      {stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37]},
      {stage0_21[35]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[10],stage1_22[10],stage1_21[19],stage1_20[23]}
   );
   gpc615_5 gpc103 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[36]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[11],stage1_22[11],stage1_21[20],stage1_20[24]}
   );
   gpc615_5 gpc104 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[37]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[12],stage1_22[12],stage1_21[21],stage1_20[25]}
   );
   gpc615_5 gpc105 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[38]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[13],stage1_22[13],stage1_21[22],stage1_20[26]}
   );
   gpc615_5 gpc106 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43]},
      {stage0_22[54]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[9],stage1_23[14],stage1_22[14],stage1_21[23]}
   );
   gpc615_5 gpc107 (
      {stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48]},
      {stage0_22[55]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[10],stage1_23[15],stage1_22[15],stage1_21[24]}
   );
   gpc615_5 gpc108 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_22[56]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[11],stage1_23[16],stage1_22[16],stage1_21[25]}
   );
   gpc615_5 gpc109 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58]},
      {stage0_22[57]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[12],stage1_23[17],stage1_22[17],stage1_21[26]}
   );
   gpc615_5 gpc110 (
      {stage0_21[59], stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63]},
      {stage0_22[58]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[13],stage1_23[18],stage1_22[18],stage1_21[27]}
   );
   gpc615_5 gpc111 (
      {stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63]},
      {stage0_23[30]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[14],stage1_23[19],stage1_22[19]}
   );
   gpc606_5 gpc112 (
      {stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[6],stage1_24[15],stage1_23[20]}
   );
   gpc2135_5 gpc113 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10]},
      {stage0_25[6], stage0_25[7], stage0_25[8]},
      {stage0_26[0]},
      {stage0_27[0], stage0_27[1]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[7],stage1_24[16]}
   );
   gpc606_5 gpc114 (
      {stage0_24[11], stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16]},
      {stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5], stage0_26[6]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[8],stage1_24[17]}
   );
   gpc606_5 gpc115 (
      {stage0_24[17], stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22]},
      {stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11], stage0_26[12]},
      {stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[9],stage1_24[18]}
   );
   gpc615_5 gpc116 (
      {stage0_24[23], stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27]},
      {stage0_25[9]},
      {stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17], stage0_26[18]},
      {stage1_28[3],stage1_27[4],stage1_26[5],stage1_25[10],stage1_24[19]}
   );
   gpc615_5 gpc117 (
      {stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31], stage0_24[32]},
      {stage0_25[10]},
      {stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24]},
      {stage1_28[4],stage1_27[5],stage1_26[6],stage1_25[11],stage1_24[20]}
   );
   gpc615_5 gpc118 (
      {stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36], stage0_24[37]},
      {stage0_25[11]},
      {stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29], stage0_26[30]},
      {stage1_28[5],stage1_27[6],stage1_26[7],stage1_25[12],stage1_24[21]}
   );
   gpc615_5 gpc119 (
      {stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42]},
      {stage0_25[12]},
      {stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35], stage0_26[36]},
      {stage1_28[6],stage1_27[7],stage1_26[8],stage1_25[13],stage1_24[22]}
   );
   gpc606_5 gpc120 (
      {stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17], stage0_25[18]},
      {stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5], stage0_27[6], stage0_27[7]},
      {stage1_29[0],stage1_28[7],stage1_27[8],stage1_26[9],stage1_25[14]}
   );
   gpc606_5 gpc121 (
      {stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23], stage0_25[24]},
      {stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11], stage0_27[12], stage0_27[13]},
      {stage1_29[1],stage1_28[8],stage1_27[9],stage1_26[10],stage1_25[15]}
   );
   gpc615_5 gpc122 (
      {stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_26[37]},
      {stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17], stage0_27[18], stage0_27[19]},
      {stage1_29[2],stage1_28[9],stage1_27[10],stage1_26[11],stage1_25[16]}
   );
   gpc615_5 gpc123 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34]},
      {stage0_26[38]},
      {stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23], stage0_27[24], stage0_27[25]},
      {stage1_29[3],stage1_28[10],stage1_27[11],stage1_26[12],stage1_25[17]}
   );
   gpc615_5 gpc124 (
      {stage0_25[35], stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39]},
      {stage0_26[39]},
      {stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29], stage0_27[30], stage0_27[31]},
      {stage1_29[4],stage1_28[11],stage1_27[12],stage1_26[13],stage1_25[18]}
   );
   gpc615_5 gpc125 (
      {stage0_25[40], stage0_25[41], stage0_25[42], stage0_25[43], stage0_25[44]},
      {stage0_26[40]},
      {stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35], stage0_27[36], stage0_27[37]},
      {stage1_29[5],stage1_28[12],stage1_27[13],stage1_26[14],stage1_25[19]}
   );
   gpc615_5 gpc126 (
      {stage0_25[45], stage0_25[46], stage0_25[47], stage0_25[48], stage0_25[49]},
      {stage0_26[41]},
      {stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41], stage0_27[42], stage0_27[43]},
      {stage1_29[6],stage1_28[13],stage1_27[14],stage1_26[15],stage1_25[20]}
   );
   gpc615_5 gpc127 (
      {stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53], stage0_25[54]},
      {stage0_26[42]},
      {stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47], stage0_27[48], stage0_27[49]},
      {stage1_29[7],stage1_28[14],stage1_27[15],stage1_26[16],stage1_25[21]}
   );
   gpc615_5 gpc128 (
      {stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_26[43]},
      {stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53], stage0_27[54], stage0_27[55]},
      {stage1_29[8],stage1_28[15],stage1_27[16],stage1_26[17],stage1_25[22]}
   );
   gpc615_5 gpc129 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], 1'b0},
      {stage0_26[44]},
      {stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59], stage0_27[60], stage0_27[61]},
      {stage1_29[9],stage1_28[16],stage1_27[17],stage1_26[18],stage1_25[23]}
   );
   gpc606_5 gpc130 (
      {stage0_26[45], stage0_26[46], stage0_26[47], stage0_26[48], stage0_26[49], stage0_26[50]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[10],stage1_28[17],stage1_27[18],stage1_26[19]}
   );
   gpc606_5 gpc131 (
      {stage0_26[51], stage0_26[52], stage0_26[53], stage0_26[54], stage0_26[55], stage0_26[56]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[11],stage1_28[18],stage1_27[19],stage1_26[20]}
   );
   gpc606_5 gpc132 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[0],stage1_30[2],stage1_29[12],stage1_28[19]}
   );
   gpc606_5 gpc133 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[1],stage1_30[3],stage1_29[13],stage1_28[20]}
   );
   gpc606_5 gpc134 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[2],stage1_30[4],stage1_29[14],stage1_28[21]}
   );
   gpc606_5 gpc135 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[3],stage1_30[5],stage1_29[15],stage1_28[22]}
   );
   gpc606_5 gpc136 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[4],stage1_30[6],stage1_29[16],stage1_28[23]}
   );
   gpc606_5 gpc137 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[5],stage1_30[7],stage1_29[17],stage1_28[24]}
   );
   gpc606_5 gpc138 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[6],stage1_30[8],stage1_29[18],stage1_28[25]}
   );
   gpc615_5 gpc139 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58]},
      {stage0_29[0]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[7],stage1_30[9],stage1_29[19],stage1_28[26]}
   );
   gpc615_5 gpc140 (
      {stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63]},
      {stage0_29[1]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[8],stage1_30[10],stage1_29[20],stage1_28[27]}
   );
   gpc606_5 gpc141 (
      {stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5], stage0_29[6], stage0_29[7]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[9],stage1_30[11],stage1_29[21]}
   );
   gpc606_5 gpc142 (
      {stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[10],stage1_30[12],stage1_29[22]}
   );
   gpc606_5 gpc143 (
      {stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[11],stage1_30[13],stage1_29[23]}
   );
   gpc606_5 gpc144 (
      {stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[12],stage1_30[14],stage1_29[24]}
   );
   gpc606_5 gpc145 (
      {stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[13],stage1_30[15],stage1_29[25]}
   );
   gpc606_5 gpc146 (
      {stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[14],stage1_30[16],stage1_29[26]}
   );
   gpc606_5 gpc147 (
      {stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[15],stage1_30[17],stage1_29[27]}
   );
   gpc606_5 gpc148 (
      {stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[16],stage1_30[18],stage1_29[28]}
   );
   gpc606_5 gpc149 (
      {stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[17],stage1_31[17],stage1_30[19],stage1_29[29]}
   );
   gpc1_1 gpc150 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc151 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc152 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc153 (
      {stage0_0[54]},
      {stage1_0[14]}
   );
   gpc1_1 gpc154 (
      {stage0_0[55]},
      {stage1_0[15]}
   );
   gpc1_1 gpc155 (
      {stage0_0[56]},
      {stage1_0[16]}
   );
   gpc1_1 gpc156 (
      {stage0_0[57]},
      {stage1_0[17]}
   );
   gpc1_1 gpc157 (
      {stage0_0[58]},
      {stage1_0[18]}
   );
   gpc1_1 gpc158 (
      {stage0_0[59]},
      {stage1_0[19]}
   );
   gpc1_1 gpc159 (
      {stage0_0[60]},
      {stage1_0[20]}
   );
   gpc1_1 gpc160 (
      {stage0_0[61]},
      {stage1_0[21]}
   );
   gpc1_1 gpc161 (
      {stage0_0[62]},
      {stage1_0[22]}
   );
   gpc1_1 gpc162 (
      {stage0_0[63]},
      {stage1_0[23]}
   );
   gpc1_1 gpc163 (
      {stage0_1[60]},
      {stage1_1[16]}
   );
   gpc1_1 gpc164 (
      {stage0_1[61]},
      {stage1_1[17]}
   );
   gpc1_1 gpc165 (
      {stage0_1[62]},
      {stage1_1[18]}
   );
   gpc1_1 gpc166 (
      {stage0_1[63]},
      {stage1_1[19]}
   );
   gpc1_1 gpc167 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc168 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc169 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc170 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc171 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc172 (
      {stage0_3[55]},
      {stage1_3[23]}
   );
   gpc1_1 gpc173 (
      {stage0_3[56]},
      {stage1_3[24]}
   );
   gpc1_1 gpc174 (
      {stage0_3[57]},
      {stage1_3[25]}
   );
   gpc1_1 gpc175 (
      {stage0_3[58]},
      {stage1_3[26]}
   );
   gpc1_1 gpc176 (
      {stage0_3[59]},
      {stage1_3[27]}
   );
   gpc1_1 gpc177 (
      {stage0_3[60]},
      {stage1_3[28]}
   );
   gpc1_1 gpc178 (
      {stage0_3[61]},
      {stage1_3[29]}
   );
   gpc1_1 gpc179 (
      {stage0_3[62]},
      {stage1_3[30]}
   );
   gpc1_1 gpc180 (
      {stage0_3[63]},
      {stage1_3[31]}
   );
   gpc1_1 gpc181 (
      {stage0_4[58]},
      {stage1_4[29]}
   );
   gpc1_1 gpc182 (
      {stage0_4[59]},
      {stage1_4[30]}
   );
   gpc1_1 gpc183 (
      {stage0_4[60]},
      {stage1_4[31]}
   );
   gpc1_1 gpc184 (
      {stage0_4[61]},
      {stage1_4[32]}
   );
   gpc1_1 gpc185 (
      {stage0_4[62]},
      {stage1_4[33]}
   );
   gpc1_1 gpc186 (
      {stage0_4[63]},
      {stage1_4[34]}
   );
   gpc1_1 gpc187 (
      {stage0_5[52]},
      {stage1_5[23]}
   );
   gpc1_1 gpc188 (
      {stage0_5[53]},
      {stage1_5[24]}
   );
   gpc1_1 gpc189 (
      {stage0_5[54]},
      {stage1_5[25]}
   );
   gpc1_1 gpc190 (
      {stage0_5[55]},
      {stage1_5[26]}
   );
   gpc1_1 gpc191 (
      {stage0_5[56]},
      {stage1_5[27]}
   );
   gpc1_1 gpc192 (
      {stage0_5[57]},
      {stage1_5[28]}
   );
   gpc1_1 gpc193 (
      {stage0_5[58]},
      {stage1_5[29]}
   );
   gpc1_1 gpc194 (
      {stage0_5[59]},
      {stage1_5[30]}
   );
   gpc1_1 gpc195 (
      {stage0_5[60]},
      {stage1_5[31]}
   );
   gpc1_1 gpc196 (
      {stage0_5[61]},
      {stage1_5[32]}
   );
   gpc1_1 gpc197 (
      {stage0_5[62]},
      {stage1_5[33]}
   );
   gpc1_1 gpc198 (
      {stage0_5[63]},
      {stage1_5[34]}
   );
   gpc1_1 gpc199 (
      {stage0_6[58]},
      {stage1_6[22]}
   );
   gpc1_1 gpc200 (
      {stage0_6[59]},
      {stage1_6[23]}
   );
   gpc1_1 gpc201 (
      {stage0_6[60]},
      {stage1_6[24]}
   );
   gpc1_1 gpc202 (
      {stage0_6[61]},
      {stage1_6[25]}
   );
   gpc1_1 gpc203 (
      {stage0_6[62]},
      {stage1_6[26]}
   );
   gpc1_1 gpc204 (
      {stage0_6[63]},
      {stage1_6[27]}
   );
   gpc1_1 gpc205 (
      {stage0_8[54]},
      {stage1_8[25]}
   );
   gpc1_1 gpc206 (
      {stage0_8[55]},
      {stage1_8[26]}
   );
   gpc1_1 gpc207 (
      {stage0_8[56]},
      {stage1_8[27]}
   );
   gpc1_1 gpc208 (
      {stage0_8[57]},
      {stage1_8[28]}
   );
   gpc1_1 gpc209 (
      {stage0_8[58]},
      {stage1_8[29]}
   );
   gpc1_1 gpc210 (
      {stage0_8[59]},
      {stage1_8[30]}
   );
   gpc1_1 gpc211 (
      {stage0_8[60]},
      {stage1_8[31]}
   );
   gpc1_1 gpc212 (
      {stage0_8[61]},
      {stage1_8[32]}
   );
   gpc1_1 gpc213 (
      {stage0_8[62]},
      {stage1_8[33]}
   );
   gpc1_1 gpc214 (
      {stage0_8[63]},
      {stage1_8[34]}
   );
   gpc1_1 gpc215 (
      {stage0_9[60]},
      {stage1_9[24]}
   );
   gpc1_1 gpc216 (
      {stage0_9[61]},
      {stage1_9[25]}
   );
   gpc1_1 gpc217 (
      {stage0_9[62]},
      {stage1_9[26]}
   );
   gpc1_1 gpc218 (
      {stage0_9[63]},
      {stage1_9[27]}
   );
   gpc1_1 gpc219 (
      {stage0_10[60]},
      {stage1_10[25]}
   );
   gpc1_1 gpc220 (
      {stage0_10[61]},
      {stage1_10[26]}
   );
   gpc1_1 gpc221 (
      {stage0_10[62]},
      {stage1_10[27]}
   );
   gpc1_1 gpc222 (
      {stage0_10[63]},
      {stage1_10[28]}
   );
   gpc1_1 gpc223 (
      {stage0_11[61]},
      {stage1_11[26]}
   );
   gpc1_1 gpc224 (
      {stage0_11[62]},
      {stage1_11[27]}
   );
   gpc1_1 gpc225 (
      {stage0_11[63]},
      {stage1_11[28]}
   );
   gpc1_1 gpc226 (
      {stage0_12[41]},
      {stage1_12[21]}
   );
   gpc1_1 gpc227 (
      {stage0_12[42]},
      {stage1_12[22]}
   );
   gpc1_1 gpc228 (
      {stage0_12[43]},
      {stage1_12[23]}
   );
   gpc1_1 gpc229 (
      {stage0_12[44]},
      {stage1_12[24]}
   );
   gpc1_1 gpc230 (
      {stage0_12[45]},
      {stage1_12[25]}
   );
   gpc1_1 gpc231 (
      {stage0_12[46]},
      {stage1_12[26]}
   );
   gpc1_1 gpc232 (
      {stage0_12[47]},
      {stage1_12[27]}
   );
   gpc1_1 gpc233 (
      {stage0_12[48]},
      {stage1_12[28]}
   );
   gpc1_1 gpc234 (
      {stage0_12[49]},
      {stage1_12[29]}
   );
   gpc1_1 gpc235 (
      {stage0_12[50]},
      {stage1_12[30]}
   );
   gpc1_1 gpc236 (
      {stage0_12[51]},
      {stage1_12[31]}
   );
   gpc1_1 gpc237 (
      {stage0_12[52]},
      {stage1_12[32]}
   );
   gpc1_1 gpc238 (
      {stage0_12[53]},
      {stage1_12[33]}
   );
   gpc1_1 gpc239 (
      {stage0_12[54]},
      {stage1_12[34]}
   );
   gpc1_1 gpc240 (
      {stage0_12[55]},
      {stage1_12[35]}
   );
   gpc1_1 gpc241 (
      {stage0_12[56]},
      {stage1_12[36]}
   );
   gpc1_1 gpc242 (
      {stage0_12[57]},
      {stage1_12[37]}
   );
   gpc1_1 gpc243 (
      {stage0_12[58]},
      {stage1_12[38]}
   );
   gpc1_1 gpc244 (
      {stage0_12[59]},
      {stage1_12[39]}
   );
   gpc1_1 gpc245 (
      {stage0_12[60]},
      {stage1_12[40]}
   );
   gpc1_1 gpc246 (
      {stage0_12[61]},
      {stage1_12[41]}
   );
   gpc1_1 gpc247 (
      {stage0_12[62]},
      {stage1_12[42]}
   );
   gpc1_1 gpc248 (
      {stage0_12[63]},
      {stage1_12[43]}
   );
   gpc1_1 gpc249 (
      {stage0_14[43]},
      {stage1_14[24]}
   );
   gpc1_1 gpc250 (
      {stage0_14[44]},
      {stage1_14[25]}
   );
   gpc1_1 gpc251 (
      {stage0_14[45]},
      {stage1_14[26]}
   );
   gpc1_1 gpc252 (
      {stage0_14[46]},
      {stage1_14[27]}
   );
   gpc1_1 gpc253 (
      {stage0_14[47]},
      {stage1_14[28]}
   );
   gpc1_1 gpc254 (
      {stage0_14[48]},
      {stage1_14[29]}
   );
   gpc1_1 gpc255 (
      {stage0_14[49]},
      {stage1_14[30]}
   );
   gpc1_1 gpc256 (
      {stage0_14[50]},
      {stage1_14[31]}
   );
   gpc1_1 gpc257 (
      {stage0_14[51]},
      {stage1_14[32]}
   );
   gpc1_1 gpc258 (
      {stage0_14[52]},
      {stage1_14[33]}
   );
   gpc1_1 gpc259 (
      {stage0_14[53]},
      {stage1_14[34]}
   );
   gpc1_1 gpc260 (
      {stage0_14[54]},
      {stage1_14[35]}
   );
   gpc1_1 gpc261 (
      {stage0_14[55]},
      {stage1_14[36]}
   );
   gpc1_1 gpc262 (
      {stage0_14[56]},
      {stage1_14[37]}
   );
   gpc1_1 gpc263 (
      {stage0_14[57]},
      {stage1_14[38]}
   );
   gpc1_1 gpc264 (
      {stage0_14[58]},
      {stage1_14[39]}
   );
   gpc1_1 gpc265 (
      {stage0_14[59]},
      {stage1_14[40]}
   );
   gpc1_1 gpc266 (
      {stage0_14[60]},
      {stage1_14[41]}
   );
   gpc1_1 gpc267 (
      {stage0_14[61]},
      {stage1_14[42]}
   );
   gpc1_1 gpc268 (
      {stage0_14[62]},
      {stage1_14[43]}
   );
   gpc1_1 gpc269 (
      {stage0_14[63]},
      {stage1_14[44]}
   );
   gpc1_1 gpc270 (
      {stage0_15[52]},
      {stage1_15[20]}
   );
   gpc1_1 gpc271 (
      {stage0_15[53]},
      {stage1_15[21]}
   );
   gpc1_1 gpc272 (
      {stage0_15[54]},
      {stage1_15[22]}
   );
   gpc1_1 gpc273 (
      {stage0_15[55]},
      {stage1_15[23]}
   );
   gpc1_1 gpc274 (
      {stage0_15[56]},
      {stage1_15[24]}
   );
   gpc1_1 gpc275 (
      {stage0_15[57]},
      {stage1_15[25]}
   );
   gpc1_1 gpc276 (
      {stage0_15[58]},
      {stage1_15[26]}
   );
   gpc1_1 gpc277 (
      {stage0_15[59]},
      {stage1_15[27]}
   );
   gpc1_1 gpc278 (
      {stage0_15[60]},
      {stage1_15[28]}
   );
   gpc1_1 gpc279 (
      {stage0_15[61]},
      {stage1_15[29]}
   );
   gpc1_1 gpc280 (
      {stage0_15[62]},
      {stage1_15[30]}
   );
   gpc1_1 gpc281 (
      {stage0_15[63]},
      {stage1_15[31]}
   );
   gpc1_1 gpc282 (
      {stage0_16[62]},
      {stage1_16[19]}
   );
   gpc1_1 gpc283 (
      {stage0_16[63]},
      {stage1_16[20]}
   );
   gpc1_1 gpc284 (
      {stage0_17[57]},
      {stage1_17[28]}
   );
   gpc1_1 gpc285 (
      {stage0_17[58]},
      {stage1_17[29]}
   );
   gpc1_1 gpc286 (
      {stage0_17[59]},
      {stage1_17[30]}
   );
   gpc1_1 gpc287 (
      {stage0_17[60]},
      {stage1_17[31]}
   );
   gpc1_1 gpc288 (
      {stage0_17[61]},
      {stage1_17[32]}
   );
   gpc1_1 gpc289 (
      {stage0_17[62]},
      {stage1_17[33]}
   );
   gpc1_1 gpc290 (
      {stage0_17[63]},
      {stage1_17[34]}
   );
   gpc1_1 gpc291 (
      {stage0_18[42]},
      {stage1_18[21]}
   );
   gpc1_1 gpc292 (
      {stage0_18[43]},
      {stage1_18[22]}
   );
   gpc1_1 gpc293 (
      {stage0_18[44]},
      {stage1_18[23]}
   );
   gpc1_1 gpc294 (
      {stage0_18[45]},
      {stage1_18[24]}
   );
   gpc1_1 gpc295 (
      {stage0_18[46]},
      {stage1_18[25]}
   );
   gpc1_1 gpc296 (
      {stage0_18[47]},
      {stage1_18[26]}
   );
   gpc1_1 gpc297 (
      {stage0_18[48]},
      {stage1_18[27]}
   );
   gpc1_1 gpc298 (
      {stage0_18[49]},
      {stage1_18[28]}
   );
   gpc1_1 gpc299 (
      {stage0_18[50]},
      {stage1_18[29]}
   );
   gpc1_1 gpc300 (
      {stage0_18[51]},
      {stage1_18[30]}
   );
   gpc1_1 gpc301 (
      {stage0_18[52]},
      {stage1_18[31]}
   );
   gpc1_1 gpc302 (
      {stage0_18[53]},
      {stage1_18[32]}
   );
   gpc1_1 gpc303 (
      {stage0_18[54]},
      {stage1_18[33]}
   );
   gpc1_1 gpc304 (
      {stage0_18[55]},
      {stage1_18[34]}
   );
   gpc1_1 gpc305 (
      {stage0_18[56]},
      {stage1_18[35]}
   );
   gpc1_1 gpc306 (
      {stage0_18[57]},
      {stage1_18[36]}
   );
   gpc1_1 gpc307 (
      {stage0_18[58]},
      {stage1_18[37]}
   );
   gpc1_1 gpc308 (
      {stage0_18[59]},
      {stage1_18[38]}
   );
   gpc1_1 gpc309 (
      {stage0_18[60]},
      {stage1_18[39]}
   );
   gpc1_1 gpc310 (
      {stage0_18[61]},
      {stage1_18[40]}
   );
   gpc1_1 gpc311 (
      {stage0_18[62]},
      {stage1_18[41]}
   );
   gpc1_1 gpc312 (
      {stage0_18[63]},
      {stage1_18[42]}
   );
   gpc1_1 gpc313 (
      {stage0_20[53]},
      {stage1_20[27]}
   );
   gpc1_1 gpc314 (
      {stage0_20[54]},
      {stage1_20[28]}
   );
   gpc1_1 gpc315 (
      {stage0_20[55]},
      {stage1_20[29]}
   );
   gpc1_1 gpc316 (
      {stage0_20[56]},
      {stage1_20[30]}
   );
   gpc1_1 gpc317 (
      {stage0_20[57]},
      {stage1_20[31]}
   );
   gpc1_1 gpc318 (
      {stage0_20[58]},
      {stage1_20[32]}
   );
   gpc1_1 gpc319 (
      {stage0_20[59]},
      {stage1_20[33]}
   );
   gpc1_1 gpc320 (
      {stage0_20[60]},
      {stage1_20[34]}
   );
   gpc1_1 gpc321 (
      {stage0_20[61]},
      {stage1_20[35]}
   );
   gpc1_1 gpc322 (
      {stage0_20[62]},
      {stage1_20[36]}
   );
   gpc1_1 gpc323 (
      {stage0_20[63]},
      {stage1_20[37]}
   );
   gpc1_1 gpc324 (
      {stage0_23[37]},
      {stage1_23[21]}
   );
   gpc1_1 gpc325 (
      {stage0_23[38]},
      {stage1_23[22]}
   );
   gpc1_1 gpc326 (
      {stage0_23[39]},
      {stage1_23[23]}
   );
   gpc1_1 gpc327 (
      {stage0_23[40]},
      {stage1_23[24]}
   );
   gpc1_1 gpc328 (
      {stage0_23[41]},
      {stage1_23[25]}
   );
   gpc1_1 gpc329 (
      {stage0_23[42]},
      {stage1_23[26]}
   );
   gpc1_1 gpc330 (
      {stage0_23[43]},
      {stage1_23[27]}
   );
   gpc1_1 gpc331 (
      {stage0_23[44]},
      {stage1_23[28]}
   );
   gpc1_1 gpc332 (
      {stage0_23[45]},
      {stage1_23[29]}
   );
   gpc1_1 gpc333 (
      {stage0_23[46]},
      {stage1_23[30]}
   );
   gpc1_1 gpc334 (
      {stage0_23[47]},
      {stage1_23[31]}
   );
   gpc1_1 gpc335 (
      {stage0_23[48]},
      {stage1_23[32]}
   );
   gpc1_1 gpc336 (
      {stage0_23[49]},
      {stage1_23[33]}
   );
   gpc1_1 gpc337 (
      {stage0_23[50]},
      {stage1_23[34]}
   );
   gpc1_1 gpc338 (
      {stage0_23[51]},
      {stage1_23[35]}
   );
   gpc1_1 gpc339 (
      {stage0_23[52]},
      {stage1_23[36]}
   );
   gpc1_1 gpc340 (
      {stage0_23[53]},
      {stage1_23[37]}
   );
   gpc1_1 gpc341 (
      {stage0_23[54]},
      {stage1_23[38]}
   );
   gpc1_1 gpc342 (
      {stage0_23[55]},
      {stage1_23[39]}
   );
   gpc1_1 gpc343 (
      {stage0_23[56]},
      {stage1_23[40]}
   );
   gpc1_1 gpc344 (
      {stage0_23[57]},
      {stage1_23[41]}
   );
   gpc1_1 gpc345 (
      {stage0_23[58]},
      {stage1_23[42]}
   );
   gpc1_1 gpc346 (
      {stage0_23[59]},
      {stage1_23[43]}
   );
   gpc1_1 gpc347 (
      {stage0_23[60]},
      {stage1_23[44]}
   );
   gpc1_1 gpc348 (
      {stage0_23[61]},
      {stage1_23[45]}
   );
   gpc1_1 gpc349 (
      {stage0_23[62]},
      {stage1_23[46]}
   );
   gpc1_1 gpc350 (
      {stage0_23[63]},
      {stage1_23[47]}
   );
   gpc1_1 gpc351 (
      {stage0_24[43]},
      {stage1_24[23]}
   );
   gpc1_1 gpc352 (
      {stage0_24[44]},
      {stage1_24[24]}
   );
   gpc1_1 gpc353 (
      {stage0_24[45]},
      {stage1_24[25]}
   );
   gpc1_1 gpc354 (
      {stage0_24[46]},
      {stage1_24[26]}
   );
   gpc1_1 gpc355 (
      {stage0_24[47]},
      {stage1_24[27]}
   );
   gpc1_1 gpc356 (
      {stage0_24[48]},
      {stage1_24[28]}
   );
   gpc1_1 gpc357 (
      {stage0_24[49]},
      {stage1_24[29]}
   );
   gpc1_1 gpc358 (
      {stage0_24[50]},
      {stage1_24[30]}
   );
   gpc1_1 gpc359 (
      {stage0_24[51]},
      {stage1_24[31]}
   );
   gpc1_1 gpc360 (
      {stage0_24[52]},
      {stage1_24[32]}
   );
   gpc1_1 gpc361 (
      {stage0_24[53]},
      {stage1_24[33]}
   );
   gpc1_1 gpc362 (
      {stage0_24[54]},
      {stage1_24[34]}
   );
   gpc1_1 gpc363 (
      {stage0_24[55]},
      {stage1_24[35]}
   );
   gpc1_1 gpc364 (
      {stage0_24[56]},
      {stage1_24[36]}
   );
   gpc1_1 gpc365 (
      {stage0_24[57]},
      {stage1_24[37]}
   );
   gpc1_1 gpc366 (
      {stage0_24[58]},
      {stage1_24[38]}
   );
   gpc1_1 gpc367 (
      {stage0_24[59]},
      {stage1_24[39]}
   );
   gpc1_1 gpc368 (
      {stage0_24[60]},
      {stage1_24[40]}
   );
   gpc1_1 gpc369 (
      {stage0_24[61]},
      {stage1_24[41]}
   );
   gpc1_1 gpc370 (
      {stage0_24[62]},
      {stage1_24[42]}
   );
   gpc1_1 gpc371 (
      {stage0_24[63]},
      {stage1_24[43]}
   );
   gpc1_1 gpc372 (
      {stage0_26[57]},
      {stage1_26[21]}
   );
   gpc1_1 gpc373 (
      {stage0_26[58]},
      {stage1_26[22]}
   );
   gpc1_1 gpc374 (
      {stage0_26[59]},
      {stage1_26[23]}
   );
   gpc1_1 gpc375 (
      {stage0_26[60]},
      {stage1_26[24]}
   );
   gpc1_1 gpc376 (
      {stage0_26[61]},
      {stage1_26[25]}
   );
   gpc1_1 gpc377 (
      {stage0_26[62]},
      {stage1_26[26]}
   );
   gpc1_1 gpc378 (
      {stage0_26[63]},
      {stage1_26[27]}
   );
   gpc1_1 gpc379 (
      {stage0_27[62]},
      {stage1_27[20]}
   );
   gpc1_1 gpc380 (
      {stage0_27[63]},
      {stage1_27[21]}
   );
   gpc1_1 gpc381 (
      {stage0_29[56]},
      {stage1_29[30]}
   );
   gpc1_1 gpc382 (
      {stage0_29[57]},
      {stage1_29[31]}
   );
   gpc1_1 gpc383 (
      {stage0_29[58]},
      {stage1_29[32]}
   );
   gpc1_1 gpc384 (
      {stage0_29[59]},
      {stage1_29[33]}
   );
   gpc1_1 gpc385 (
      {stage0_29[60]},
      {stage1_29[34]}
   );
   gpc1_1 gpc386 (
      {stage0_29[61]},
      {stage1_29[35]}
   );
   gpc1_1 gpc387 (
      {stage0_29[62]},
      {stage1_29[36]}
   );
   gpc1_1 gpc388 (
      {stage0_29[63]},
      {stage1_29[37]}
   );
   gpc1_1 gpc389 (
      {stage0_30[54]},
      {stage1_30[20]}
   );
   gpc1_1 gpc390 (
      {stage0_30[55]},
      {stage1_30[21]}
   );
   gpc1_1 gpc391 (
      {stage0_30[56]},
      {stage1_30[22]}
   );
   gpc1_1 gpc392 (
      {stage0_30[57]},
      {stage1_30[23]}
   );
   gpc1_1 gpc393 (
      {stage0_30[58]},
      {stage1_30[24]}
   );
   gpc1_1 gpc394 (
      {stage0_30[59]},
      {stage1_30[25]}
   );
   gpc1_1 gpc395 (
      {stage0_30[60]},
      {stage1_30[26]}
   );
   gpc1_1 gpc396 (
      {stage0_30[61]},
      {stage1_30[27]}
   );
   gpc1_1 gpc397 (
      {stage0_30[62]},
      {stage1_30[28]}
   );
   gpc1_1 gpc398 (
      {stage0_30[63]},
      {stage1_30[29]}
   );
   gpc1_1 gpc399 (
      {stage0_31[54]},
      {stage1_31[18]}
   );
   gpc1_1 gpc400 (
      {stage0_31[55]},
      {stage1_31[19]}
   );
   gpc1_1 gpc401 (
      {stage0_31[56]},
      {stage1_31[20]}
   );
   gpc1_1 gpc402 (
      {stage0_31[57]},
      {stage1_31[21]}
   );
   gpc1_1 gpc403 (
      {stage0_31[58]},
      {stage1_31[22]}
   );
   gpc1_1 gpc404 (
      {stage0_31[59]},
      {stage1_31[23]}
   );
   gpc1_1 gpc405 (
      {stage0_31[60]},
      {stage1_31[24]}
   );
   gpc1_1 gpc406 (
      {stage0_31[61]},
      {stage1_31[25]}
   );
   gpc1_1 gpc407 (
      {stage0_31[62]},
      {stage1_31[26]}
   );
   gpc1_1 gpc408 (
      {stage0_31[63]},
      {stage1_31[27]}
   );
   gpc606_5 gpc409 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc410 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc411 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc412 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc413 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[3],stage2_4[4]}
   );
   gpc606_5 gpc414 (
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[4],stage2_4[5]}
   );
   gpc606_5 gpc415 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[5],stage2_4[6]}
   );
   gpc606_5 gpc416 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[3],stage2_6[3],stage2_5[6],stage2_4[7]}
   );
   gpc606_5 gpc417 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[4],stage2_6[4],stage2_5[7]}
   );
   gpc606_5 gpc418 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[5],stage2_7[5],stage2_6[5],stage2_5[8]}
   );
   gpc606_5 gpc419 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[6],stage2_7[6],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc420 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[3],stage2_8[7],stage2_7[7]}
   );
   gpc606_5 gpc421 (
      {stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[1],stage2_9[4],stage2_8[8]}
   );
   gpc606_5 gpc422 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[2],stage2_9[5],stage2_8[9]}
   );
   gpc606_5 gpc423 (
      {stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[3],stage2_9[6],stage2_8[10]}
   );
   gpc606_5 gpc424 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[4],stage2_10[4],stage2_9[7],stage2_8[11]}
   );
   gpc606_5 gpc425 (
      {stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], 1'b0},
      {stage2_12[4],stage2_11[5],stage2_10[5],stage2_9[8],stage2_8[12]}
   );
   gpc606_5 gpc426 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[6],stage2_10[6],stage2_9[9]}
   );
   gpc606_5 gpc427 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[7],stage2_10[7],stage2_9[10]}
   );
   gpc606_5 gpc428 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[8],stage2_10[8],stage2_9[11]}
   );
   gpc615_5 gpc429 (
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22]},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[3],stage2_12[8],stage2_11[9]}
   );
   gpc615_5 gpc430 (
      {stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27]},
      {stage1_12[1]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[1],stage2_13[4],stage2_12[9],stage2_11[10]}
   );
   gpc606_5 gpc431 (
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[2],stage2_14[2],stage2_13[5],stage2_12[10]}
   );
   gpc606_5 gpc432 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[3],stage2_14[3],stage2_13[6],stage2_12[11]}
   );
   gpc606_5 gpc433 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[4],stage2_14[4],stage2_13[7],stage2_12[12]}
   );
   gpc606_5 gpc434 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[5],stage2_14[5],stage2_13[8],stage2_12[13]}
   );
   gpc606_5 gpc435 (
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[6],stage2_14[6],stage2_13[9],stage2_12[14]}
   );
   gpc606_5 gpc436 (
      {stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[7],stage2_14[7],stage2_13[10],stage2_12[15]}
   );
   gpc606_5 gpc437 (
      {stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[8],stage2_14[8],stage2_13[11],stage2_12[16]}
   );
   gpc606_5 gpc438 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[9],stage2_14[9],stage2_13[12]}
   );
   gpc615_5 gpc439 (
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[8],stage2_15[10]}
   );
   gpc615_5 gpc440 (
      {stage1_15[11], stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[9],stage2_15[11]}
   );
   gpc615_5 gpc441 (
      {stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19], stage1_15[20]},
      {stage1_16[2]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[2],stage2_17[3],stage2_16[10],stage2_15[12]}
   );
   gpc606_5 gpc442 (
      {stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6], stage1_16[7], stage1_16[8]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[3],stage2_18[3],stage2_17[4],stage2_16[11]}
   );
   gpc606_5 gpc443 (
      {stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13], stage1_16[14]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[4],stage2_18[4],stage2_17[5],stage2_16[12]}
   );
   gpc606_5 gpc444 (
      {stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[5],stage2_18[5],stage2_17[6],stage2_16[13]}
   );
   gpc606_5 gpc445 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[3],stage2_19[6],stage2_18[6],stage2_17[7]}
   );
   gpc606_5 gpc446 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[4],stage2_19[7],stage2_18[7],stage2_17[8]}
   );
   gpc615_5 gpc447 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage1_19[12]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[5],stage2_19[8],stage2_18[8]}
   );
   gpc615_5 gpc448 (
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27]},
      {stage1_19[13]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[3],stage2_20[6],stage2_19[9],stage2_18[9]}
   );
   gpc615_5 gpc449 (
      {stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31], stage1_18[32]},
      {stage1_19[14]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[4],stage2_20[7],stage2_19[10],stage2_18[10]}
   );
   gpc615_5 gpc450 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22]},
      {stage1_21[0]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[0],stage2_22[3],stage2_21[5],stage2_20[8]}
   );
   gpc606_5 gpc451 (
      {stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5], stage1_21[6]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[1],stage2_22[4],stage2_21[6]}
   );
   gpc606_5 gpc452 (
      {stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11], stage1_21[12]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[2],stage2_22[5],stage2_21[7]}
   );
   gpc606_5 gpc453 (
      {stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17], stage1_21[18]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[3],stage2_22[6],stage2_21[8]}
   );
   gpc606_5 gpc454 (
      {stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23], stage1_21[24]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[4],stage2_23[4],stage2_22[7],stage2_21[9]}
   );
   gpc615_5 gpc455 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10]},
      {stage1_23[24]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[5],stage2_23[5],stage2_22[8]}
   );
   gpc615_5 gpc456 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage1_24[6]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[1],stage2_25[5],stage2_24[6],stage2_23[6]}
   );
   gpc615_5 gpc457 (
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34]},
      {stage1_24[7]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[2],stage2_25[6],stage2_24[7],stage2_23[7]}
   );
   gpc615_5 gpc458 (
      {stage1_23[35], stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39]},
      {stage1_24[8]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[3],stage2_25[7],stage2_24[8],stage2_23[8]}
   );
   gpc606_5 gpc459 (
      {stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13], stage1_24[14]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[3],stage2_26[4],stage2_25[8],stage2_24[9]}
   );
   gpc606_5 gpc460 (
      {stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19], stage1_24[20]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[4],stage2_26[5],stage2_25[9],stage2_24[10]}
   );
   gpc606_5 gpc461 (
      {stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25], stage1_24[26]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[5],stage2_26[6],stage2_25[10],stage2_24[11]}
   );
   gpc606_5 gpc462 (
      {stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30], stage1_24[31], stage1_24[32]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[6],stage2_26[7],stage2_25[11],stage2_24[12]}
   );
   gpc615_5 gpc463 (
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4]},
      {stage1_28[0]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[0],stage2_28[4],stage2_27[7]}
   );
   gpc615_5 gpc464 (
      {stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage1_28[1]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[1],stage2_29[1],stage2_28[5],stage2_27[8]}
   );
   gpc615_5 gpc465 (
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14]},
      {stage1_28[2]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[2],stage2_29[2],stage2_28[6],stage2_27[9]}
   );
   gpc2135_5 gpc466 (
      {stage1_28[3], stage1_28[4], stage1_28[5], stage1_28[6], stage1_28[7]},
      {stage1_29[18], stage1_29[19], stage1_29[20]},
      {stage1_30[0]},
      {stage1_31[0], stage1_31[1]},
      {stage2_32[0],stage2_31[3],stage2_30[3],stage2_29[3],stage2_28[7]}
   );
   gpc606_5 gpc467 (
      {stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13]},
      {stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6]},
      {stage2_32[1],stage2_31[4],stage2_30[4],stage2_29[4],stage2_28[8]}
   );
   gpc606_5 gpc468 (
      {stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19]},
      {stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12]},
      {stage2_32[2],stage2_31[5],stage2_30[5],stage2_29[5],stage2_28[9]}
   );
   gpc606_5 gpc469 (
      {stage1_29[21], stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25], stage1_29[26]},
      {stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7]},
      {stage2_33[0],stage2_32[3],stage2_31[6],stage2_30[6],stage2_29[6]}
   );
   gpc615_5 gpc470 (
      {stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage1_31[8]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[4],stage2_31[7],stage2_30[7]}
   );
   gpc615_5 gpc471 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22]},
      {stage1_31[9]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[2],stage2_32[5],stage2_31[8],stage2_30[8]}
   );
   gpc615_5 gpc472 (
      {stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27]},
      {stage1_31[10]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[3],stage2_32[6],stage2_31[9],stage2_30[9]}
   );
   gpc606_5 gpc473 (
      {stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[3],stage2_33[4],stage2_32[7],stage2_31[10]}
   );
   gpc1_1 gpc474 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc475 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc476 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc477 (
      {stage1_0[9]},
      {stage2_0[4]}
   );
   gpc1_1 gpc478 (
      {stage1_0[10]},
      {stage2_0[5]}
   );
   gpc1_1 gpc479 (
      {stage1_0[11]},
      {stage2_0[6]}
   );
   gpc1_1 gpc480 (
      {stage1_0[12]},
      {stage2_0[7]}
   );
   gpc1_1 gpc481 (
      {stage1_0[13]},
      {stage2_0[8]}
   );
   gpc1_1 gpc482 (
      {stage1_0[14]},
      {stage2_0[9]}
   );
   gpc1_1 gpc483 (
      {stage1_0[15]},
      {stage2_0[10]}
   );
   gpc1_1 gpc484 (
      {stage1_0[16]},
      {stage2_0[11]}
   );
   gpc1_1 gpc485 (
      {stage1_0[17]},
      {stage2_0[12]}
   );
   gpc1_1 gpc486 (
      {stage1_0[18]},
      {stage2_0[13]}
   );
   gpc1_1 gpc487 (
      {stage1_0[19]},
      {stage2_0[14]}
   );
   gpc1_1 gpc488 (
      {stage1_0[20]},
      {stage2_0[15]}
   );
   gpc1_1 gpc489 (
      {stage1_0[21]},
      {stage2_0[16]}
   );
   gpc1_1 gpc490 (
      {stage1_0[22]},
      {stage2_0[17]}
   );
   gpc1_1 gpc491 (
      {stage1_0[23]},
      {stage2_0[18]}
   );
   gpc1_1 gpc492 (
      {stage1_1[18]},
      {stage2_1[4]}
   );
   gpc1_1 gpc493 (
      {stage1_1[19]},
      {stage2_1[5]}
   );
   gpc1_1 gpc494 (
      {stage1_2[6]},
      {stage2_2[4]}
   );
   gpc1_1 gpc495 (
      {stage1_2[7]},
      {stage2_2[5]}
   );
   gpc1_1 gpc496 (
      {stage1_2[8]},
      {stage2_2[6]}
   );
   gpc1_1 gpc497 (
      {stage1_2[9]},
      {stage2_2[7]}
   );
   gpc1_1 gpc498 (
      {stage1_2[10]},
      {stage2_2[8]}
   );
   gpc1_1 gpc499 (
      {stage1_2[11]},
      {stage2_2[9]}
   );
   gpc1_1 gpc500 (
      {stage1_2[12]},
      {stage2_2[10]}
   );
   gpc1_1 gpc501 (
      {stage1_2[13]},
      {stage2_2[11]}
   );
   gpc1_1 gpc502 (
      {stage1_2[14]},
      {stage2_2[12]}
   );
   gpc1_1 gpc503 (
      {stage1_2[15]},
      {stage2_2[13]}
   );
   gpc1_1 gpc504 (
      {stage1_2[16]},
      {stage2_2[14]}
   );
   gpc1_1 gpc505 (
      {stage1_2[17]},
      {stage2_2[15]}
   );
   gpc1_1 gpc506 (
      {stage1_2[18]},
      {stage2_2[16]}
   );
   gpc1_1 gpc507 (
      {stage1_2[19]},
      {stage2_2[17]}
   );
   gpc1_1 gpc508 (
      {stage1_2[20]},
      {stage2_2[18]}
   );
   gpc1_1 gpc509 (
      {stage1_2[21]},
      {stage2_2[19]}
   );
   gpc1_1 gpc510 (
      {stage1_2[22]},
      {stage2_2[20]}
   );
   gpc1_1 gpc511 (
      {stage1_2[23]},
      {stage2_2[21]}
   );
   gpc1_1 gpc512 (
      {stage1_3[18]},
      {stage2_3[4]}
   );
   gpc1_1 gpc513 (
      {stage1_3[19]},
      {stage2_3[5]}
   );
   gpc1_1 gpc514 (
      {stage1_3[20]},
      {stage2_3[6]}
   );
   gpc1_1 gpc515 (
      {stage1_3[21]},
      {stage2_3[7]}
   );
   gpc1_1 gpc516 (
      {stage1_3[22]},
      {stage2_3[8]}
   );
   gpc1_1 gpc517 (
      {stage1_3[23]},
      {stage2_3[9]}
   );
   gpc1_1 gpc518 (
      {stage1_3[24]},
      {stage2_3[10]}
   );
   gpc1_1 gpc519 (
      {stage1_3[25]},
      {stage2_3[11]}
   );
   gpc1_1 gpc520 (
      {stage1_3[26]},
      {stage2_3[12]}
   );
   gpc1_1 gpc521 (
      {stage1_3[27]},
      {stage2_3[13]}
   );
   gpc1_1 gpc522 (
      {stage1_3[28]},
      {stage2_3[14]}
   );
   gpc1_1 gpc523 (
      {stage1_3[29]},
      {stage2_3[15]}
   );
   gpc1_1 gpc524 (
      {stage1_3[30]},
      {stage2_3[16]}
   );
   gpc1_1 gpc525 (
      {stage1_3[31]},
      {stage2_3[17]}
   );
   gpc1_1 gpc526 (
      {stage1_4[24]},
      {stage2_4[8]}
   );
   gpc1_1 gpc527 (
      {stage1_4[25]},
      {stage2_4[9]}
   );
   gpc1_1 gpc528 (
      {stage1_4[26]},
      {stage2_4[10]}
   );
   gpc1_1 gpc529 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1_1 gpc530 (
      {stage1_4[28]},
      {stage2_4[12]}
   );
   gpc1_1 gpc531 (
      {stage1_4[29]},
      {stage2_4[13]}
   );
   gpc1_1 gpc532 (
      {stage1_4[30]},
      {stage2_4[14]}
   );
   gpc1_1 gpc533 (
      {stage1_4[31]},
      {stage2_4[15]}
   );
   gpc1_1 gpc534 (
      {stage1_4[32]},
      {stage2_4[16]}
   );
   gpc1_1 gpc535 (
      {stage1_4[33]},
      {stage2_4[17]}
   );
   gpc1_1 gpc536 (
      {stage1_4[34]},
      {stage2_4[18]}
   );
   gpc1_1 gpc537 (
      {stage1_5[18]},
      {stage2_5[10]}
   );
   gpc1_1 gpc538 (
      {stage1_5[19]},
      {stage2_5[11]}
   );
   gpc1_1 gpc539 (
      {stage1_5[20]},
      {stage2_5[12]}
   );
   gpc1_1 gpc540 (
      {stage1_5[21]},
      {stage2_5[13]}
   );
   gpc1_1 gpc541 (
      {stage1_5[22]},
      {stage2_5[14]}
   );
   gpc1_1 gpc542 (
      {stage1_5[23]},
      {stage2_5[15]}
   );
   gpc1_1 gpc543 (
      {stage1_5[24]},
      {stage2_5[16]}
   );
   gpc1_1 gpc544 (
      {stage1_5[25]},
      {stage2_5[17]}
   );
   gpc1_1 gpc545 (
      {stage1_5[26]},
      {stage2_5[18]}
   );
   gpc1_1 gpc546 (
      {stage1_5[27]},
      {stage2_5[19]}
   );
   gpc1_1 gpc547 (
      {stage1_5[28]},
      {stage2_5[20]}
   );
   gpc1_1 gpc548 (
      {stage1_5[29]},
      {stage2_5[21]}
   );
   gpc1_1 gpc549 (
      {stage1_5[30]},
      {stage2_5[22]}
   );
   gpc1_1 gpc550 (
      {stage1_5[31]},
      {stage2_5[23]}
   );
   gpc1_1 gpc551 (
      {stage1_5[32]},
      {stage2_5[24]}
   );
   gpc1_1 gpc552 (
      {stage1_5[33]},
      {stage2_5[25]}
   );
   gpc1_1 gpc553 (
      {stage1_5[34]},
      {stage2_5[26]}
   );
   gpc1_1 gpc554 (
      {stage1_6[24]},
      {stage2_6[7]}
   );
   gpc1_1 gpc555 (
      {stage1_6[25]},
      {stage2_6[8]}
   );
   gpc1_1 gpc556 (
      {stage1_6[26]},
      {stage2_6[9]}
   );
   gpc1_1 gpc557 (
      {stage1_6[27]},
      {stage2_6[10]}
   );
   gpc1_1 gpc558 (
      {stage1_7[23]},
      {stage2_7[8]}
   );
   gpc1_1 gpc559 (
      {stage1_8[31]},
      {stage2_8[13]}
   );
   gpc1_1 gpc560 (
      {stage1_8[32]},
      {stage2_8[14]}
   );
   gpc1_1 gpc561 (
      {stage1_8[33]},
      {stage2_8[15]}
   );
   gpc1_1 gpc562 (
      {stage1_8[34]},
      {stage2_8[16]}
   );
   gpc1_1 gpc563 (
      {stage1_9[24]},
      {stage2_9[12]}
   );
   gpc1_1 gpc564 (
      {stage1_9[25]},
      {stage2_9[13]}
   );
   gpc1_1 gpc565 (
      {stage1_9[26]},
      {stage2_9[14]}
   );
   gpc1_1 gpc566 (
      {stage1_9[27]},
      {stage2_9[15]}
   );
   gpc1_1 gpc567 (
      {stage1_11[28]},
      {stage2_11[11]}
   );
   gpc1_1 gpc568 (
      {stage1_13[18]},
      {stage2_13[13]}
   );
   gpc1_1 gpc569 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc570 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc1_1 gpc571 (
      {stage1_13[21]},
      {stage2_13[16]}
   );
   gpc1_1 gpc572 (
      {stage1_13[22]},
      {stage2_13[17]}
   );
   gpc1_1 gpc573 (
      {stage1_14[42]},
      {stage2_14[10]}
   );
   gpc1_1 gpc574 (
      {stage1_14[43]},
      {stage2_14[11]}
   );
   gpc1_1 gpc575 (
      {stage1_14[44]},
      {stage2_14[12]}
   );
   gpc1_1 gpc576 (
      {stage1_15[21]},
      {stage2_15[13]}
   );
   gpc1_1 gpc577 (
      {stage1_15[22]},
      {stage2_15[14]}
   );
   gpc1_1 gpc578 (
      {stage1_15[23]},
      {stage2_15[15]}
   );
   gpc1_1 gpc579 (
      {stage1_15[24]},
      {stage2_15[16]}
   );
   gpc1_1 gpc580 (
      {stage1_15[25]},
      {stage2_15[17]}
   );
   gpc1_1 gpc581 (
      {stage1_15[26]},
      {stage2_15[18]}
   );
   gpc1_1 gpc582 (
      {stage1_15[27]},
      {stage2_15[19]}
   );
   gpc1_1 gpc583 (
      {stage1_15[28]},
      {stage2_15[20]}
   );
   gpc1_1 gpc584 (
      {stage1_15[29]},
      {stage2_15[21]}
   );
   gpc1_1 gpc585 (
      {stage1_15[30]},
      {stage2_15[22]}
   );
   gpc1_1 gpc586 (
      {stage1_15[31]},
      {stage2_15[23]}
   );
   gpc1_1 gpc587 (
      {stage1_17[30]},
      {stage2_17[9]}
   );
   gpc1_1 gpc588 (
      {stage1_17[31]},
      {stage2_17[10]}
   );
   gpc1_1 gpc589 (
      {stage1_17[32]},
      {stage2_17[11]}
   );
   gpc1_1 gpc590 (
      {stage1_17[33]},
      {stage2_17[12]}
   );
   gpc1_1 gpc591 (
      {stage1_17[34]},
      {stage2_17[13]}
   );
   gpc1_1 gpc592 (
      {stage1_18[33]},
      {stage2_18[11]}
   );
   gpc1_1 gpc593 (
      {stage1_18[34]},
      {stage2_18[12]}
   );
   gpc1_1 gpc594 (
      {stage1_18[35]},
      {stage2_18[13]}
   );
   gpc1_1 gpc595 (
      {stage1_18[36]},
      {stage2_18[14]}
   );
   gpc1_1 gpc596 (
      {stage1_18[37]},
      {stage2_18[15]}
   );
   gpc1_1 gpc597 (
      {stage1_18[38]},
      {stage2_18[16]}
   );
   gpc1_1 gpc598 (
      {stage1_18[39]},
      {stage2_18[17]}
   );
   gpc1_1 gpc599 (
      {stage1_18[40]},
      {stage2_18[18]}
   );
   gpc1_1 gpc600 (
      {stage1_18[41]},
      {stage2_18[19]}
   );
   gpc1_1 gpc601 (
      {stage1_18[42]},
      {stage2_18[20]}
   );
   gpc1_1 gpc602 (
      {stage1_19[15]},
      {stage2_19[11]}
   );
   gpc1_1 gpc603 (
      {stage1_19[16]},
      {stage2_19[12]}
   );
   gpc1_1 gpc604 (
      {stage1_19[17]},
      {stage2_19[13]}
   );
   gpc1_1 gpc605 (
      {stage1_19[18]},
      {stage2_19[14]}
   );
   gpc1_1 gpc606 (
      {stage1_19[19]},
      {stage2_19[15]}
   );
   gpc1_1 gpc607 (
      {stage1_20[23]},
      {stage2_20[9]}
   );
   gpc1_1 gpc608 (
      {stage1_20[24]},
      {stage2_20[10]}
   );
   gpc1_1 gpc609 (
      {stage1_20[25]},
      {stage2_20[11]}
   );
   gpc1_1 gpc610 (
      {stage1_20[26]},
      {stage2_20[12]}
   );
   gpc1_1 gpc611 (
      {stage1_20[27]},
      {stage2_20[13]}
   );
   gpc1_1 gpc612 (
      {stage1_20[28]},
      {stage2_20[14]}
   );
   gpc1_1 gpc613 (
      {stage1_20[29]},
      {stage2_20[15]}
   );
   gpc1_1 gpc614 (
      {stage1_20[30]},
      {stage2_20[16]}
   );
   gpc1_1 gpc615 (
      {stage1_20[31]},
      {stage2_20[17]}
   );
   gpc1_1 gpc616 (
      {stage1_20[32]},
      {stage2_20[18]}
   );
   gpc1_1 gpc617 (
      {stage1_20[33]},
      {stage2_20[19]}
   );
   gpc1_1 gpc618 (
      {stage1_20[34]},
      {stage2_20[20]}
   );
   gpc1_1 gpc619 (
      {stage1_20[35]},
      {stage2_20[21]}
   );
   gpc1_1 gpc620 (
      {stage1_20[36]},
      {stage2_20[22]}
   );
   gpc1_1 gpc621 (
      {stage1_20[37]},
      {stage2_20[23]}
   );
   gpc1_1 gpc622 (
      {stage1_21[25]},
      {stage2_21[10]}
   );
   gpc1_1 gpc623 (
      {stage1_21[26]},
      {stage2_21[11]}
   );
   gpc1_1 gpc624 (
      {stage1_21[27]},
      {stage2_21[12]}
   );
   gpc1_1 gpc625 (
      {stage1_22[11]},
      {stage2_22[9]}
   );
   gpc1_1 gpc626 (
      {stage1_22[12]},
      {stage2_22[10]}
   );
   gpc1_1 gpc627 (
      {stage1_22[13]},
      {stage2_22[11]}
   );
   gpc1_1 gpc628 (
      {stage1_22[14]},
      {stage2_22[12]}
   );
   gpc1_1 gpc629 (
      {stage1_22[15]},
      {stage2_22[13]}
   );
   gpc1_1 gpc630 (
      {stage1_22[16]},
      {stage2_22[14]}
   );
   gpc1_1 gpc631 (
      {stage1_22[17]},
      {stage2_22[15]}
   );
   gpc1_1 gpc632 (
      {stage1_22[18]},
      {stage2_22[16]}
   );
   gpc1_1 gpc633 (
      {stage1_22[19]},
      {stage2_22[17]}
   );
   gpc1_1 gpc634 (
      {stage1_23[40]},
      {stage2_23[9]}
   );
   gpc1_1 gpc635 (
      {stage1_23[41]},
      {stage2_23[10]}
   );
   gpc1_1 gpc636 (
      {stage1_23[42]},
      {stage2_23[11]}
   );
   gpc1_1 gpc637 (
      {stage1_23[43]},
      {stage2_23[12]}
   );
   gpc1_1 gpc638 (
      {stage1_23[44]},
      {stage2_23[13]}
   );
   gpc1_1 gpc639 (
      {stage1_23[45]},
      {stage2_23[14]}
   );
   gpc1_1 gpc640 (
      {stage1_23[46]},
      {stage2_23[15]}
   );
   gpc1_1 gpc641 (
      {stage1_23[47]},
      {stage2_23[16]}
   );
   gpc1_1 gpc642 (
      {stage1_24[33]},
      {stage2_24[13]}
   );
   gpc1_1 gpc643 (
      {stage1_24[34]},
      {stage2_24[14]}
   );
   gpc1_1 gpc644 (
      {stage1_24[35]},
      {stage2_24[15]}
   );
   gpc1_1 gpc645 (
      {stage1_24[36]},
      {stage2_24[16]}
   );
   gpc1_1 gpc646 (
      {stage1_24[37]},
      {stage2_24[17]}
   );
   gpc1_1 gpc647 (
      {stage1_24[38]},
      {stage2_24[18]}
   );
   gpc1_1 gpc648 (
      {stage1_24[39]},
      {stage2_24[19]}
   );
   gpc1_1 gpc649 (
      {stage1_24[40]},
      {stage2_24[20]}
   );
   gpc1_1 gpc650 (
      {stage1_24[41]},
      {stage2_24[21]}
   );
   gpc1_1 gpc651 (
      {stage1_24[42]},
      {stage2_24[22]}
   );
   gpc1_1 gpc652 (
      {stage1_24[43]},
      {stage2_24[23]}
   );
   gpc1_1 gpc653 (
      {stage1_25[18]},
      {stage2_25[12]}
   );
   gpc1_1 gpc654 (
      {stage1_25[19]},
      {stage2_25[13]}
   );
   gpc1_1 gpc655 (
      {stage1_25[20]},
      {stage2_25[14]}
   );
   gpc1_1 gpc656 (
      {stage1_25[21]},
      {stage2_25[15]}
   );
   gpc1_1 gpc657 (
      {stage1_25[22]},
      {stage2_25[16]}
   );
   gpc1_1 gpc658 (
      {stage1_25[23]},
      {stage2_25[17]}
   );
   gpc1_1 gpc659 (
      {stage1_26[24]},
      {stage2_26[8]}
   );
   gpc1_1 gpc660 (
      {stage1_26[25]},
      {stage2_26[9]}
   );
   gpc1_1 gpc661 (
      {stage1_26[26]},
      {stage2_26[10]}
   );
   gpc1_1 gpc662 (
      {stage1_26[27]},
      {stage2_26[11]}
   );
   gpc1_1 gpc663 (
      {stage1_27[15]},
      {stage2_27[10]}
   );
   gpc1_1 gpc664 (
      {stage1_27[16]},
      {stage2_27[11]}
   );
   gpc1_1 gpc665 (
      {stage1_27[17]},
      {stage2_27[12]}
   );
   gpc1_1 gpc666 (
      {stage1_27[18]},
      {stage2_27[13]}
   );
   gpc1_1 gpc667 (
      {stage1_27[19]},
      {stage2_27[14]}
   );
   gpc1_1 gpc668 (
      {stage1_27[20]},
      {stage2_27[15]}
   );
   gpc1_1 gpc669 (
      {stage1_27[21]},
      {stage2_27[16]}
   );
   gpc1_1 gpc670 (
      {stage1_28[20]},
      {stage2_28[10]}
   );
   gpc1_1 gpc671 (
      {stage1_28[21]},
      {stage2_28[11]}
   );
   gpc1_1 gpc672 (
      {stage1_28[22]},
      {stage2_28[12]}
   );
   gpc1_1 gpc673 (
      {stage1_28[23]},
      {stage2_28[13]}
   );
   gpc1_1 gpc674 (
      {stage1_28[24]},
      {stage2_28[14]}
   );
   gpc1_1 gpc675 (
      {stage1_28[25]},
      {stage2_28[15]}
   );
   gpc1_1 gpc676 (
      {stage1_28[26]},
      {stage2_28[16]}
   );
   gpc1_1 gpc677 (
      {stage1_28[27]},
      {stage2_28[17]}
   );
   gpc1_1 gpc678 (
      {stage1_29[27]},
      {stage2_29[7]}
   );
   gpc1_1 gpc679 (
      {stage1_29[28]},
      {stage2_29[8]}
   );
   gpc1_1 gpc680 (
      {stage1_29[29]},
      {stage2_29[9]}
   );
   gpc1_1 gpc681 (
      {stage1_29[30]},
      {stage2_29[10]}
   );
   gpc1_1 gpc682 (
      {stage1_29[31]},
      {stage2_29[11]}
   );
   gpc1_1 gpc683 (
      {stage1_29[32]},
      {stage2_29[12]}
   );
   gpc1_1 gpc684 (
      {stage1_29[33]},
      {stage2_29[13]}
   );
   gpc1_1 gpc685 (
      {stage1_29[34]},
      {stage2_29[14]}
   );
   gpc1_1 gpc686 (
      {stage1_29[35]},
      {stage2_29[15]}
   );
   gpc1_1 gpc687 (
      {stage1_29[36]},
      {stage2_29[16]}
   );
   gpc1_1 gpc688 (
      {stage1_29[37]},
      {stage2_29[17]}
   );
   gpc1_1 gpc689 (
      {stage1_30[28]},
      {stage2_30[10]}
   );
   gpc1_1 gpc690 (
      {stage1_30[29]},
      {stage2_30[11]}
   );
   gpc1_1 gpc691 (
      {stage1_31[17]},
      {stage2_31[11]}
   );
   gpc1_1 gpc692 (
      {stage1_31[18]},
      {stage2_31[12]}
   );
   gpc1_1 gpc693 (
      {stage1_31[19]},
      {stage2_31[13]}
   );
   gpc1_1 gpc694 (
      {stage1_31[20]},
      {stage2_31[14]}
   );
   gpc1_1 gpc695 (
      {stage1_31[21]},
      {stage2_31[15]}
   );
   gpc1_1 gpc696 (
      {stage1_31[22]},
      {stage2_31[16]}
   );
   gpc1_1 gpc697 (
      {stage1_31[23]},
      {stage2_31[17]}
   );
   gpc1_1 gpc698 (
      {stage1_31[24]},
      {stage2_31[18]}
   );
   gpc1_1 gpc699 (
      {stage1_31[25]},
      {stage2_31[19]}
   );
   gpc1_1 gpc700 (
      {stage1_31[26]},
      {stage2_31[20]}
   );
   gpc1_1 gpc701 (
      {stage1_31[27]},
      {stage2_31[21]}
   );
   gpc1_1 gpc702 (
      {stage1_33[6]},
      {stage2_33[5]}
   );
   gpc1_1 gpc703 (
      {stage1_33[7]},
      {stage2_33[6]}
   );
   gpc1_1 gpc704 (
      {stage1_33[8]},
      {stage2_33[7]}
   );
   gpc615_5 gpc705 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc706 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc707 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[2]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc708 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[3],stage3_3[3]}
   );
   gpc606_5 gpc709 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc710 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[0]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[5],stage3_3[5]}
   );
   gpc135_4 gpc711 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_5[18], stage2_5[19], stage2_5[20]},
      {stage2_6[0]},
      {stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[6]}
   );
   gpc135_4 gpc712 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_6[1]},
      {stage3_7[4],stage3_6[4],stage3_5[4],stage3_4[7]}
   );
   gpc135_4 gpc713 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[24], stage2_5[25], stage2_5[26]},
      {stage2_6[2]},
      {stage3_7[5],stage3_6[5],stage3_5[5],stage3_4[8]}
   );
   gpc615_5 gpc714 (
      {stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[6],stage3_6[6]}
   );
   gpc615_5 gpc715 (
      {stage2_6[8], stage2_6[9], stage2_6[10], 1'b0, 1'b0},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[1],stage3_7[7],stage3_6[7]}
   );
   gpc615_5 gpc716 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[2],stage3_7[8]}
   );
   gpc615_5 gpc717 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], 1'b0},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[3]}
   );
   gpc606_5 gpc718 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[4],stage3_9[4]}
   );
   gpc1163_5 gpc719 (
      {stage2_10[6], stage2_10[7], stage2_10[8]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[5]}
   );
   gpc207_4 gpc720 (
      {stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3]}
   );
   gpc207_4 gpc721 (
      {stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[2], stage2_14[3]},
      {stage3_15[1],stage3_14[2],stage3_13[3],stage3_12[4]}
   );
   gpc615_5 gpc722 (
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_14[4]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[0],stage3_15[2],stage3_14[3],stage3_13[4]}
   );
   gpc615_5 gpc723 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10]},
      {stage2_14[5]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[1],stage3_15[3],stage3_14[4],stage3_13[5]}
   );
   gpc615_5 gpc724 (
      {stage2_13[11], stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15]},
      {stage2_14[6]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[2],stage3_15[4],stage3_14[5],stage3_13[6]}
   );
   gpc615_5 gpc725 (
      {stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_15[18]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[3],stage3_15[5],stage3_14[6]}
   );
   gpc615_5 gpc726 (
      {stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[4],stage3_15[6]}
   );
   gpc117_4 gpc727 (
      {stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11], stage2_16[12], stage2_16[13]},
      {stage2_17[6]},
      {stage2_18[0]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[5]}
   );
   gpc606_5 gpc728 (
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[2],stage3_18[3],stage3_17[6]}
   );
   gpc615_5 gpc729 (
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage2_19[6]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[3],stage3_18[4]}
   );
   gpc615_5 gpc730 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[7]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[2],stage3_20[2],stage3_19[4],stage3_18[5]}
   );
   gpc615_5 gpc731 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[8]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[3],stage3_20[3],stage3_19[5],stage3_18[6]}
   );
   gpc615_5 gpc732 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[9]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[4],stage3_20[4],stage3_19[6],stage3_18[7]}
   );
   gpc606_5 gpc733 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[4],stage3_21[5]}
   );
   gpc615_5 gpc734 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10]},
      {stage2_22[0]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[5],stage3_21[6]}
   );
   gpc615_5 gpc735 (
      {stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[6]}
   );
   gpc615_5 gpc736 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[7]}
   );
   gpc615_5 gpc737 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[8]}
   );
   gpc615_5 gpc738 (
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[3],stage3_25[5],stage3_24[5]}
   );
   gpc606_5 gpc739 (
      {stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[4],stage3_25[6]}
   );
   gpc606_5 gpc740 (
      {stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[5],stage3_25[7]}
   );
   gpc606_5 gpc741 (
      {stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], 1'b0},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], 1'b0},
      {stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[6],stage3_25[8]}
   );
   gpc606_5 gpc742 (
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[7]}
   );
   gpc606_5 gpc743 (
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[4],stage3_28[5]}
   );
   gpc606_5 gpc744 (
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[1],stage3_30[2],stage3_29[5],stage3_28[6]}
   );
   gpc606_5 gpc745 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[2],stage3_31[2],stage3_30[3],stage3_29[6]}
   );
   gpc606_5 gpc746 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[3],stage3_31[3],stage3_30[4],stage3_29[7]}
   );
   gpc606_5 gpc747 (
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[4],stage3_31[4],stage3_30[5],stage3_29[8]}
   );
   gpc2135_5 gpc748 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4]},
      {stage2_34[0], stage2_34[1], stage2_34[2]},
      {stage2_35[0]},
      {1'b0, 1'b0},
      {stage3_37[0],stage3_36[0],stage3_35[0],stage3_34[0],stage3_33[3]}
   );
   gpc1_1 gpc749 (
      {stage2_0[15]},
      {stage3_0[3]}
   );
   gpc1_1 gpc750 (
      {stage2_0[16]},
      {stage3_0[4]}
   );
   gpc1_1 gpc751 (
      {stage2_0[17]},
      {stage3_0[5]}
   );
   gpc1_1 gpc752 (
      {stage2_0[18]},
      {stage3_0[6]}
   );
   gpc1_1 gpc753 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc754 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc755 (
      {stage2_1[5]},
      {stage3_1[5]}
   );
   gpc1_1 gpc756 (
      {stage2_2[18]},
      {stage3_2[3]}
   );
   gpc1_1 gpc757 (
      {stage2_2[19]},
      {stage3_2[4]}
   );
   gpc1_1 gpc758 (
      {stage2_2[20]},
      {stage3_2[5]}
   );
   gpc1_1 gpc759 (
      {stage2_2[21]},
      {stage3_2[6]}
   );
   gpc1_1 gpc760 (
      {stage2_3[17]},
      {stage3_3[6]}
   );
   gpc1_1 gpc761 (
      {stage2_4[16]},
      {stage3_4[9]}
   );
   gpc1_1 gpc762 (
      {stage2_4[17]},
      {stage3_4[10]}
   );
   gpc1_1 gpc763 (
      {stage2_4[18]},
      {stage3_4[11]}
   );
   gpc1_1 gpc764 (
      {stage2_7[7]},
      {stage3_7[9]}
   );
   gpc1_1 gpc765 (
      {stage2_7[8]},
      {stage3_7[10]}
   );
   gpc1_1 gpc766 (
      {stage2_9[13]},
      {stage3_9[5]}
   );
   gpc1_1 gpc767 (
      {stage2_9[14]},
      {stage3_9[6]}
   );
   gpc1_1 gpc768 (
      {stage2_9[15]},
      {stage3_9[7]}
   );
   gpc1_1 gpc769 (
      {stage2_12[15]},
      {stage3_12[5]}
   );
   gpc1_1 gpc770 (
      {stage2_12[16]},
      {stage3_12[6]}
   );
   gpc1_1 gpc771 (
      {stage2_13[16]},
      {stage3_13[7]}
   );
   gpc1_1 gpc772 (
      {stage2_13[17]},
      {stage3_13[8]}
   );
   gpc1_1 gpc773 (
      {stage2_14[12]},
      {stage3_14[7]}
   );
   gpc1_1 gpc774 (
      {stage2_17[13]},
      {stage3_17[7]}
   );
   gpc1_1 gpc775 (
      {stage2_19[10]},
      {stage3_19[7]}
   );
   gpc1_1 gpc776 (
      {stage2_19[11]},
      {stage3_19[8]}
   );
   gpc1_1 gpc777 (
      {stage2_19[12]},
      {stage3_19[9]}
   );
   gpc1_1 gpc778 (
      {stage2_19[13]},
      {stage3_19[10]}
   );
   gpc1_1 gpc779 (
      {stage2_19[14]},
      {stage3_19[11]}
   );
   gpc1_1 gpc780 (
      {stage2_19[15]},
      {stage3_19[12]}
   );
   gpc1_1 gpc781 (
      {stage2_21[11]},
      {stage3_21[7]}
   );
   gpc1_1 gpc782 (
      {stage2_21[12]},
      {stage3_21[8]}
   );
   gpc1_1 gpc783 (
      {stage2_22[16]},
      {stage3_22[9]}
   );
   gpc1_1 gpc784 (
      {stage2_22[17]},
      {stage3_22[10]}
   );
   gpc1_1 gpc785 (
      {stage2_23[15]},
      {stage3_23[5]}
   );
   gpc1_1 gpc786 (
      {stage2_23[16]},
      {stage3_23[6]}
   );
   gpc1_1 gpc787 (
      {stage2_24[23]},
      {stage3_24[6]}
   );
   gpc1_1 gpc788 (
      {stage2_31[18]},
      {stage3_31[5]}
   );
   gpc1_1 gpc789 (
      {stage2_31[19]},
      {stage3_31[6]}
   );
   gpc1_1 gpc790 (
      {stage2_31[20]},
      {stage3_31[7]}
   );
   gpc1_1 gpc791 (
      {stage2_31[21]},
      {stage3_31[8]}
   );
   gpc1_1 gpc792 (
      {stage2_32[0]},
      {stage3_32[5]}
   );
   gpc1_1 gpc793 (
      {stage2_32[1]},
      {stage3_32[6]}
   );
   gpc1_1 gpc794 (
      {stage2_32[2]},
      {stage3_32[7]}
   );
   gpc1_1 gpc795 (
      {stage2_32[3]},
      {stage3_32[8]}
   );
   gpc1_1 gpc796 (
      {stage2_32[4]},
      {stage3_32[9]}
   );
   gpc1_1 gpc797 (
      {stage2_32[5]},
      {stage3_32[10]}
   );
   gpc1_1 gpc798 (
      {stage2_32[6]},
      {stage3_32[11]}
   );
   gpc1_1 gpc799 (
      {stage2_32[7]},
      {stage3_32[12]}
   );
   gpc1_1 gpc800 (
      {stage2_33[5]},
      {stage3_33[4]}
   );
   gpc1_1 gpc801 (
      {stage2_33[6]},
      {stage3_33[5]}
   );
   gpc1_1 gpc802 (
      {stage2_33[7]},
      {stage3_33[6]}
   );
   gpc1_1 gpc803 (
      {stage2_34[3]},
      {stage3_34[1]}
   );
   gpc606_5 gpc804 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc805 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc2135_5 gpc806 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2]}
   );
   gpc606_5 gpc807 (
      {stage3_4[5], stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5], stage3_6[6]},
      {stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3]}
   );
   gpc2223_5 gpc808 (
      {stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[7], 1'b0},
      {stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1]},
      {stage4_9[0],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc809 (
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[2]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[3],stage4_7[3]}
   );
   gpc1163_5 gpc810 (
      {stage3_9[6], stage3_9[7], 1'b0},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_11[0]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1],stage4_9[2]}
   );
   gpc1163_5 gpc811 (
      {stage3_11[1], stage3_11[2], stage3_11[3]},
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[2]}
   );
   gpc615_5 gpc812 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[1]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc813 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc606_5 gpc814 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[2]}
   );
   gpc135_4 gpc815 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4]},
      {stage3_19[6], stage3_19[7], stage3_19[8]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[1],stage4_19[1],stage4_18[2]}
   );
   gpc615_5 gpc816 (
      {stage3_19[9], stage3_19[10], stage3_19[11], stage3_19[12], 1'b0},
      {stage3_20[1]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[2],stage4_19[2]}
   );
   gpc623_5 gpc817 (
      {stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[6], stage3_21[7]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[3],stage4_20[3]}
   );
   gpc1325_5 gpc818 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[0], stage3_23[1]},
      {stage3_24[0], stage3_24[1], stage3_24[2]},
      {stage3_25[0]},
      {stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[2],stage4_22[2]}
   );
   gpc615_5 gpc819 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[3]},
      {stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage4_27[0],stage4_26[1],stage4_25[1],stage4_24[2],stage4_23[3]}
   );
   gpc606_5 gpc820 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[2]}
   );
   gpc615_5 gpc821 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4]},
      {stage3_28[6]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[1],stage4_29[1],stage4_28[1],stage4_27[2]}
   );
   gpc623_5 gpc822 (
      {stage3_30[0], stage3_30[1], stage3_30[2]},
      {stage3_31[0], stage3_31[1]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[2]}
   );
   gpc623_5 gpc823 (
      {stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[2], stage3_31[3]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[1],stage4_32[1],stage4_31[2],stage4_30[3]}
   );
   gpc606_5 gpc824 (
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], 1'b0},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[2],stage4_32[2],stage4_31[3]}
   );
   gpc1_1 gpc825 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc826 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc827 (
      {stage3_3[6]},
      {stage4_3[2]}
   );
   gpc1_1 gpc828 (
      {stage3_4[11]},
      {stage4_4[4]}
   );
   gpc1_1 gpc829 (
      {stage3_7[9]},
      {stage4_7[4]}
   );
   gpc1_1 gpc830 (
      {stage3_7[10]},
      {stage4_7[5]}
   );
   gpc1_1 gpc831 (
      {stage3_8[3]},
      {stage4_8[4]}
   );
   gpc1_1 gpc832 (
      {stage3_13[6]},
      {stage4_13[3]}
   );
   gpc1_1 gpc833 (
      {stage3_13[7]},
      {stage4_13[4]}
   );
   gpc1_1 gpc834 (
      {stage3_13[8]},
      {stage4_13[5]}
   );
   gpc1_1 gpc835 (
      {stage3_14[7]},
      {stage4_14[3]}
   );
   gpc1_1 gpc836 (
      {stage3_17[6]},
      {stage4_17[3]}
   );
   gpc1_1 gpc837 (
      {stage3_17[7]},
      {stage4_17[4]}
   );
   gpc1_1 gpc838 (
      {stage3_18[5]},
      {stage4_18[3]}
   );
   gpc1_1 gpc839 (
      {stage3_18[6]},
      {stage4_18[4]}
   );
   gpc1_1 gpc840 (
      {stage3_18[7]},
      {stage4_18[5]}
   );
   gpc1_1 gpc841 (
      {stage3_21[8]},
      {stage4_21[4]}
   );
   gpc1_1 gpc842 (
      {stage3_24[4]},
      {stage4_24[3]}
   );
   gpc1_1 gpc843 (
      {stage3_24[5]},
      {stage4_24[4]}
   );
   gpc1_1 gpc844 (
      {stage3_24[6]},
      {stage4_24[5]}
   );
   gpc1_1 gpc845 (
      {stage3_25[7]},
      {stage4_25[2]}
   );
   gpc1_1 gpc846 (
      {stage3_25[8]},
      {stage4_25[3]}
   );
   gpc1_1 gpc847 (
      {stage3_26[6]},
      {stage4_26[3]}
   );
   gpc1_1 gpc848 (
      {stage3_26[7]},
      {stage4_26[4]}
   );
   gpc1_1 gpc849 (
      {stage3_29[6]},
      {stage4_29[2]}
   );
   gpc1_1 gpc850 (
      {stage3_29[7]},
      {stage4_29[3]}
   );
   gpc1_1 gpc851 (
      {stage3_29[8]},
      {stage4_29[4]}
   );
   gpc1_1 gpc852 (
      {stage3_32[12]},
      {stage4_32[3]}
   );
   gpc1_1 gpc853 (
      {stage3_33[6]},
      {stage4_33[3]}
   );
   gpc1_1 gpc854 (
      {stage3_34[0]},
      {stage4_34[3]}
   );
   gpc1_1 gpc855 (
      {stage3_34[1]},
      {stage4_34[4]}
   );
   gpc1_1 gpc856 (
      {stage3_35[0]},
      {stage4_35[1]}
   );
   gpc1_1 gpc857 (
      {stage3_36[0]},
      {stage4_36[0]}
   );
   gpc1_1 gpc858 (
      {stage3_37[0]},
      {stage4_37[0]}
   );
   gpc1423_5 gpc859 (
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0], stage4_3[1]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc1343_5 gpc860 (
      {stage4_5[1], stage4_5[2], stage4_5[3]},
      {stage4_6[0], stage4_6[1], stage4_6[2], 1'b0},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1]}
   );
   gpc1343_5 gpc861 (
      {stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1]}
   );
   gpc623_5 gpc862 (
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0], stage4_12[1]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[0],stage5_11[1]}
   );
   gpc135_4 gpc863 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc215_4 gpc864 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4]},
      {stage4_18[0]},
      {stage4_19[0], stage4_19[1]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[1]}
   );
   gpc615_5 gpc865 (
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[2]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], 1'b0, 1'b0},
      {stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[1]}
   );
   gpc135_4 gpc866 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0]},
      {stage5_24[0],stage5_23[0],stage5_22[1],stage5_21[1]}
   );
   gpc1163_5 gpc867 (
      {stage4_23[1], stage4_23[2], stage4_23[3]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_25[0]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[1]}
   );
   gpc1343_5 gpc868 (
      {stage4_25[1], stage4_25[2], stage4_25[3]},
      {stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4]},
      {stage4_27[0], stage4_27[1], stage4_27[2]},
      {stage4_28[0]},
      {stage5_29[0],stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1]}
   );
   gpc2135_5 gpc869 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4]},
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0]},
      {stage4_32[0], stage4_32[1]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[0],stage5_29[1]}
   );
   gpc623_5 gpc870 (
      {stage4_31[1], stage4_31[2], stage4_31[3]},
      {stage4_32[2], stage4_32[3]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], 1'b0, 1'b0},
      {stage5_35[0],stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1]}
   );
   gpc2135_5 gpc871 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[0], stage4_35[1], 1'b0},
      {stage4_36[0]},
      {stage4_37[0], 1'b0},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[1]}
   );
   gpc1_1 gpc872 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc873 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc874 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc875 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc876 (
      {stage4_3[2]},
      {stage5_3[1]}
   );
   gpc1_1 gpc877 (
      {stage4_4[4]},
      {stage5_4[1]}
   );
   gpc1_1 gpc878 (
      {stage4_10[1]},
      {stage5_10[1]}
   );
   gpc1_1 gpc879 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc880 (
      {stage4_28[1]},
      {stage5_28[1]}
   );
   gpc1_1 gpc881 (
      {stage4_30[3]},
      {stage5_30[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor_CLA64_32 compressor_CLA64_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h747cf5c1a18c8da11efd87cb84eb22fef4fed272f578ed74426efd8cbe56bce49bc4e499e62ac551dba0e6bcb565e67db232e4630adbb9815d4cda810fdbbca39e412d05370ecc09818cc71e01c76a55967f5b8535f1a10ccad062ef1445f5ce1c11d607b5bc79de4917df49c98726057f48f39b970ce35e304ca8f25c59b3aa6948fb5d1c50d0ffab01db1e1a7a461190096825ddee3f58298f824ffad2c86cae3e71062ffb24bf09cc63b1a8c7ca0811b917b8d698f654df0046c5d1ffaba26bdd82c67e6699e2b2911ad300b090b50c9a8e4db0128775bac0fb9c69f7f21175256fe3e0ab77fee3d568c5af46885d712a73861f1cc36cc29f1479d45c990;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hab8becedd3f9f531b4bd36fbbf453f173b582281a0c2a4d67ef7101efb2f89ae9cce36980dcba11e154528be4bd4912615cd3ab0f8fb1ce3d39ac3379de33b0d79957a61679d64836662c3b9c9828302c869fd64be9191950dbeecff3456f7ddd85da5715f97f15853922e3cdb0b904c07e37a1e6798c176de88eb53331dce28077f89f544e994ab33db289199ee51a1e0acb0e844ebf2c67d0ab93526166112e25792f7131449ad65a974e61c68dcab542b65f722e5fe1c107494326223f3a8e1fba6d7f51b6239258deaf8c0c4efc8d6bc34a0b62f0184bad922b34fd66b70da3e93f5bad6628c89899a523e3b73427d6a8a6db595f5dcdfd7a6e4d2698bf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h42c9c7d8ac401ae5374344111d4e4a9552d456dcee3dbda767d17179d736255cb5a864667be24341d7aedc9fa4021d2a00543b89641a882408dd3b9c60e6e18b411f4e9eb46abe9bc1cdb2b25febbbfcad620365da3d42eb4a0879157299cd8398bb516604b9062b9aa4e8eeec8368d745865732a64275d488a41afacbd7988d079a078600511721203f23b48df934ddc18c60aa24798efe099b63b9d669abfd00102fc50e37fab32ffa9aee0190ff873c9da83cb1aed3729471a7c92e734224edb324ae53d6a8a6823d86c83fce35fd755b9b08e3ce7ea65ae96f7d5223ba73081d178bc156dffb94fa0b143387516969649c80f1403b1f651f81b389dfa675;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc20d9035c21e1afd482c1b44d84606ba1fcfd7b1f268257e9356cc2931421dae49eee367d3c2bff0a3903be24b12c2e14b4b53d20e0006eb98e44c80a40fbde7026876d0b06ace67fa85910147b4a3f187275473415ecf39c79f129e9f2365a30f8a90a8f84587d353de3c9776db562900948000aad4cb3b31d2482bee73481f67fd3c97c134d3aaf85a03aa272c0da74fda81bb9b7255ab4f9ff030d228818519dc6e6fc03ed416d22f2676d84b4ddc406e9bcfc450bff3326f8fe01932ac9cfd2f83bf7602efe048a1ae03c1eb5569123778316986d158b63b51627cec32996c8edeb2db60b64c693cd2bb8c171b24c647ac58cafd14eac5fb61f9745c7a39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he4f5e75401658b570932b60a434e4bf20fc3aae76b85e6dda7ac395654bcdc8c762e64ed55f21c291ea38838efc10f669d7666b8844a9f3c244403beadb1126ab7f116b3ebf82e6af542458ebe9f5c8c1b3dbf80f867b1251d2e7759a8c96bfb6c3b60370130eed1abd167fcdb0f697e9056318cff8a64d5b7d05774fe830a66475caf043d13954b45f21b4b066013d264bdaf571d43b76fcc5d82c3dcfe1e7ebce49b07b77aacb376e1aed9b0c593dabb84a9218e1861d040e1972b57c8b0f7b36ad757486bd3f0901e8efafd571b62591f23172bd906685b84fc2ee10c8931640c16f58c67a81d7f0229a934a2e1de087a9e43401366249bfae049a2c0673;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfc746384690c9177965742fccf95c7462da6cf3e3a0b944ca525b3b9c5ccb8469340c5bce55bbeb9c7b5af6f11c8fb8b1af3b5dd40d48adecd342133491c0ce8e22072c91446ebbc8ddaa3b1d0cb09d705fa44c81f77d837a91f1b46b9cbcdef4b5378aa16feae5725914a6f20e3be8fdf9c0c3172947fbe8beb454d275693eb847fc5d2738b48de8328d430b62db3bbfadce186cd5c670a5f33c1a8fed2fe5fc64c29092ca3b2cfa4bc3e814bc3214ec4edfd107ae5683e08eb03587b4100aa16884f0b43571cbfd6d5317c0825a82c760d81ffadbd89f4a3759653a9d7d1475d48051f99c01e6a228e2e528242e556c52ea70b82f55d604a88dc4ccce6bc99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbad0a5bb186914b19bebdb7fd5d77a79ccc92e19ebc76cd5cfa25295d4b0a1b5b8e837bc767837d68f30726e84b444b7682f01c2bc1468694f8b97df25d765247ed7f5c0201a507f515c31f540d1416c5cd13dd5d4d1f980848b78b51e3ed7757a854edc08b51f2af51036352df6b1c64308f42d5bfc3c1f5152d414a258396889c3b207f63542f93e4e5c78303b0cd67f13992ad15cbcd60263ef0c5c397f03e4076e731f12685489576b6337259b825e90758f9c436c38bd2301e14819de5473d7645ce500148e6725c785bb57fd8863d710f479705b8309299a9affa034fdfc77a5309df7a9d089f25f9892f0ec11edf1f2903893c88b3fb08c83440c1ba6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h229a60f924b2c44e9796e4f7386988c33eb40b0c0af60426d36d76f84f33da0337851f758b4bfe1d4519c164194eabd2d52ae03b8795927cf396909aa1b839f90bdec344cddeae6b82f2c42e8da7a63fd2eccabf6d0b18ed4ff85a094953d416481f7a303d1610cbec06ee4ec572dd958b2b1468468a304ac437ce78b406db838dbaadd4f767265996149b1eeb595d04dc8c6aa3956fbaca2e787d426f3e3fbf0ff004c098493296d256e9594de9aabbe81f0228f9519c5d27b9b1a374d604db1f4a9ac11bc492f94068eaec7ae46f66ae1c92bafc0db0f01d02a9393d0c63c4e91d293d006a76e8ead1efe292903e15dd9f964c5337cbf25f69e771f7f24c33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4fa03979cd95c6eb97ecab6c6975fe8a693ed3f177369b72984fb56c02557a562833b04d474e643f3c5631a32658d167043dcff5f5604918210d2350f1bb2c5c42fc0ada335733c517bbd990514900c7508df464769c2604d1ab04b78d67e9b4618e77d3ac82f28cc8d1121028a420897c8d8668b81bad779311868e8684ad12562a6261b30d3b5c4cb84c4d2860ce0958cfbb2cb462bc5ec2170f6eae25c581d448393b8913c2e75958b9f747b5f58654ed4a16aafdeeff5af4657bb339eabe1bba3efef7ef42e4d57fb88193e8fee1780ac46adbedbc730b2f0582c79e957bd36cc82af729c91b4a7232688bf883d68c52767933f71dfdce5f0d84565dad41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffefbfcf380aa0dee501641b7eab117903bf1f8f1dddbc8eac7ebad759a76bb679579629044b7aeb057cb55c3ad7c8e65f34c0f056a957708b6ff30ae4bc5176620149fee7594e5832b3067e7e5e842c1947f196d0ba3f7b59c8384834ef271138d8b293648830ac847dbf43cc2cc7dc6d09518c2f7c8c12afbf34ed377eb277f28033b90421f56053e6ace463433105202a8b5349355eef054993d26ec76c5b99f4408e26c9223afc42c5e4bfea013442def148d6725f3da86ac58de07e97746aec3d1bf01ac5002318d966a8dfd7802d48f72cef89c9d6e299db06321cf96b2078df1bdf3b48168e4010565567dfeb06b9c554e126a87cd91d0c993e63888b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfad581f44d35535ca91cc851ee969ed54e0864e57d05f8d8e8677c566b940da23f668b3bc8e20f09589c02121506b67b907de719b105901e940ebe3b4bd57b481915ef885ebc97eee4f37d23a57696edd5a42273fdfc00604be45b61c2ab9e30433208c1f53ce14da4d22661d328ad0b7247ed837a4816f7ee92277d2f0f75fa2f3d59ef45110bd95dcada54dcc7425457dd8c36f9db39389af80274da4f11c95b80feadcd073fe0f4fe17ec44485fe9578754265ae7894923a503b79bcec3f39e47fbdd8aeafaba31afe3ab76d8b42fc5e018ddeff78a49b5066aa042e89e8e24780c78739d010ec50f85639025a9b4c3b26a8e06c85858629ec7ddd0149779;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h466df0be8ffa336258970027b2a1e27b882a1c475883c519c4de23e2306c0b411ad93ae7bc165dc7a0c06704771bac2260a16edb89c2ae98fd1bc46a2bfacfe351453217461da79afd9d184f59ba0364552c48595ca3890740ed8ed0024bb476f0492616d2943941049ce4e341d1eea53ed4da956d615595d980b0297b236ff7189d0bbc58f7739f8adede16ed919d695ea5fad426f18f7864428c361167ef6b6eaea4bb600bcdfbdd4fe424188c13195759521da8cac02e605324701f24e401869eeb833f02c194397cd9d7cfc48148e06bf0e20d5b49fa5a4340b0759553c9205dda6a89976789051d953f97cecf98b3e25ca331641eae350efeda5f55d7a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h85a0dc43be0736954d2156d1be4e563cba921ae38721993558c29f2c725304b4dbde5d7c052fb97ecda331c1458ba1199b0b8050185390e7a0dcc1d7eae4405f0e9a0f884a0f5a9c90a5cdefbc71ca26efabc8acd261d5cf8da69be9c6512fd6cd77baaf614d9d12b7bad83b9234ec05a61ce5257fee456c2f413b579ba669bbca56f14d8f7d130becf4007ec498b1fa3ee8b12e6965c1dbc050df4f657b31ae92bab65591718ec8e50a682f3bc115d5d2b55ab8b2b4a4d1a7e2f6a16a5ba14f4a19f744c4b53288343c6f112f1456a2f4e0b8997c789678b9182bd89827ce38344014adea00b4e404ec4970fc657ac25ce9140362400f4a1aabda496ed5298c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hab143f66b106a39a54152f1a38e0289577a16d3216ae2c49d067dc4f76f4d773a52c8b5b8eea08fbd0afaaec42bb393241b17ac4ebe139e6b843544762945fc3c1c51455d2258c43a0b8f6f1bfa048678a259997f09ce085836a2f84dd7853fdee4ed3cb3b2fca798c04c3d57f29b87bab8cad52af63b9c6480c3fe8a7bd0831c7b5b590f7634c94124c56dc3107ade55f5056797237ec2ce52fa10e95bf15577087344b9580b9a3cd399b69e9669b3aab67929cad8f78b4dd6fb2333b7f9055e85210716181649738be1866d7cd979eea24598f8050c3dff09134a30071464d4d76b973bd47b8a6e0c45120aa4c82a0a07c7bd6d34eeda98ad3b3280c68ca89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9c8c24d6acec40a186b446dbe184352eb6920a76610f12271f96271430ff164939415c2689045786db831a97fdd1b50358bdc4565f5a45ac1e6a0a2061f3b5c488a98372d56819c461b61ad89f159285c7e993606da2859522eb33862fe1c70b2e26fc28ff00c6427072d378404a0b774229340d4102bd35fe762a8271f4ef128b5dbaefd2161373f2613285ae8471bd43a8b0be576ff7a46ba47e749b4568734f877e10e58987976218729619c70f77d98d952555abac3d02e69503b9443859ce254427c238e501a7f8280b79231a608777712e823a4e6c60c176b2ef3919e195f873dd1dbcba0b8d6d8a26facec41de0ba961cad077e2f017e691f74552e72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf53d1c96377e4fa143681a4edb39f196360e25d8fde72e6b8bcd32677dde34cb067057423e68542d10a8e2cab1f54f16cb410f4705469ff72ab3c63a6d877901cc15d8c81d56ca325c55e2c3cc6caf39834b12f7cae704e6317715ac8bf81feef466881f3028a5bdef80339633135c86043c8885f6d3a64ed00bc12dfaca1d108cc079a42bc3b5ebc731ec0bdef42298847b9608351909ef976e5ea9b241cd456729b4eadee2a938d9abdb1ecaa3560d8deaea8741723a6da176e2f30d01f314bed683f57e52150f34ab74dfe560ccc5bbb47df767dfc93abeb6e2976555d142aaf5ceedabd379c09b450ad8c784fbfacc817a5ab9991d81030f8f58e9b82686;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1a4cc7d4a890c3822e90d9010a57658328c48eb999ea39319627a1a59337e878878cc7ed637b44981351a1e3c3e38df0684254a145e42135652c008c24d2855e812cafa5640c0ad5c6c6f9c32d35012697097e9fcc11271c25c27816356d8eddb77d9c546e6581897266972e0bece98ce2f9f3df6c7f0549d0f7a36a53c424dabcdc678aec00a2da901908d7a160e5f19e32d95930e9b16f14a1cbf23fa618ec73198ae40052f5f00c3900741c475b187024f8491723e43320b14096ba4ff4e92f630887b69fa878c05a9f4f92d8b3157dd7f285ad033a69e1cd29f15ae034e21e07576cf328a592bec8401e2d7540e7b3f6c25a017c33acaad2afa5f92d4bef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h73065dcd70e8bbe6c24ecfa7d33e7cb943c774392cf9491bce027f4dbba0e2cef760a20fa968b0497f67ca962e5f7c9b5ab33bd83150d119abcadc8b8487fa718ab7bebab4e46b76bb4f4ac572c9d7cbca846aacd4d27d5a368367d28e0c3ddcd21910945719efccce541797472d11bb57ba5e403e9c7ece3236794343aad1fa72ebc4dedf658b54297777f9f4dbe8b18b9428bca282651ae44745541418845d26188beaa8db61c8c14a034e09098eb077de15dd60d8a5dee3981d5bedae04b4d15c8c70fdeef28670cd44e4f11ccde434f4789a2059b5d13d9df0788563a1bc46fde8efde0bec6cb233e9b8da91b59ac51eb13fdb03d331f689bd412324865f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36c3bbf3ee89e0a19a4c2ed95f735984e3e11da277bedc3e832ad87ff5eca35d6e60416a0e86cd8df01974823fbfc5a6b0c2bef66b3dcdf3f9a986e4eac50a2cc0003bd95e1f06d8e5133b99d7e0a12fdfaf05587f6b560b22e45465ee64264f7025731868dd129522a596e3de0b26700b99d0c5235b418dfd9dfbfc1ad744a7c15a1c602961e3c075f31b5db2f1838457942bc69b082d98f73586591be943dbddc782a666c1cd9f3bf74fdded883e43cf6611e5f3c1dfc2dc4b08fefb8e106fddba7bb91b3fcc658b925a616127a34810e054bbf320cbd83381fa63f547a59dcbc7260312c9bd737d2bd35c81fc596062a4e189898bf634def7c9017add70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h285f0bd895943ed6da077c879d6f1aaa20503239b2efb5695a0885e8d62f4d9842331e73a6014a65d763a62d9f301f87eb7b9cbc28026b52d538a9dbc8d768fd04bbed1ac8759038b1871a3c471bc507b313af3e2dc29cb834f0c0efd737868fca439c79474724446515ed283ce206792772ce24e76fad621e7bfcb8a6cd6649a3b7b8faec3d5c98deda181f897f56fdaecc225944b24ca08366bb8a12d7a383d64103994f1de243b450721df7069031c60b0ec8115a800aca56d1f2db5023a947a62e5425276423d7e185b57a9266fd47dc4d2ffbe46b8de578687ad83fd550b91c12167c07b1d3ef5c1eded44381197d29bccdf2fc8877f18ef84b5227e556;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he92d9c277b5ac00d914e206276b12a267f060ab0751ecababe6f4493f15465fa23b6401a4201792e54f72fd0a3daab5b574585e0e2a465d0a1ad0e17850b8e59f79f8c19abc9dff97ba8dfaff5c80f56fd0665e8fb5bbf29bc7ee26ffbbf25c8890bd3832b87d65c3f32a124fc269e5af86bb8e84dd4af34e33d058e6ea2fa024edbf09a04eb16f83527785dc22013408ff70d42e6eeba4a915ee73a5c41ad282c2fe9643f1cf23f84591dbd6dbdc2305bd09856e7dc2a085e367ce956593b32b2999782e4c170109a73bf3a20e858a53e29ea15ae96bdad285eae2aeed637bef97673cb685d34efabba61e2f289bc818552ef14d40111fb9afbb475aef16c6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h63a15b126ae0c2a4a53ec5773ddf7827c794e532f7843b606e44e2e23c9a042d86779f495bc416c85c3cbc69d0840efe2c07c2ee84e9733e7aaca27d92de04575630c270258cb4ed105b056d53bfa1535a04c1c626af40cbe6501623037a73f11ec11d2995278d00da9111a462d96b102bcd23651d23d36409b3d59168d40e9830be995c70d8db0f06522ea844957dd47ae31158b5af0808f8f0d507fb6ba67e800b36bc513c7dfb5bbfc8c4e61e24aad6d399450a185fef90ccf4e00cb62f5b1211d2ab4a01a973642abdde8a395b98434c1f6c98957c4414a4e03d79c7e26f97bdfdb8c2e08fa73e5f113b1033d1b2f313b6fa16937f55871d86d880b2f6ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h268a293d601e6a61e5f3ca36553cb2ca18ddb4d0802b2257c2cf8477f5f9af333e36956eacbff533a12b7f3bc4a60a5a2ae7e905d498999e6cd736acdacad19d076933f4bd6df70f6b8ebce584529ccb385f9fa4fcb2423cab3af8597213808ea57a80ccb52efd426eb370478b7a2e723018b87555c64da4b3fcbdaec4622e996466bedd1dbcbb18e841333a7e952f457fdacab07e549bf3856ad71137fe6ff40b0d94dd6499765f034b91cc4813826ef6f7f3735a496146f83ebf892baf8d6674a15ae00e1968f3b6cc1c2b34d34d69a79fa3d99b770632a9a5cc3ad0a8441842feeed445685ddd54e662cbee75ad65862f032f673d3e2df5cbfbf570968812;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha3b46309d3a5c3ccd8798470ca8d4ec87d6f5090f54193cefc3ad3295c69f776cdc7ad1cf22c240ca5a83fa3d7c59ee7ca361525378e725b7e61513b07df24895e9be4b5a874104e6c5400e55c06b4b5ee21c372eee6e11229707c0ca9ce30252e899fdd88aec3830c50c45d5d22594c3353fdfaa6693861d7680eeb2ecc76b1fc3e03b7665881eed2a7e23269059cd77b98deb49a5fef3cf2ce7f4d28df4c7b898607e30b340f9b5bd6b5b40a50ffa73752d2c99dfc197129fc090378bd209ed1ea5f24fa662fd9eea2d170f2ed5d47243ef38c6c7d9ee55ef739b2dc1ac28c291fca1b34551a926e2df5d303171cc418a87aa3aad1d9af569a71b28e45f8d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h706d17e9df5f40b5751538f75053924cfadeded715bcd6c03ec12f07de22e6b365379d767e1416e50d234191dfe9d7c87489925709a13c6bce82ca3095b95c39df5c4daca4d4d7d996e61dba93d94e869ba7e556ccf7176568bca664c736b266c8e412821b960ac3b19d73bce648911cc1f39600234249965aa8f66dfdc38e8a885988fce4ee089115cfefdc669aa51a20054736237efbcb49e13cc09d0d8d7f1324f2adfd323bece9e9ac4b865658b73fa5ccc848268a927f854979b61d682ae3b3e427e24f3894f1166d3088254b3b74c3aa2ce06bbf96e5c6e5c8010fcd287bb791b201b41dec67b9c7d3440242699011dea3b7d7c6124a99d8a2f37704b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1d04380b264dbc6a2d974d81b6fe43e6037f6615b561e6c93b3bbf9d2902dbd87a5525d210e28b6c66e39a1e8e697ca17022535e8e4ed0884085484430da9ef1850f6384a08832160f79276d0044edca81ad81a50b6aa1191c75689b3c989d2bed874a17c28222ec3ddba1d2c358846cad148f7ad799817d84c8a8c3011cb930e81683d32dc54e36bea7e800e0fc1f35a378ef00d96134608c55ccc3d939ed3d0d4d6f56e88a404fd24a2cf15d74e8b84562e88ad6d163c6cf2d82f5f34b4100413fc1d369df6905076af7e68d2a381ad55b55ff63a66c85a1a3c1d997f014fe43357c1bb4211537c2fd1e1a5f356c3fa9a473cb9dd7beb0612b9045024835fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7c8eb784324668cce374c5589de4fb1479f720bb3c2bffcbda622c9034dce4b36afbbc4ae7e3d50cc8637bb26acbb1b42a5d8926f22c74fc8bfd2f61a9dd4cbd38febb95cec734ac9799fae64ee5d48c44351e6d8251a7da4091ec94780b193a9799ed0e3cdc8f93828dceae17732ebfb2b9bad44311e560073fd006d3260d836df73937fce4243194fb75a118a4a56eb92d38b7ad06f0e7435e253b53abf065fa1dc41e59d95f453ac7ccfb3cbc26ba51195a5d85b4fa35431789a43175dee0f1c52036ac4295d79954940746bd3bcd93eaf2f82991328b7aace596514205934a461c667213a89b7dc22cfa61b9c9ce932a1861135faa3d66d826dca29ab6d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf6e0df6191ea76817d10e3c43cdf5ace3bcd4a8c99321e2cb8798e588cfb5545c8050da9b23ff4e06585424498d5adfbc574524c4b75f26a4263fdc6659a31469cb4b6df693ef04cb523b1eeda2f6d5931cd6efcef73fed62591c6c3ded609e8557495ab855c67ed5e05b31349cc2385e5bc58042363df04af1d57cf8a8426d31c4b240f7241075ec52c614e448e34d694cbc539172b00fc4e46dc95b5d7386de78353043dee519533b3c51fdf4ac6d3f2086ceb55632ae5fbc62792e8412223d5ad316b77cd2dac4e0ee280fee7e98aa5dd3a806d01aaa086a70c5a3fe98f931826bed89ab9b91c3d4b28fcc245ae3053e917ec23e8c409c580865963eb5550;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha6f8b6fa05c78ed54a4f9dcdfc49211006b093d0ac105ab7787bd115f2f95602113594616df52568bca02a67a682a3d7e4caf0d861fefb206eb2716ef134468ddf40a39f99079acaa8e2955ae9aca2039c3fa762e19839c0b0de928cc6f58f8d898e3d81262dce9c2740386781b2d8be7cf0f5831f1ed5554dac56d0d2d841669bbde0dee7d10400cfb2bf9141d97155237ed8da24add2d509d77a90b456d07234398d737183308fde4ff6ced30a28be2b8c391de9f3f001fdbf1779d56399ed933747b6c3941e13a2b7869b10bf033e2f0265d63f2a8b01ce4e7b14961878cdf5bcea509d9710eb37650286c799cbb55a73563738e78096379da2077608cb5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha5cebc9ddb35ac205e5f27b32b563092c5a036718bca47bf1886bf16944d84830071c7e070ff15ef1694f30ac2fbccb107e1039467bd3e2da2f8924fc336524b8eff1e7b754eae904631eb236797cb54d890011040f443e725d4cc3908dc905d52a113909023178eb1245a922b46dcb2689b6cf5458eb4dcbe8f8226f44056b6954bd7e35b7abcd533808f0ff1e0fb6c5340c8d0b2e0ddebc62d203bad0a31fe4779d864c6ca16d20fa412ed71f293ed652b01bb2a4a800b858768eeef6d7a9aebf241b92990f573386ded0d23aa5d982bb88be63ce243d3289b6fa26a5ace46d931ac7b7e71fec91869e4dde4eca515914b65f1b688b05e48b9b6accf508587;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5c56b0a8d4acd546f4f1c97734f009618da08f418b7b66ec683e6c381391413ece0b875942129015036208c47e46155e27eac2871330c99d5f6e1646baf23713987fe9cafd15bd617adfed8f343d494d2e1cdfa14a18a35d54264d457ff5229d3a2f808f8dce0e31076fc652a351c63779cde74b5975e7ea22d068bb2560cbdbbc502e9f73f6558abce7f79197ea9bb2dae2cffa77c5c842e4582f2359cbae34d65e1951ba92c7dda23469321aa9910f23548f77d4c2632d9447dc349cec5400cb1457230dc1e06d1ca74ddf90593014c751b79f0a2692a4d3997d586ca5060ee07c5f78ab7205453b652b7e2a9ac795d2f901c7a30da62a6fc848ced3eef2d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1fb9a27d4e8828d085b2e088d32ef7a9df280a72ac49fcf3efcdf76332a974e60c825f85f21604c5b32965495e56a87495b49ecb79ce180bc80d16d1ce2f51fce82a2c9e22bf7af09b98461bf3edd85682e53fa3f11eb1d55c2336dd0a3a4bfcef5f442732837b8b607ffdf81d95f56b4b30808b5be2c768b7ff560b203b63b692cb5ee93cdb09514d3f295e0d43245cfea052874805c73b589a8bae5bbd0c3bf3626fc09924c5524c9b3a59eff3395527d64de777b85394493dbc9b9703325e74037fe2faeff7f0ed71a3a8537a90928971a55ec5e422556308f57191d7fc816489bba1b9f2939dbe9b9248a2219befeb83d79024b41c9074a3268a0ef8b7a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbf4e4dae55f2af8cb068d8f766dfbaef31e6d1d76f234ab85c9282dcdcb0638f9f6fbfed8aaafa843e122491cb4bebd4c40d2e41cd413db5a7dd6e1aa6d00a71cb6d47e3351f633275634d155e3a290a5640ea9ee665fc2dbe79a5fc1a4f2108a55a0904cd469a386d60a8833dcd582c1b44605dc4f0f0ee0fa686f000b945e616f00b882030e4c2d4af7643afb922e09c880fcf5408ba48562f66d225d71720bd8e93beb8387c809acca2891bea40f6ad270215b0a66595d4c130dfeae8f4655adca05902313e4250ac1ae703271f5d895fe8c0f1792071280c2f0481b44fb7385c42f07bcb017270da0ecbf5f062cc50ed113b9158f911312f2fb81676be77;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcc6157084dbe5207941cb734e60bb7a4e1eb23bf83f002b9d30f4f0b4ac12b8d603e707ae1fc6b0ec06cf688a9322a12df30ce201b8d7cde04bce81c1e73a496cea0bd2132912f1b247513a92f1ab749665ec735796a5f8b751b6719b16ec68e5c8a7dff0d624db8875906671faf46f94e026d1b89906d0cda419ae25e03f8540b17452fbbf9d961934452b44d0113b2435cbcb616be9e3932ffa3a59ffd225322bb748d7e3946ca88a6170903f03298b38098cdb027909ebcada82e303c04e2f405e36cbd8b6a6b5be3b7bfe5a52ee5eb018d6f05b79e257401d87bba0c77c9b8e6ffcb2ffd1a122dcb32b1c412cef237d5c948605ef12e534e1d1267e12b4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc8070cafaf5c0b2db4b911adaf56cc16e1fe79d0363a50eef51b7a6de5f79152b6d00d2e36a21104fd73484747dddc9b57afcef896d3075bac0fc5dccc40973656c750326156a5661e608d4f93c101c033a957e87ec147b8c808a6c733e1377b7d215b6987cb9de2171c0e865e61c3eeb628091e3237e631b7ab52a58e4dab6c53aba4a805507b9530d41e887892dfb7771134e479a52bb52e4e15dd4cb129e6ba3ad8febe76b276b883706e705158a582bb918ddebc831aae6a22a2851aaf5844d170664ed827ff18f4dac68498e59c44ffbc616a146e83490b3a3471ab0903b80b8d42678b6b05f397d92d9fe79631c26f7c8d725fe8ec167c705b31d9b193;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcc51ae6b295dbd57922aff7b642c8f57483e4b8396b7b6a2ac651d9bd1a33e0e84f9359d1facfc6294cefc208dd67c4699b407c056f732ba0d505c8e5f0eeffdd3f04165a901601899399e9903d4cbf2ba52bd7c283af7c379c674aaa407a72ad20a799b4ebc0682101aa49a723d5dfdeb2991ef7661e2e6ce166278c5e4ee55c8c8cb191c9607418f9302196f799aee076b6dfeba9a32ee608fb5f8e3614c968ed9f06aa6d13fb983b13a59157eeedaf49e231be60e4ce646b5a36ef3072535d142eb297e00d0925a375e318652f14ea9217dc615dd431d15ca990d7653c5001bee8d4eb858c8eb9331ae03d37bce3e1ed17577d586b2c5e692a9699933d1cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb41054ed37c82289dcecdd1167336a10caf3bb3471b054f760f2a7966e6c4f22d42b0eba7fa9f3f2ffb749dca1aecca826cbe90e0ba0f9d1362a0d2ddb2c04f2f1be5c557ff4b018961234dcd954dba187bd15694711ccfef82aa5d8d19b33c6dfcd02e56f7a2d818f488f0be7de43e88287f088cf470d4f1319466cb933edfd2d6d00259f2c8049958d672f20d554ab9586ef4f32dd167c31383aacd4c2834f387f25ca51bbecdc1866107f74c469081099cc6a307495249ac3ee2c80cbaa9288338d2b01b7668b7961fb57c15e39a81f3ffd6169eeb2143f98a18660cbd2f1dc1ebd8040a36b32b51dd76f0686b35c3404c0217f6c705d12cf04ffd4cab561;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd01fe3e86b7fa2d12d299272e71078f007f984a5305c4c020e275d92387c94a5fa580f20663a3485c1cf767eb97484f4b7ae17e42e8df8a94cfaf7b5df6bbbf1710f2c6ad2f3ff9d763384b1bb29f8a0c0b7c0d49e2314d86f2af844122c9b819c4559f56559806027f2f838572f96b8abb1c9ea21805975fa8210d1f82583ab60f94729fa2a27f5a71c22e20cb46a0d18257d7a3fbdd92d6e7185ebdb4833cfacac6ddf38bc5b1e49d64c3fd26cf9fc8e6c80eb44fd9627572136087cb11cd71f2cd3d813d21c0a52f2bb3941ee8761a3174d46d066052aca86970e499e6b58e7855e73a40b7ece72843e89fc68ac2651922570b2ff1dbfedc7163aa9fdc0ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1a42a61494cca4226861e4ea3c5e5e41d23df7080aca7fab8b122fe018242e16d8d3198142b434e083c8bf8ec163955f4cdbd16a240589d580c359582dc16662ca808cfce227da6a296d263a73c9a2051eff40807ca4063188e4bcc40ab7f7417916da000070bf98d7bd6fcb68025165059f3699345bd41e2103894f91d720fe76ec5cc3512e9e359e85e8ceef4f1279e532767948477ad51d1693fa5eec156a095fc244cb1c55c415e9a741ccf9112ef4db3ba3974d294009870b393d649b8e1757dfa2cf4c83e02d5dec7fe4af974d59cadb69852bccd8b8812b6aacb0ec5db972acbf87c5795bb407e1f0a526d571b081d7a1432002a573d6e4440b050c6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9275f6e8bae14f1050124dba57d714b488e13f9de321857773702e7c60a7143acea78431b4be825372c868ff5f2b22576ddbbc8069392952c546aa1eee82e59a6ea48aea91873d3ecae2c1e923e7a260aacd2b8944e5fed0c9e90d67c9ae388fba77f8debe40c3e1c0d205af1ec56c7d2a717b3a30299ef4b75042556a99ad65abd8fe688a37cebd763623fb18af607ef58f40171580685e6fb55b51eae86408df748fdac1fd60c2af594880eea4a654b8c1068e3ffd3dc8b4805b0b8dda1eefdf5bc7df9a5d67490e1c7b57b7509bd9e2055ecc220aeba5a8198d1e7f171b89cd9b019b687e085975d1bcff8840696ac2e6f8ace208d4ff25845566862e5334;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'habc35c6bb6460271e57e46ca2dae580a31d2df4a9426efecf88fef3cc285e9987821c344d711b1452f76a34f3193aecff1116229ff9311c037e253caa97d5b3b10eb6be0942ac8344a7b3320875ebbb052e8feaa234dc1a6f25fd4624421e634aa342631349f1935887b3a9629a0b567b238df5c9af9aa586d16bdb31707f1777faa6dd7566778f93124a9cf0af9f53625ac0dc59dc85635519e7cd1848929f048edaa7aa0eb1fd6cefa53bf0e050eb0e54640492641bedfd1dc3e6ddbb9dd1e135fc824e2c20e03aa0fa84ab900f746904550dfc9e07f9606affcba9d8457584af24dad01580eaa4cfe2e518649758a743c3d2c893417c1f4308db4aa0010b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8eef40405ca68312c36c4f72e7de9d9006224b803ce986d1267bb16b465dbfe6ca78765916c85e011051a9d6d9ea1885dfb49b3866e1c28654f44e233315f6a36937156d48bf375f32d0d432d2ed7274ac8873b16d16567aff48c7d16bdc972d83c193fe9054500a1a476352238872a4eaf0b5423bfcbced73397560ef5884dc88e875a8b969ff60a9010baf6064bd81df3898284db85ab72d67d60960f7f1d6d71abed437e025875e96bd7f30ddc770d12ebdad068ad3991b1b87c120f9aa62a31e421adc06df35533361da9be17dd3732a2924cb46ee0883601ab789d0132d32eb2358e9da2cd1ac2311784323a060ce3ea02c472cb98d504be9e281867911;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hde3047ac65d8af824aedf86773a12ae1f409ad41367a8e7d63ea1d5b0832b922f62d823030d4f977fcf30e6609542da491dcbb13ee0633fee3684bdcf31eeac2f8944fefc10e8928b1025b56ded2633084600de2fec032bec324572c13b8387e8b453e1f5bbd0449f4e94d54878e20b61d132ad32028ddd93ce8eb6d7afa3643f524a06749f786fa6bd3c64132d582f8f0db48126f128aebc729998e306f005a797bd6bbb3ddf828c80c5697c975a652ac6a8703979427241da9f7fd13d2344c461c17b7d728637932c8df15604733eda33e9c47114aac6e25fa0d8d5d23eaa090e2bc82d84f6633c89a8bac2582c9d7a3f971f966e75a4d616bca3a8ab93d86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2b6c11223771191b602d243b6f5f1f5d207819daadfa9459c2eb08de399ca7f1d98d748e398be336421e07572c42774f013cc18819f78f13fc28002a0ff3d000bc4618c4fe206b86ab6c5aa2998bfef6c130e7936642eda75820475479d9428486d429920a2f7d778774ea90ffd126cb1fa12e94c7772162eb6970bc060ebb56ed1535dc183aee38bf510f7b96352f7f7a11cca6a04ce05d6f59cf29b07fa82ded6b2c2e0d42e05b571075eb1cd1cfeb2dae7d0d06120c8f600d3088b63b92ac5c8820ec4ff4d9d39a54d9a9d246bf2c5526d29d09f0530d93ea01f596e16db8718609383f1697b31414c74bf7eb473bb64226a9dd6dd477fd2b24814d6dbb8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8cd0e14bae3446a62f09c844f38a0282ff6756cf24dfaccea7c1d3b1d7292ea22526e7a43a8061fb930a711d01ecf40d518bd575a2206ddceddb4f562d4181a2fe20364419b30cf621e9f380ec36b2fea76677416f60d1ec8e04c37a57dcb53b93c8d762b2317d4fc082cb5f4cb7a8c0b62c0c74e6ee47a5540b7a7324caf85088a49680e8dea66309eb0eda4bde691ec359d0ceb659e44cd5a08dc1d9109bd50cea5bdf05c7e53d5632b81c19f84427ea0799c1193737c2316db911e4cc0a6ba043a7199d7299b202cf557f6da78143027700b123ef402cd12db753716f9712be37ec0257feae95dc76d56e3cef3140d5ee88b0d904036a8d57e79dc96aba44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8ea4dd03c83d5e2de4fe13635fe63337d40fe4e162ab0c4bc6e4ec6161a9fe7333459ffaa0d7a73d8b1ce67b9750cd1850b399774e27c9c2e434bab4c789666e82027190a61db2a4915461e1e7a3cce87343fe9f4b159bb16be757eef5ca84819c163674bc23fd86fca5e43094f727e1ecc5e9da93e32bd1b7733cac86949b9b430fd7b65e6a14df25b35a762adb2fda0d985c1fa882301ecec59cf7a483450286269afeae0bad6089e67cd83f8440e706373b43a13f71d2ebb81854467e987faa05eb2cf271bcd8bb9cc359a1ff9ecbec51ad28e12251b8d1680784edb434a06bd132f8863f0f48b9ff60b9329ab890cfe8f94355c5fdb97cc057e28ac463b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h97cd2da606e1063d93b25e95578074e8bf399331b1622f1906d55504e6ca23ff92e1c967af92101d69169fd8472a8176573970d12b225c8bd466b35db8d83c67a79d86b6aef7385112616e87cf197128f80ade5e795a280c25580b40ae4cf5832b31a341a1a6e133532f1146e63dfb3f1be94838789d31a4b894e48fa6869d85bbbfd6c2e033889bcc79984b31c950611c181e5e458a0755bb56551c3ec0075f44da371b1615a72a4a25d340f668b25533cfc470d1f1c345ebe3e71d32bf74b1e901bc94d00f6583a3f430d69458e26c48b34624ac8affd20a5eb8344cc75453bafb088647db777173a7d3fc3c4ee7133cc8785397e6f6bd951bcccfc39dce0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h880b7c88e416cde2c5dc03d892c913c3b2e53f3b56529deef1479bce85bd97723244489bdddff649e470deeda19705c958a65bf0b2d01caa9a7b9f2fbfbad03399d0cf4acd9f546461bd12853817ae60868c8df55e2cb65b60bbbed483b7e4a4d8b04361416baa763e658fb73727139b4353dbab3072f0544cebbd0ae072ef9107a41de5122010db56a4ed0eb7dcee22e39024617d537736da512406a96731b780ada37b70d4ad80e799d5f2843d49485205438b3711a5e33e19264ac0246f1d28631b9ebeb3749128ce209b687aada219ec830aa7c38dc2dcb245d1e1e3fd946d569f2f0413acd6963dd4f570790477ab7bdebffeed48b08c7ee2d39b32c77a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1761e05beb2e225e551c45ae819a144fc7cea2147cbdf4be0bc38f0547581bb117d5ff4ea46beda02c44ea9e5f0d3452a02a205a2d9b5a65d031d515688ac73a982994e038132a401154424eca0c00c53a22e813cb6df60b40489f5991ac4679133124ac64cef65f1207fa16c19ab440b91982859f2bda25f4971bfa06276d235ddd8f88dd63a680b91adf7941d08ec0bb6b56ed8eeebb2a1e4fc4dbb321bfa08ffa2704fa7bbf3becb8510ed820f3d316a6cfd65b1f348737d22725fd47c391d3d23a87899c3662fa64d6d37091197ee504012b6ec53b12b5b4e004ce0bb7c9504d31994312c311ecee2c9e20f0b4e457c85f87f096d84d2bc2667e92f40297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h40184d5f22c69de641bab38b58e681725ef8885340f4aa02c74a2044d7abc38f9639bf582f0794093fe76f629541b7ef1d28ed3f604020fbd9594fc5e88d78711b9cc535bac2e3c93203eaf8d426fe34c317e81500fbc11f9b12cc58f486e74f632860687f0e5c4207db449ac7c5366a642201d57e276ceef5843fa3b89baa2e3fb31e20d928e2f4eafff757036240c590ca5851ba3a599c7dc296393cc0690bcd0f268ba13a04274348343d7af4bf93a2e067ad3079ac064a5a003701bad172e75134a3d2581ffae1a4955bbc29c0dc737460af57994a804dc82ed69212fb3a855858cd886e93c6acdb4d689bdd155c6f443265f6d29b7fb401a8e573e83428;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbfe227472d61d5b630560fb42301a735a6704e295b3ea822702bfde019458cc69cfb812eb1c36c625174d0743c2367c1cd72886648f76244cffe77f1d569eed8a25a942421c843336fd131c5ed48355d5201f3a7b38049f7d488d820fa119a5e80fa17853b6afd986ab20f8706ca895bba20ac0cba8141ff543276742bfd8d3c3402f848df0a52a9dbf3bfd16388f231e6a5880f8fb2cba8171893d00d28d9113100680ae03482135beb29838454c8f1e161325d6ffd9c7cd394d9876ce35dcf9f679325a974eb0c77c9cfbcfa17462d5e74c68e0ba5d27c53713691dee20138c37122d1e54edf1b41baf1a099c90a850682a508918a92275c71f05aee73602e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he5a956c52b0df343ffb7d232fb4926483e5f9a8701551306f17451537aac6a41224c6f198146829f615b6593e59aebf9b255a1c95eafac67d026c09b9f38b7faea4541b32f3c52688accb7e0c4f8c77a8a2647aa55969795e5babded54d3fd49865a1d7c29311217d5de8c08f4ed1e398d84ae8699116f25f8aac4b229c883480af23cd205a08e5060bda8bcbc926b2079b7a6a42f627d4dca6cfa30604d5b6838beae48140259f35a62cada1fda75530786e663af3b07ab415074977ce5ea29e35427e91f7be18798f98a58f5ef1a2d365928b8b4f5d27f766fd26a591ae15eb04ef10c22e9644a960a502e7863cd4be9d1d28fc0c724a9dc4a40425418e61b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h101e67c1fb619ee6ee14e377f0af78660614c1613f9f7e68e2ac07e0e82c7cfb4cd6a31a1515ed172dc92ea44f60ecef919270d70227101e00fef15ff0e3908047a0ea1cacb789897b649c56cb9a812b59f93ecd822e3eef66be19adb9f14ffb6a1e6187d4f3362cee12f61df6a19d6dde5a0cdf33900d30d6b2f804705a0343e8973b1914508dc5fd4f82327ec4602a52f52b5c839aa9467f9d43fcada37c448ddd110b7adde112f9fc947474bcd4d9b128fcb8647d62d9da758b8d5fc1002e214e8db71ae61c1794e0a7ae866d03e76b50d632f5bed93765a22e46c9b9c3d35058a6ac8736ade4d6aa74049b6d2a92fe931e21a865beaab9d6aeaed36c6699;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3b9a897dc239e4697592f608fe403418c4aa866140ee6b271bd99b1aa1257a021fcf05f8e4447c398d903879b35110c6867efb91788c0cbb004ac5bfe5c583bff83c65b04dfb08a5c2b87b469e36e439c3cd296b51ae241b80ac3c9933e610ce3b671dfdce357be46487cbdd69284e33a840253aa4520f6d768bccbd7f7a8d717513dddb95f68b85339f6a979b4e24fc633afef544d00d19a9b33fb62dae75da664441f786da0351a639c2a2e0ac3759bbfb5336ecaf82d98fdc9678fe8306f029e1f5cbc2115668927bccdfdeb802e65c1cdfc2873514fd4871aaa1fa9951d522ca415682c5ade4bbf329966d266b0af0631402400aed9f3a682feaeac239fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h871351215d5ac183a965b86fff78f61c5e4b99ee21dca65995589cf6ce6c26a8d9996d794419260717443eed20446e5ccf8cf98fdb928ed58b064a4b3c2a1710dffd88a5fab2e3b5ee583fb67f6f8ee0cfd2c2f4bb765a24542175e46ff153cf0490ab51d8a94eca838971a1e269b125c147e7c1d493290ecac97e87d567d0f2a2f12da1bf936d8e1957d10ea099c6ee488d9d25e52331472771012e4226e0c1f83ba40d42eafef42f9f7ed41ca03d7a2f254c8f92204bb5c60c791afdbad613a43a499752ccda6384a3baaf271e9e7f6cb7be7989bf221b33ea6f4a6d4ba02b0e99d02c8296f1e4ab57911bbb27ee10e97bbb7f1194035e3e17c3d2e54da26b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5024e856822f8cf4693d21bcf870076c9e864d4efd4c48e937bb757013e9bc5e3eedc5da611a87a652f48fdb0a0f0a0a7e09ba31edeff2993d2df04e063ec2c758180efe52381e8e3899dd74d9f2fe6486e5485e0d7c8ef330aff539142335c84f394d002800f7c9f2159b9160a7fe86a47f794934ea610454647b2964efc1b6cfe11efb1229e14064f7197cbd778fe110091e4d18ab62936ccb181ea3179a85a89fea14b5f38afe14b928677cac5213763caeaf11aa9cfabb8163f33a06f9f50b117681d2896e56a40c8bb751fc8367b9b8de7ced06d95f1f4a7528f82ca175916f17c0f9e8833cab9da22e5cf6f78df9d3175763619857099a1c334e5cefae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haa67ccae35b244275ddf5e1944bf0547f264e027c97d12a97edff5306c3af694fbbd72338fcb4a63d61e32679db4eeef576e74b95bdfd5e8279381650e4c3a43b93ab6421f5f9c877f56766208d20f46e7d8c04598c51c05873883f58a21284019dcea93b7b424cf8ce120e8374ea23354eef6f18bcb68f7ddc2c23c36234d2306a092b9c6268f490a62db406eca79224815f2e25b58a79109ab166801966f16b72fe878e76560eddf131ddb554dde8a38239aaff0707bbdd66d7dfdbb9b461fafba3d448c71b9817a0bc88af05e344f954eec031ff0ffff5d8514bc1a4c60cf81435a39d1866b4b86ed12d304bf712c64589d413486e82fe24df880268fdafd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7cb953a1f72b20b9327778fba801723b7b9d2007ad3b5bd4e90b98889337714bf6631fcd9fe78fc44c4705f8ba59c99c2183fb3cd3ce67b5511c5bec293b77ffea37951dba277913c937bd2bc7e557f1c9df69b62af788450a6a368bc11e620a5c1f690cbf7e076acc1d22fcdc997c6d768b9fd91502d3c3ae7f2f9df13892acc68f88d905abfe64261724d260001138c6cd294b50bc8ddbd14718e17f26d0b84dcc44e4757c967f510c3c09311ab8f64e3c41c6f2662acee3bc36224190f4898bbe6ec1c3a23268a828f4beb31d7426ff0ea2a42231802e9021e4a9c9dda7fc7352c52b38bf5e1312eb73b5da1801fb219ee51674dec45b8693468bf693045b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h62f1e61df185ea85b38518f80d4407661c81e4d7aed94611a360cef9f489088fef800b16ef176b0f00ba1e3ddaba7b56f726f024e9fc8f4b439bdf2ab0c1d9f38ceb6848b0fdc217629092a03422c8f99da9971448f71e129d888c6f0c4ddf5bc0a799abd20eea355bad523fe8b64d238f1d5423c6632d69c7c0416e9bb50b9f51bad94449448cb1366aed497002863696dda31a7c511d35b9a2c35bf17f2846c704716031c638cf2e34adc331022270c614e021f377c49afdee2f0a0562c3d8ef6dfcab8c38192fe38bc4702a34cc0421ea5c1640bc78ff5e735905d6c583b653960b597d0619896eeb73ad8b49604991557ccf2e24f4e7ed9c7f8e4482f584;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h77030788cf040e5e32a3453175ce1cf7e0bce626d685bb4f2a84a9c8635e369cc7d25596788ec50b8e56cb02e0209b73752f3a27bb9402912bc75a01d9a396972fc500362c4926f0725ed7ab9be7a7254b21251284e09a1049a897284577fd8db8edb04b0c4d3abf2a6df5b6ea4bd4fea527e3b5c966a9fc602998b5613790bf9459d9f91077226c689e0d98be8a28f77dc152a215d233152aa09f1a89758578adc07690e2345a635819f6e677105acba1220ddbd17d01ab17eac9209788f6a4d3f5b6ac67e1e93ece9a30c18a3c6ce03357f75eec18c5a9823f551c33cd853fade8e582ca4e6b0cc0932019c0150b38499311ef82b20bdb3a229f0dc150d47b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6d22fa780254efc415a20b478cab973e918f8f55260d8037ba9eaa85563edae28346bf78888a66767507a38a577bc2abd6a6b929b530c27d5542a503fbf6993489bca5c3c80705b192562fb6c7a370a4430cea255be7b40efb93626fb9a3b36a22b2fc3e1ed9d93c5f58cd7bd67862426bbb544fdb85f367a41c666fcc2a80317adc58518af99ab0907d942fc6208fcfd84d8a90c15af8e2a2c68a2035e769360968aca17238245bf99f8899e830cfd2a64dadcad717837a6e6f396930d980f824558b68539cdbdf29c403661a197730b71196e401b81a7809a4c98256ed9366127a59b99ac7b5ce7a2de4c3e40f5545c48a01df1433609f4736a6673c892a5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8c0924a0db35bd72e0275457e5a8fdfa59ccf449de1dcab84013e4475cfbd66b5089d3b31c84345b0e52fe4f378cb2f03b5635bff183e5538418d104cca10b7f841546e26889fda424beb57fb16e5bf987f4c5424599af8319dcf072f4042d412bf652fd4b441bec3d25549e59a461b753bfa55682dfa58eebd729fc4d17d4cb2fbca0f0cdcc9d5d5e36571d85c1425713d87b602b79ddf5846c998c4b6481bac4e9f41275b64f6382fc2bd152fa032ca4a9f9dc464c2eb49580cbb6a53effb10cada2160c3e682809f0fe7b7285704a03ab362968283d80e2ac4177fada4037d4bd4680aedb779f31934b1a4e05e73bc0f75107c5d316a7a2541de72ef673df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h52a2f6a8dccb7092014d639175d41e1c3ff0edac7a8e764571ef7ae1f49f5b22944cc6577ead61d8a4eb02a3593bba9fa541cbf0560e962feb508ba94da0ee58333d04ecb512ea1e92f506687c41b70e76fb27653dfb47c6f85edec59bb79506fc5f85af1cfd3ad1aa70624066b7072556c1d734b24e3ffa41782729537596d5e14f2bef385ffb809be165435e4855c451795388f859658ecb98f6c0593096799724374af9be1f3913ef33bd0ad96f61e7370a4fa95153fd0341c98836fd743b055e6980aa6ce87fb45414ce05ac2b103f80151037975d1fea035b7d4d6ede10b38fa3a39e2774167a8704bf9c8292e308393c53ee157e47e88f1e66f3da4d6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd578032c88120fcf93ce1167c97e4420ada25fbb1a3502e6862b2ab22a032f5ab49f7e2c3756b635e734b9b0f362d1630ea2aa530215f9c43020a60f3ebeb204fd1ec62bc3e0acbc500326150505b2b7d74f0b60f749ec46d9392a75b22b32542f2be6b10c9e2854e2525df710a872dcfd9096606e68d236db293f12741929dfa345ae529d969f1c6c900460c6e285e9258c5886d831935bce4a47accf2f13e402e37e865fe2f7a42a68f271bdf362932abb545d2c48e61c53f3cfd028a9098757f715269890b83aa12beb6686586700b98a3b3bba371ff28d538aa7de76a6ac89c44ac8848d650cf07a0f5c41e31d06b8105bcb3b6fc4087b0e589fe9a7491c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcca3ad7fa0258e92cbdd194fa5b2974e583153b9cf22668c7d23c2b18fe7960e5bf7b0f4251b6ca5eb055dbdec43b71274929eb2c37dde5e98a719b71418f83c9d1162650b407687ec66fbdda458014694c1e805a71379c1849ee691716200037041d14f5e95cc468a091b03666f1a310ba364e96e925772f5ab27c384ebf5636769715ca9b13bb20c502c61f2a3501ddbb0da330fdf34aed645a2bebbc1b631380760e0db4fdbdd7356f20b98207b2f584ff374b645dd71d9886689a291a05d009ebb9532bedf489ea0605bb5552cb6b6cf58ea3a446fd1be39ffc7dbd2b5d38b30e39378ae7822d8938e3adfb182ae2a5f86b5daf0e7050d9c1a30b74738d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h78d4fe9947d45eb08abce2add7acaa0387ea7b15cc07ff97e5edab5414b362e3fa80ab87ca0b2bf7a529eb646f68bfeed634ab3535046a1f25387d13b03df655afbdbd31660ebbc882319762977466a9a6cb4355f8829e043f2aaf32e9e89f4a581790c7f1e6343150ae435c9e775308b3a9a4ddcee3ab3487c2a6d5322f669492010dd189e953e9178df633837325d0d61b09807786fdf30c627a2cfa7ad3fd3645f7ce304291814477641a91c94e223b3c071a1fb9365a5fa5f65bd2be733bc5c0d8c408593b0ab3cc7083d646c81394f01020350c7fcffcef2e701e145609d3006d5f8f72091fccd89bab6a8fc95ae7f224755b19f4767049b1fb1f78c4ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf707aad4b28b5027594e5efa1f2980737ce312557d193b268b90cf045f32351cc110890d261be488d1d694992fd54f4244c1ad8597ceaadbe9621f3b3a225a0f0c5c5afecb0e04edd8ff9e1dbad715c3b3f1f6432707220d61a04881e02f2d49fce03e7b123ee03a45fc174f8a7f678cdc62cc91fa17c19366503e0a48db2e07a5f26d985f4f096ec02985065ee38b8244bee29ba60cba58d57da58deff197d0d3cd8c859e0b50be03b9b3229f62d86214f292d57bd9d4c8f1680a1845239a1137f2e558fd8925607bb0ce9756ade4462fc38371327175d8486db495e342007c9f8f909a5f0660e6b0b0e93bb60782ea7b10af34d263b0037b09ae083e613fcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb872c468b5a2ebcb5ec6f49d3c4678e08812ee73f4368239e92b06d6667bdaf63a47d610e1a80932766793e59dc18507af6405ea8413016f628a25ff47a4117141fb5befb69ee46dfe76fe8209ab609a00afc5bb0342d51e53e2811574b33624feeefaaff05d019baf0cef1f85401dd4d9a554ab2be242ff6e7a940500fde9fa0636fa7256622b450c82b65f82ff6d3938c754a77e4dc1af1bc82ba74fd045fcea35fcee0013725cbb93760a53ac314350dbb79ed7ded9432008e82b2a0b2244997ee11cbd346a6c6caea0652a8be0ddb64a565133cbc5a4cfa69ccbf46ee92c5d4ec122a635f075353ffd7df31b04d089d3c2db18ce943f8faf8bee216cc330;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb88f65755cfc6645928081f7b0b1ba893a0c8b80e340b70a274933695534cf32d5bb9702fb42d2e647330785e953acfcc323f5585950de04ce4228104112f8ddf70aa7ecb2a9d18c6427d6d52fd5f2f4186dc5b6ea65ce43e8fb2563278ee3e74929f9561d9ff794d22dc0f6edf2b1d75b368f09bc4aefbcd53c7ef7747329d1aca8ae3ddeb8d32a72182a04187cc9d7af2f3e74e2689d9bcc36f6eb8444ce979c36ebf13c26bdf9fe4825490b73f814f68f8d431ff1f55e2fb7ebbd6d25c68be59cdd193c1b74a3af493839fc5e8e690f291e200fca1c33a7b93a69874989bbcbd876bc66bbaaf577394753675cc679af40954a9490dc60967daf059b3768c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h57abbf19a759214e41b05d494b90413753b750044c3bd08b5dc83b62028001eaf9eb0bed35515135e3622d312dae81d09b17b3395d7331c94194a117f026f8479250caa320c4ef956bef4d05f283a00025e3321bf07f3b072388c827a9c66abb9bdb4784e59604dd370ff58f59c1598e8b1250be2f0d910b90e4cca1f74e32df5499faea3cb759c3636704cfe2c7a4665e3acd120077a245cc9afd3ce0790f82c3b8c3ac8c69164271250bb088579144a4541af9067b6f924280322e5a988176697897a370311ab8bf592315916923a1f2c3f312d3652deb090b9c6702e295fd046262489a4e239233bc8ef33543e3a52ca6e4455eb4b919339a1f601d22da27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h16f55cd2a2d08017b78a3f4c73522d2fcf107cafab0e27060d6774972b8eb36c740b635d4e9f831c567a11069b520a1c4977f8df81d986856c5754baaa8a0c595ade51128fe3629798527daf297d9d5875a026539fb0721cecac89d0a0b32026cd06a5531d05ca7cdb805456de732f18a6f599bc25be55a169369d80975331b71862648d98b6d0de58edf4ecf44affb1a4bd558bbb1604d82161b6b0137c9375ced8fefce398d82fdb90f0be0b3944cb544b55704c3c54e7d667087cb83aec2a382d496cb2e4c1bf699ac6575357bd73947fe7d3d8affbcdfc38cf372d1d5b8a3b82217748144eceaaad8aaf7ec428d0c1efd02751cf7b0a173c26b2d5fc4eba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2e00926fa2f8c95b9937b9f6f7d536d920df87816e95d9238d12dc7df669027303201f0f966565d770ba69ff2e014a12138f3d3498612933badfab490e0a6b9a962030fc41648031dea92e528c857ee54e7ee5a51be6145cf106221562015b26b8f846f9ca1e0d03a766b9126c6f237eb960099e65bb26e535781e201bf2735e5180f9e7f9812fdd034b64b70e01a2a55848096d712b829dd6a61ad7e8b3f8ac3dce7385ae3975f77e28b2ee3229f8eb592b889402c19003619d66c39ad8c4458a46fdb828b722e54c80f449cbba97d31d01b16f04f7b879037bedcdf4ada946c76ba19a0c20617753fb8ce42d5c066d76575845d439b542a206a04366ffaca5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h99a76d9959adac5cce28bda19b3b2a7f31c01c2737638df8546f7724f2fa7ca8ab2df96b69251df2ae0d09b094e45a2f35e27e4f7adda269c9de5c594b69515a1f0119c1486e97457925081e4af49fae89b5e44ddfbb483334583ceb520ed9bcf9fd397225f50795acb481429600e0c0773f2eae71192799d4d3e80c2cb40e5e23dd8c63b175321cb086b4a2ac2addfe755494fd699715d9386bda86d409d5ceb92d338042dd7caaeeb79ec0e2466839100afcaf3609b2600f061da7c37a5ee224c5a2a86eb2217928f85ac5a1fdbec8335eae70f1655b701d5e121ad55cf06a70c4da49030f86fcb70996ec56ae37d62123d473a5f5b9cef5d395f61b835b02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h66cd3a0e7d7fcde884df1e2c79190f52ed0a3d909c87a1db04ee1b7c7b030d917da187b636e1cda05e93d57fbd08faf81b709c7ef29c7c625c739fcd749fa074a9fb3d5405b61098d8a336ad6184c578de35fce53e8d65f9e61a7a11f7415156b39488212ab61a9f9b37a9ea11649a218cdfc6c2f286e2c6279718abeb36a542ee1887c91c2443b2533e66e76c4b053928d6e25d0eadecb32ad9348a6e81ad298907a886d6aaf1a17eb6b4a42d5021476f6fa80c8d0cf1fc7ee623f1fc2d74048940ca33dd650e3c10b57a7b225826caf391b52ac521d5b44f8bf3fb4deb5103224dadd6093d07e50b241053e71d5fb744d91a68bd804d96f193ed5d6e8cd911;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'heff909aeae7ccb10252ab8e8e38dd5f2b7ea73eed80894568a7096f69daf71a13b8bf6a7af1aad7ab00492d230fc278440cc7e3f2f4ebe457b3a5ab05c8eb906e3fb75355572146b76c2fdaa5b42e2a76aa5fc007e5b92854629ff386619a6e1636763abf17dad174967457203769ce5e940045c05002d422756d828a12c375070e922e9d093b7f73aa51bdf75f1ab733f619abcc5ccc25317d7aff5e4a5ca83883c9cb664e9fd14d205ddddd89ff5000f4dc2f600867842c9699cf7d64f4dc62d98d148ff8fde8e4e0ff9f5d10e7b3b4d1ca4494cd0fe68d91661135a3cea647b2333b26e9fb56e76ea95f8a8924a599b89bf5c94d4901db6e0f2b997b1d192;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf2f22170a4e905da88c91f4814472d67c478dd83d00ab16687f54eca4c2af913c37360f9db3fe7fe0ef8317cf056f23ffa98dc68e43306b7c1ee65a507381b66b4d78383fe8ddaf12eabf8227fecffcd7f7e3fb202b78d2be9a76fb8321922b1b35415e0b2239613ebe3fc694470683c38b3f11472214569d7f903309dc7736090645c741dcecee12d0de3a35865da34d0e1f06b187e86b7d320f2df7ed9ab444c60c705ec32cb8af6c1defeb23733bb555ed50cd39dc44d7037b49cb4eaba2e7c5a72c763f7a1d976b26a89e702fcf5705f3078755b24cd9789c74025f2f34e4b352f5440357d810ed4f0d22b6cb0fefc6d25de7c64553e1b11471a185706f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5edc1b59bb758e5b33b32fbf832df6e00dd5e1bcecc69f1a4bbdd51794045816c7a448e2284d862f49cdf4156996ee412e2688f47d690f239ddf59bc52d3f392b03f77342538510596b64899c4e995ae536372d406aa8f0643c377c1afcac9acac3fbfc2f45aff7d2d3c09ac0f7470f6bcc6ede3fdd5be3e4fb8859d820a79a6b3ed419e8a15d23ec8463c38cec572ed4ecae8cca87af9143426819bee324fd664cc03e0aec8781eb76e18450461238e0e9bc47ea78ad4dc61413b8d173ae25331c758c7286746f63ee605ded7501c2ef0f0d66b578a90602489796bd8dbff11346ba37fe3be81124825ca388e9de00822eca3f74a5a3b30533993e7034a1913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3c5dad3cdd8fd3f7d72d308ed8333157e1bfbdae8df9f020cc2f1fc6826cf3b0d513ec6d85e248ca8a0a86905808e9f7bd0c096f08aeecc70bb0aceb85881d2bc7f91eae64ec5a0a3427ad1b2eb519c13b88a5eb44d76d8022feba2b77fac5097dc7909c07956e69b0e2fada40dab1cdbab6898a7bb52eb644a70ed8ea12552f0b7ba8b2c77cc8ed1c3cfb63b7a0142e02c1603d92beb0c2b2b169c516e0a8d6853193b93a67f58a65777c1a08f4e262fd06655e4e67839e50da6e54b0b213a91b1ea5dbec105efbc1480d8f6010c997d721876470d7edb7427430d00efa79bb99dce81c78d0167ea6206a6fe8f0313659a6321a1b2018ae80e68c141c0ee8f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h51d929ef6d242e8e67c04e2a93724a16af08643a9237866824bb7a79548db0fa376280b85467fb7443542ebfddd41ace4c20fd45fc7f99f7b2e9ea67db21bfcb90a3eb118502871697cfc7246a60e18a56878cb010ad2f28ec8d21f5e50b9df476f21eb0d6f352f84300ca2f1331a8a87b89902eebdee1dae774b5e8422df90d7c2a42da3037f6b78b8947b227bdcca08f660589b2334c52a7ba7a69c8da64b5962205f2332349e7d19df1670e73b341684a466dac88115909e3476b41d70598d03d935f38797c5096702e0a73a3321197ded7ff13fa9def8f6ac4b4fa49e262a290bb316849878fdbdd24f5b0fbb9bef2333ea61308ebb9be8010487fb602d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1c32786063f9a5d07bbb64d772320b94e66b2df07587d4169036e8b6c2699905e98656826950bd645b5fc24e3905b2a1f2695b77e3e906081e3d67eaf4e521128a48ffa57ccbc931a6800b093a42cd6eb7b6cbe08b8c0b567fef9ee94227ad515f190324a475c6e8fba59e892f9c09ddfff289efd50788fb48f9b8b14b1dcdd28b3561c97891da799daef8ff48fe390ae57da70a82b7fd893207bd88f68445ad67e347528b39c66fe0997908ca8347b6487b55d98ba3b2d13856fb2a8d6f8de57bc2ff80af8294978b177ad2270c68ba00efac9d48ce838ddf94c44f0afe65a795d7aed697f228a515ee063aa8c2f60c799b7c84c4754b2e4fa93056fcc807e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h306c5824f6658dec146ba1b46a63c2de353a7e3fe9702e956e16d30e2e464fdf5a4a59e487764cca2e729f8277ecdec5773a78d858e000b4eff2a7eb8151fb681a037ef48bab73062cd6a18576fad3481f0d74ddfc9da3d88c46b6ab523b76ba68d908343abe7a8cf0dc1a67e2a88562c0bb8de2de028982dc3ab7beb4f568d9ef5fcc07929a11716127b2715f4bdff522b4b4e1d36c2ffabee1a5fba35a321dfe16d3e5b75bcb4023161f25050d53740664933733068b2927eaa0ed70fa492db5c46638efabcf63b493c866274248fb94b47aac7bfb76a2d2ca0a1b485dbe8542a70b966e6e7481b05d28d64bf84fb59257104748a162345e3cdd1319a15f62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h87f800339a5ccc67e5aeff566cb370cf903fc5150afa6b512651fa38272997904af95df3a939f8616b97dc104143daf13344a2acbeea02b779de7eeaaee5720fc2118cd9189be14bba0e4daf19c3b3fe76d3714a2bd1335dfdc9c87e38b7c12f23e4fdc7fbfd6f06dc530bdb419766f650420dcb7057a41b154daf5482e36b65ee3b3e8644f323b79797416e86f0f73471d6232e680c7c1aedeef60be021def1e6ed9a36ad70f95385c1ea496f7f0a27d7e6be6bc86290d8766b13a059cff9d8aea105e889cc13e2135118594ae554fd9120d39e4b7db98f5b87497230fd703c8fbea6a0987f8ff49994cf6930ae06fb53876d85290548fd7e58dea441684a86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb80e58667d9e9d081b2a5326203d8ac8b5df35fb94dd2bdb2686cb8439c9f7719ce6c4ba5746545f364c3cf0d8befda39db454377f09de6a0a275c0a45ebbf3451c4b4fd406653692982ca2bda4c631b5b9e14fa27f2f7ddc9a0b1410acf051f85ca46a0740ed88e6ade7c9c137ab32bc6b4f4bccd337370b355f0d5b5cc401471c0edd7ad771e8451b4f208e3231eb43133d04a3d6b24ca9cf59d58d10f114fe5c12493b29befe0d057fc7ff28e296773dbbcf37b3ad7f0c980fbd8c082370ae72b4bb7032d0224104c63f62c16f28a8987b86abc48d0ae647661fdba48fa6900b50d90ce2e85d9e87c6531f8cf84e8a0c2de9772d450bb26e794e48b63a868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h32fc060ab9e813c60302a07109b298e4e6acc593ae1b087082aae51510eb0b00495a946af01565c120e3d78f380270c7d165f4659c36a9c4fa7d15bade644073df8238c6b9add6f168428c212ac75850a849a5f74f47fd84c81796260eb9bc57eae915eab1b68efb0cc76c735ffa91b897576f3fe57c23392dd3fb6d0607db41bfc920f31a72b8adee161478eb7b66fe52981cc1e3bb25d3d2e44d5e41328cb7d105c16c4fe170eb931c428db0a40dee48d3947771cc16592fa38435c0ed118d36e156f308e9af94379cbef43da202b19fb036b46fa1e9990bf6331a544990c1a8a61dba6f389ed9881391d9957888500acebe94e1a6e1d06e58e9d8921b1099;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd50b23f526f7bd75db5dbd2aa9d99f8d2e6fd92a5b13d047b543c9dd946361bb8a14309aadc5761af4c55c32605d9935d2b12d6a62dfbfb9e7564a308d453dc6cbdecac5c42cfa207ebe9e9f8c7ef5f8ad3ba46146a881cb0819b6e7be76926b0f47ce195f8e6fc6cb134897fe917caabd17dbe14cc479949fbd98968434391d57515feb8cd350963d0ae4e77f8d5d0a2933ecbf1dd6b0e6fd76a14170d6f58fe6f5e991c252091a2be7f6b27d6d1a0650399377a6b35358e1b985558a2877d31231ee2018f3c62bfeb1a97a6f66e643b72a4e823262339756eff56631fc14697faea94dc186c3aede99cc03094df2aa8a5f641df7f096585cf4c250f78bf3aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he3a37c565a5af73b1210af3618ac9092f1bbf0d5af9573481c978a05c0a4aa7440e6f1fa165ada59c15558cebc69bd5dfd649a6bc21afb6e285a44af22f0c5e0c523a6d23cea54faafeee4c487973338c53955096f7827677567b115d8cc9d8b800f88e2f8676dfb1fa977903a292c0a4998b3fd221e76c99742874c129859bf58c5d58715b1f2e05a8d31ac6310ac50e7afec8ed3e914c17f56fd128493b2c2094958c88b1e6c216cfdaa5f42631d38b4187aae093ea2bb8bdc5a92a083ded51386728f0c8102056fca16b30a3c336f6919b757671c263316e4626934d99083ffbd37e94a2f0a6385a171d113f0823ac1d0689784ac6f8de2bf8c69b59c8d4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he0cfb74c4950cd41db490d162c92ef286a7bebf2a7c1a6a789a8e15af65ef4f50c30011beae5fec32ebaac89e08474370a656710ca3dd44f857107fc4825ad8b7ae1f9fcfb3fb9dbeffb256633843f11f54ee1d08e90679d95ac23255af67c524457cf82781432075cf2f696b3f2195af9f408eb3f00674034d755175734473e023738d4ff06227c87e9cb3f523b4085d0378e3df7acf08f29a9d0235590e5f9886f76ae2b6ed611ecf5a92081cc7fb9201927e75df1e16d6d110ad4d1c882aa567aaa5d4ab88b45b4dc5eef74b024e7e7bfeef71fd7675f690adcb0835414bcc268f5be7830576b650cab88231cda6f272d27b2cf4588cbd1ef85e91435db73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf5cc109a79d1b32f428380a77469a7407b9e52318c5f00f30d6e5ff0993ebaf9a8e117ca286a76a1a165a1ba7af811754f3b72fdbbbaf57ef5bef3cf2f6e1b14b1cafbe92e5955840f961b3a887a87e2c40b36a84afc8ecce42537b754e31f7f7a807deecc785e8662d3adfe53ad5a5099d60f4c07b4d9c629fd25c89cb997f728c1454cad34dd7aea379ccafd431a6354934697341dbed0955214e2f554481a2b0ba19cefc828c6bfb8e66be4ee56cb12aa7e91a25a3f81a31bd451ad5c1d9a2acdc90396a3a347e73cad006805353a499467efaf34a0d4b20ce1fbb49d9bbd848a5975504757fd1c79ed82b9d4e1ee1ad41c24c41d37555958ffa1138dd96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h33175d92738402060543e314fe0bbac11915cda9c4afce776866291976c38e759e898aedb6a5567185f25bdc3bcbd3f3eef9256824fc9da6bdddcc943935a04ea1abb8ec573fc4f5895e7fe88b7f56b6122efe9b630c397bc68cf08ea0a85f5243a691007ea8dd17777306160841a2bd0802debdab921348c19945bd5961c6c96ae83dc43321b906a38e75eef6e797a2f124d5e30534aebcb8c2cd7808ef2104ab1d8f5e0844c05426cdc7d85d61540c31268b5c0851ceb15e74b845bcbe094a0ba1a0c65a7809d7e17b57c181f6ecf9873be575df85c9fd725a77b66ced4edf3e107211ae0bf180100a65726198550b18962b0275f08f750fdb478b515efda6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hda6ddf3a14286204a50aab31f7345719f96b4ed20c9ff1270b8a173704769a40873513b67334c2b04cf116b8c18c072b068b53bf9743fcca5eb88eb8e8c65a059cb3c65e5e43c54b70be328a4407e021084141dce312f056f89bd4442031a40f15b39d4bc7ba858bc52a791073a4405b5b62e3339424e5ecd91d8f5384e4b63faf422193d6b4f668ea39d656551eb444755538e2a1ccf90577713bfb89ed48a6e8b28326ad68d2cd670770fc29f433c065d13d594c4857c7851d318b0af9cf4c9fb3bd18e4ef55fc72bddac16fcad03bad2da37cdaf580255c572b87761fd46a0570b4c2190e3854b5ec718b3881c06f574abaf28327b2dd31808652a7398bc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haadeb91a78522863b4e580ad2855e955de6ff262b313919ad5744dce2808bb597ae9f92a1331c10e518f80cc5b0e55398c397efc37df86e513a3efeca4b87c0d756812db5963e40f5fea289da83a06ba5c7502cd6df272c634a64890f8f2abd58ef867ba36c4136cdf06b21b8d817d886f7070f496522e04db438a6ac5e826140ce6afac51322e1a4c7d09b7a078e41c68ed81a51da1de630b9993c3786b12114f0021f946098c1fb8f1c7501674a63c86797bb92ef17a9202238547744efc5475828afeee01ef897d39b44d3467c60c3fc92893a7ca0e2ae369fdf4c726e485c6e0448a55941a186067860b11f8e5d2e6b927166dcbc7b3ec66a58cb5d547d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hba690a2042b4672db5f439a7589d8aa72fb25cc625d2f8395d530a12b3fb0be68367976977eaf4c5c71d769049a1d3b00ec11bf496db7d1a7ef9b88566943439c67107335f016214d142f724201f11b26862f6a5e5b7f3dd4e3ffd4245c05d5d99c816ad2c68d94b8bec5ebd8d16ad29bca4eb819a1a08e52d728d82fd83f5a55d2cd5ff03f996c2eae2e39a893ea7b6f8c5b0c0213cc7148e3b9607df5d3ee218ce324ccae4e811987da890c6e2f589c26708e19bcf44219facb6f682601059597bae90b4ff5be1d560ace2b3c43947ce02a186709411111d666b813d1488577de6ab42a61ea0a84b9631c6c6253430230132032684ba23efc861f16dc99391;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h328e147dc4d5a8cecb5152cf96d39e95831869f2ab921cde7fe21963ef518a8c46208efba45548007598e0c555a18aae3bad2757534e6f7f52be629004d824dc86f6abf2d50a5760dfaa9d4a0bcb1b0da0f43e00e9c1b1a6e385b38e36103bd5f0222b5a4acf4e2cb49bcea9db591889b2619604f44386f782c887679302cb084e04490bcc4fb2c79610f27cb457111056ff6953a3529bede6806dd68e00f171293e7b06411905ad58b1d8649bd7f66b23485c89001203ae5df95a85567cd6eaee8523f284e50d7b4e31c2c43efa1e29188f2cb142f6841e01112b76818173d149ad585f0e4f92803ae0aed0bec6cb2e6c99e3a47643a6fe3db0f3d5e704bbf8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3146bea1f127af906353c4c06e3e417dd676b6e34dba2dd6f693075d7e8902b1b413ce7456c870a31c4a2cf38713f4c9ede3f6897b83748c110eb5566c157e0c3a6d0eb5377849eaf86205074ac62b95a45c85ee37b469a12e0d2bfc1fa7bb072ed9172ae07b831af7e9bba36d542a0748c18ca23ef2eb9ab837523b9df46b984876a5e42506aa3b65412d362ed806debf818aa1b8e8d7dd64506070f4c893749150bf89c7e1d61ce11ab8b2e346e4885b4bb288ee5e95a4a796a374a5e8e9b972c42c6a17f6051e1698f3df903a05bd9700904c1eebf2aef426b8f6b23376b2483628ba68c11dccd46fd6de1f6c2917d2a048bd96e0bacc032a91fc367bb407;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3d7861da132bb940539f47ebdc33fc7e7c3376580df447fc5a5ca56ae99670bc049c3107cd6fec44931c21ec77420dbe89aa93678b8da41712d75671c0d9c0f277e57ae504bd0249badcb8efdca16c734785e1dccdb16445424e4cf26ce3552fe117fc65aea762c3cd1b4f265004a1a1194d3f3c9e364d71f373bb523ed43048f1432fcc58798ebfc262d928a2297cc28e67496c0f69065b978a526a615417b82900f04fa7125f1d6152e1a5dae2228fc62ac68619f1364c2b5e64bd1aa45ca938f631df38757581e531a65092b808784cb9cad9681e512586446bd62caf117c9b0a7ae43c81009e2b589c6ebc0eacb223bf6be1af0743f7d451402fa35baace;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h44db97fc0ba2e807a79ac1c71693e0d8f2ca4db943e34446190950c0eb7bf81b64a1dc3aace22210fdefdc39738d5e1160060b2bb8a5fa606326792d265b0afad98575f0dcae5bc5fb59600768c8342292434a8c37162054188588bd4b561c9321a95bbbeaf9a08aa832834b3059989e8dde6212a85ecc643131b2892fedc4883ed9a875ff97f0c557c1532520a3f398278a8d262168d2c61f609ac57c05627d7e2b0839984f059a5edf6f455d58382e16b7966f7191aa215867a7916a85b994f307b1db9e5dd51fa047ac86859091a3a89dfdc84782e5cbf6b58b162463d700c09840f0bfd679fc003d1f78608e127b12dc6d93742f86baea4266c3ac7926c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h895b63a6f22a109e1f378733737c142a4586f4d6b45fb8279b7362490bce1fba570c35b51e6fb29e510f15f3d9df1011cdaaa7681649713eb57fc47ca8ef30f37555a78128b89001b2d02ca89d55288f5d091dcafbb66a6332709b15075488d7033cc9b42c9db7832843cb4092c925a224dfa0f4066b180bf7650abd472ef9091f12936d8e26972207db3fac1f430f0b89c2704ad2c5b03595329d34ccc9ac4f98d41a3bcd2493163cb2e5fc15ffbfae6003827fec714ce77ddf3f474fa385da2daac293d2333741c3afa984572577919d45bd2a8a099d7bbb24bc19595fa070002dd908d5035f5a9484cd30654874985d28ee6b23f2419930e7a5c679a9c1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5c563332d16dd9c298e252257dc5990cc09278bc9247ecdf89624b3d283ab9fff98a3e50a30942e19e4666894cd281a21e0a482a1ef6afcfbfe7f05a0088cdfaafaf18595e8189a4e967d816e66bb9057c7e5b95d337dd29fd4aa9d4a76db7bbb55bd62535a0bac324de5bdcaddfdc158903d166a8b129e1196af212b1853eec8aea421e40f2e6319df878bfd0c5ce6993342a9c2c7cb462aac348a72b7fcbc8afba39334978ca30ddea1960246eb2cfe5703b81e8d33864002e081bddef74cd96a6006adb584b6464b0720b1d19fb30559a06b74609b190167d23945c422531753485a077f985ab5402cea3f6b44ba7f2dd07dc663ac0518c133d81b7010e51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haa6dfa4d095fe5dbbd08c91608c2eb48a4d3fc4a258e1c94a2ca68bf0cafaccf8501a0375412b1009534969fe20d546530a632d355fe936b43eefe00f04c60dd895684affb1f652344700f289eab6a7f52ba33b538ed1e8edf81109420d6604d17275f6e7a42a846339dc0815c337a919e454e0505fe9fee79d011b872560eb145237ac8a666d22d819c84b2ed5c2f62dbe743e0402cdc00f22c2baa39175dc13135480aec337c606fec36e9f0e49662b62085822632287e6648e217e6ea16af89f6ce9c2e4beaaeecf3cccf260f0f36500460b7e4df4addac63a44461c1054c7541ea7f1aaca4a94cff1ca8b12e730eae219758a3653e96f16936744c253680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h74d22de7048f0728a0b84a95d691702a5d20ddc948f5a65983771eba4bcaf3906605fcea927e75a41d432ccccbbbac5173c95cc4abee5bec855c720410edbc53ca1f841c6fe04bdbf31b8156e65e83f46f5eb2ace1930109e322c12566adf158548ab990b2a752ef064d8ef70f053ca57c6c649ebe61da72e2294bf73f39244f44d9f29fde81ec1ae0f2648d462ef9cd8cb6b1f9ce85618059e4e8b42231a5b40d0579b14e6aa0452da4ee13781d46ac9a9449cd8921990e252b7f027c59978e4774f473a5b476ba815bf05144c31d81b44c3e1760683a5e7664adac1ce7e886919b1484af5e36e558087d09bc2e31dc1f02021b2d5e1e4828108734a2a4f94;
        #1
        $finish();
    end
endmodule
