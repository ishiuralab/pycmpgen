module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [29:0] src31;
    reg [28:0] src32;
    reg [27:0] src33;
    reg [26:0] src34;
    reg [25:0] src35;
    reg [24:0] src36;
    reg [23:0] src37;
    reg [22:0] src38;
    reg [21:0] src39;
    reg [20:0] src40;
    reg [19:0] src41;
    reg [18:0] src42;
    reg [17:0] src43;
    reg [16:0] src44;
    reg [15:0] src45;
    reg [14:0] src46;
    reg [13:0] src47;
    reg [12:0] src48;
    reg [11:0] src49;
    reg [10:0] src50;
    reg [9:0] src51;
    reg [8:0] src52;
    reg [7:0] src53;
    reg [6:0] src54;
    reg [5:0] src55;
    reg [4:0] src56;
    reg [3:0] src57;
    reg [2:0] src58;
    reg [1:0] src59;
    reg [0:0] src60;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [61:0] srcsum;
    wire [61:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3])<<57) + ((src58[0] + src58[1] + src58[2])<<58) + ((src59[0] + src59[1])<<59) + ((src60[0])<<60);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28ccdd04e6fcd29bd83b99604d8fcba97afbeabd84098879694120ddcce4a67dd4ee47c150cb7fa59eb134947afad4760c4a414642b7a27e046a412fb2d65721307a359c519560d4ed8915d5baac473d29a178e9f334bbe6bb599945da2927e09d960213464c513cfb44094f4b04d24d424bf7468d54b2e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4c000e68fbe03d9a50f83106997011e54c94b4cd2bbce1139c6224a835e7819cac31e115194885bbe0bf9ae74f548b5f47fea947ebb7cb764fbc75c643b84a7858dc981cb358bcc2feb0bec307980438b0c2cd630b0fd4d88da31a96fc39cb6cced59fb3d8308176cf23b72cb0bf697e87ffa8ed4c65b21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1502d85c4bb0d376f9d1454d640314ea7b2970491aecaa4e5608645a45545264fb3b046ff080e64f3eb5557826fa387fedc2af59c716976d6d2e90824953d86ea41eeb845acf092cf38fd3f3cdaff83089f318bd3b1ee01692ec0ef19fe8aaace2144271de4b0936d2d2cda479a070fa40dbc5529a9cabce8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3325e4e94c00ac0ff115efd051a63633774f8243c1c5076680383d07cd0fd6503065fb0630797acdc303bc8c08475031cad8a2b5a28121212a9c8f7cd247c4137223d1e5148edd978d8b321efc06668c0cee92f036942d48f6c679961d565583c2596b1207a605c1d51ce7b620325fd9a53009f32308c04e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15034b581260cb8a2486d80cf676ef7db0a9834170c00e24d86bc6c95294858068ff62cc966d944ad46b9cea86eccfc68d9cd57cbcb0cc1b8192805bc8692674e6848cde7762d6da8f642536254f9d2a84bbbd61eb2b98643d9d5402bc9412bd6f61033e5e6e2b4291c68d62ac3e5aefed23c226dc265dde6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd22b59f7d0b5def82c8199a49bd3e235bdd8cb78fdc3a53f600dea42520f603ae679a087419ae47b1eb4a2b2f443269e48dfde8ab2652f25744adb8ffcb25216ca6f7bf9f3f08318a30c4f5d53e958ad4d898dc8beb7ba8eddeb3b33d3db6f9de838572bebe1f6070aa5af463d8b01557e01a6092ceda512;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f01468c7038918f615bfda2ff643d0857c7f1df4fefa5f48c81766256439f6e14194de94372e95bd0de25f1fc7d95b93bfec47cfeb7235ff783652639980aeacdbe228e7116d9c3f5d6a1075f791ab8346559669e35be04e0235b2a8334e501ba37eda0384c3e6be9bcef70cca45435fa9716360b86ec71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e6c384909c1ba931d0401656a37a7f2e4affc3c37482d2f2441611a7327f29ee2a834712d196e4a320ed57646a67b50f2904595555aa89e86421ec9f42eafc98a8daf4100e4f7cd2b8fd67b28dbb33d89502d2ab9ed9cbeba90b05887e06212912cf58436c7d1ba33f3eb54416b8db9305a7bed80b73eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca3a34cc93f779fd8b309cb8a00533535ba1ad76ae626da22ac2cc2bbe729635cd4308c79fb7bba2ba4b197eca39d68f0430a8708e8473c94596e827b4d2b590dc52f5b18fcb0d514cb1d27cf36f59eb19bb4a799b57b018a34ad6637230be827b5e1c37534b725ccb164462d3a727ae10a0038c60231b7a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba38527db8ed0a3970ae4e6d06f6ac3f7ac14c6072796649b268c8bf6431f6e4eabe0ff579cd454b3618fb61d1963d987f81207965b33ef81cb14880a864c63ea4d42b8e2b222e97b6a146ec948a86dd7e1a7d8527e63c60cb096b913834a38d36d3465e57b27e5e20928f391a7c1194579795ddeb24ba4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51d7f9db8ca96e5bf1b89d8edae3d75a9c177c797622cd469957f1b5f3161268f03fce3fb352e044f989cd78296a6f869d4f9c2c3a575bc6cbc2f5a828d589e359733c56ad38fdeecf8e61e20827839fd5ab67970c38920fcd53cf38654da5c2b5f853969cd5e3117e3797cf634f04a1175e8b4a21ad2fa6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99dd285a85192676996de004849fb06e499d00021cf558f8703c6b6ebb0acbb370bb400ae5153a1f5a02554ff609ba94b06941e4c08079012789455f1d250501823ad0d1f27772f4e5cc05c142876e2aadbe5d95253440345e3fb6511eefc7807b1191994e012ef44fdd701746e04175feab56f014984eee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7de55580cfa72140a22216dff24e646d7493ce628025d9ed84d7dae9fbde511ff8f39c28ea9ea0eb43b5a08dbc0647dcb4ee800778d95464b4fcfe74261e33077ebaf1e7f9ae9f80a596d3ad6775fbfab2ee27bce9ddfb70165f090c36b94883a550eb31e20de6157241cb09e09b40f681b971a426a42168;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d874a7d9622884956b7590ae614bd0d3af4dba2a0beadb4c11b21cf15b0e97da671c2606fce7ed0a401076bf61100d72933e3b9118683416bf7763534a4bb4cb12c3e5f3c297a9383e3289b619f37aeeea38f30c4d5f532ebe445f546269d0cb8870a2b51970445790b1d47cc7de1f5f980235e109ba0e29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4aefad9daf9d35d582f25f6c1e8f354fe98bb96a7a781822f01fa99e8a39836e73baf4011e63d1cd8df5bc7c644f69cf0367d8cf50f81705f10e03d885d0fb1923cade9b2afc4624a5c81e877fca764ee6042a1955bcb4c58a28e8ebe50ad3294b067c6d92060174dd001c6d1c5102de307b4746636079f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1479c9233ad1945d1edee24c8ee228a333cdf3c949067fe2dbc5d011804e2c5dbe5a016007ed73289293ed9a30f7ce5459538a4b9e04a7acc5207e30149d3c4f85bec27a56f378a176ef04ba7394b2682deb0374448155e87b91820fe1be79e131241db85aa03094222e16e23dffd82e9297abe26a440b96c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a30f1c0caf69bbd4b9d797244a1fe4f207afa4356e5953446d87f43a9ecf12905c61d9ce504db64482c3867e2942ea1b28096560ac4108d821d8c2b35e59f45255e4f0d257264e350963727d82b01082164ed82565cdcbad1c5e48ee61274878d3fdee9710e6b9fd0ce88dc20c23287f02b7e79cde469273;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9ba7f81b16b48bcaf8c08c3a101551818c04706158043959bf90dc3845df6506335744281c3d2ae5c4c5209b01f40b7e0b78026eb5286592959aecf2966c30922de47709f7b9bf4a8e75ec2cb11654db9de625990ca75cd6cbee7a0d1eba85b1d8d3cf17608462a6d266e91adbe5f88d196359b761aa43b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dbc736e63835ee3cfe8640184c99141ad9dd59a5afe44c1a4d8fa7cfc38e786ed6ce80928588db01343bd2e1df75b99a33dd25befc62e6c828d34cc8600adafa4b62187b4ecc214833628caac65fac9b8b05252b828740f45107b73d8b0f665c6568f1be750fb1689ea0305181dcb097c0c12b42a299e69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf10c76a8cf2d32e20021d2378585afc9e9d84e12b60d5ea759000a90ed7b8a81e4aea0dae1db77546deeea6a0f0514422e2565f365e3e8d8a478c2205e3f598548699314f47aae79e0ef070d0f1de3dd8f702eff75f5353b2c90a148e0f462f9fd3862baa55426c048ab9c8d95fbaa390d478f1f8d7a5283;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abe5f5751efb596bfd4244739868d60061b4fb7942951e225fc4d94811a37744ab5b7dc421ebfc5d41ea20a662bbad445c7da9bc99c003c1984e6697f267abf30a5d4fdd02e7366490c79f26287be97a0fd1ae82c4b1dfaee8b54d0974551c7bfd7dd15b7a6625327f7a6a8cd0e87072abfdd69f960ecd4a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3fd7139880e5f204642d659395c76cdf5ca78438dc28e99081c0630ca730bd3a690d5767bc9201960bde61a09be1e67f890fb47cdb6bb883f2e2705843aad2131608e9fd771da2303776c29048c7ca845536ac89de4516ca9a98f4b0faf1ebf7efd00ad2b3c9cc02c9b0d9028c8f72439776d6f3cd33b3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133a42212bd8a081dd19ec48bf438e924bb44f17a90298c073925878cffeb1d7e09ab0b13aa5b445f85890a5c49a387a7f1d66007ec047364169597bcfd6629a1ae7136da93e3108753d9f8fa3ba5244940f8cae2259da923103bc2e210934a5c6f27122c2fee2845eb415b27f2e4548f7c32dddf21c0816e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8732a839d63d370c94640101e274756aef8bbfb2a12c0ba1ec78e9756347f2ee87a92dc5e5512cbf18ef6d2d83abcb6529c00c067ceed5ea49397619baae93d4ed29cc0e994d2c36b0ca04a195843c9a6f8a225cded2d170e99ce6eb3a3b93d725ac6c2406379aa956bb09864a831823eb2925c380175893;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h895dfed209ca03cc0cfbfd9e33014122b5c6546675d52df3d1c39feb188129bce8e2dbbfb6fdd3187d66fcb758b4e267870147b664a1d7fef8721de1b9e9c9f62c7640081b234eb37e9cb2e736fab0c3cc686fe4161e53f8b9e2c6c1d95193243319a0e3a582214f4bd27f1f3d7bfc15512d29f20ab0632;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127d28678fac5b0e740bb0a7478effb4b9d2e6adf59f290c6a7efba8cb63e8085c37a3175b490fefd8cd83d9a7afc65b5fe3ce7b075488c8b473d2a23e7a15436db13d6acc7cb5f521d0100497e78a3ff0d33846dd27b506cf718a6678db9cae0cc16bad8fa2c0e3ada8fd8fd294a2399161a818d99bcfd35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181237abaebc46d691925c039f8759900f7f749588a962f6e1564c818345d0d716f75254d5f2f2ea508ffd2cb70f374423f210aa90aa91b7854c2e135e91aa53f8e9cc0e8604e3c71d14163d72f422fc52947f1491995e4d1e273d7f554f0acb62222bc2c4ff191f2a6770004c55cc65a362ff27940b7d868;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16aba36051d7b730ffa5fc1b678445a175ec3bdcdf5d55ff1e158e3c397a63c38acf176cf415a953894c7b18c7488d040ff910613b1eeed0f5d1d3a7a998ffde7335dab59f33332df80fd26c65fa816cd745659704b3be7d906cf065b2172487064a9b14318062cc22a35c58d4ef0bd700c7d59ce6f2f82c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157e67bd9a577a1996c8abec3f53ba3a1456dd8873f72bea2cc6ce05414ba57f538ad463755a02d1aebe8e269ba7101e670648ea7427dd25c3a5d3943009a013c12dc1838a1b3988584c95f955b0359226d99c8c510fb87b042d99eb9e1591f15b31275781d80a7d50848e2d4b82ac895a7467e734afab74d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3114554a8d6255f3c6fd53bf5acc75638e4f791a834134ca431e2ebd85c929cc1f4aa5a087e36ed2da44335170abe6a9c45fd77fe71ca6c79c0ebe49dd8ad7833786838e75a583c2a828f51d9bc142d94a6cf37b04fdb89a5961bfcb0704c37136127985e412cdeb1bb938573a46c5054aa10f5fc0af36e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10afd41078643ac675baf0ca3543ecfcf8b46b2c302b51911d5a5fbeac49868f1802297dbec6b6ce2f1c51c2bd4a2b4830125404bdddc170989b8fe8a916ab174864466a1fcb1cb2024ded6b6a08d33b56a2bc2d0a2f8d91698248e34e25e6d1321e5f76af4aa2cbba21e11cd0e92467c1faff5f681a6c7c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h345be4eb175c2218b123ae9eb011d039f2752f4f0c456935c0126eededb692103851b4bee054e5a1a671a26081c391f4a119224c0d000728019f3f5d68464a3faf50b15315bd63b772e63e4200e244dab2b9640de95a6de72cbb41602582426d485437e84a59b276c4cb73835ba9dd4b159a36a2e289df61;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f884d3e9c8b925b3f6bf1303ac478d86f67284a87bb1bd6bab5897576c28e10e28e8a8ab9ec3b8afdef3a903e005b36d876b2183d8f8f9494fd2cc8126b3ed81040df506f979a957367f09bf01806f87224ee543b2f458966201a17c91d6a775e33693a72261d496e0a3dddde902faa93ffcb6e4c3358bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149b79fe680b07d5cef9ca03bfbe261daf387efb2f502cabc480f626e46782f327a941269d6cd445ff4de90d2424372fbb8d964a3d025fc23538f0a5d697573bb297507a0c7d938d660e49d2e9cc4bdc21c6f9ae57f83d4d9d568778fe81f7351a2b6ef17c14a3bf32e11c13f8b4653d5fd50e40838cbbc37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66a5ba010118f914ae1505073f299cfc3c8e356183158e08378b1611c51b71a4d5582abfa939ae5e8f708157dabde7833a71a3ece7f4b41c993816c98c0b933e8773446e37189a06dcae22eb7b3ff47a299069d49b85b73918a16c229d8fdba7789d245cd184573d9c8d4dd691d2d5812871f09bae30169b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a00581e2c53e4714911e8823ab91803c2dd8bed20865e0079dd80ce0f10df3c4c1fb70498c067a6d51edd36355adb80e2b5998909ac8334e6132a65006c98f2f3ceb62dd654c01ac52b0ce7d098653e0d4cbada47403a1992f2b84d71e50edd4964fe4d195412b8e7673b12b7901382103b9a2680d3e9a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cccc659ac155d9bf1933aa1e88a572a39802f942fea58f0a0a6120b65712e226b99cc8e383e95b2f21fde93d3d836924634d2a19013bcb399c2bd7d7a64a8a627a75e08b162914e9ac9e36a1d39ad74682efb72d94b19895356d25b9ba0c0295804b863d438cf6831f2dca07d0a0705ca2b36e3153a168f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ea874e85bf81a75adf2e5cbaa219e33e2e5b7721092efa62f3a79538158a734bad7775d1eba1f72aa9a765d46e03fd64dfba8ca5fcb82da6c18e5cda045e2642e00d82801d486554ba5e58a331783717d2f63f63f8bd66e8275dfba868c0622ef8ba8ca1b95b9ecf174c54cb719ef9ddd7956e5b77ea5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1a6471fb0b9688ff6079e875792b9f06dbf11b3fa16b9d2001ab1ccc1409f63ca404c4ab2178d8fd0f06118367767118648fc6d697812b0de81e37371eb607fbd2c0deff79212aa01f8894066bfb142cc941f9c615eff7bbb08eeea5571547a1fcf9edf3dee96b3bfb879c2e087b07d849bb11c3baf0521;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5465d471c07cd58318652180decd2e41386a77e60a69c9a03fdd7521a70ca4d2cea50f53c032e7dfca0e4e7b3a6616e02c6e20c0d7913be98a006f2feded2fd19e3f59bf91d2ff778320a2f4a60aea4e2086fc36eaa36b4ce6b95ec6a2c6e87b17ef278218090bc83002a8652ca39b4ea069c062e5f9233;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1163f41935b9c1c77319527f83830697e773e511c2f21f18e58a2ceebd675299164bb7facc9ae94e4dbd3d036c317c60a04ffa385c31e03e7ae2dbe8777867126b0fa2cf384f62dc875349b983cd52be2528bca26c2532b8cad24afce732dec7e1e050491509e80219fd1303f441404844a196b37c834b11;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba62e07eb9648591adb16831af7d65c6f418827ebcc100f8c92ff3a96293980227c534b5d299bff430e5354577ca5e3d91be3d6d678547b2704cb10eb519a1d9802b746cad44ce2f46413c4e86d7c7fc034f99a2ceb087d3476936cc1962e30b02a9793d491f1ee9c5a9259c2b6c53d0242999292eff554e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9423ef46e9cdb383875c68b7c634e01fd0186c629e9bc216c07c011a45a7dd159b0b927ad46f2cab5b9e9ab07a89e0732e3005f9656f7f92445b4f58fa04de5646ef8809c7a267ab52d36082f848e1728046d323c6bd8ffee5aae35deafad051a8fe87d55f1053675db9cb3924767a5b85903c9732639218;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1c2e0cb5766501ef3029a2898a0446dc35931dc3bbe47b856a665bb11951aa95fc0d141f3e2e386e702b33acab3c689d6941e72093e4be3ab11685b98c9584f2b7b20676bc55bd973d49a1a6a22c72367970831d4eef33af131fdda8c4590f75f8894325553712b38c81fd403373430842ae0d8b13fd746;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba9895cca1c2e2922ee2c4a3de6daad47dcae0132679a2897a260fa4156da85d822153bddcac48f0517b6d09811945890c55703753cd540629459d882bb6049c9ef15fc600c845bda7a3fc6fa80026c9491119aca0bc0dffe945d20511474d34c73bf2bdeb08c1e174cbb4fe0ac265bf62ed33e1e1e3871b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fee4abcf8c93ba2e64183cf703754c59c688ee46099085038523485b9b5372f0445e0cfaffc4aa5b2b789600bd363befffa4dbfba691c057f623bf4c4d7c9a3fd0bd204de9b3112c3907f71c19fda5e71aef4f56ae9d7fb9ba943497eccd2500d82b45f0a20af8c70af474d529b50df8eff4b19428d06ccb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46be303765f23be545ec14f644c94b8788e35883c413e2de0e6615fafe2089094872554d87a4f101a78e2039354f0500bc85cbcc0b630aa02ce0f8e7e67133e491e3fee731d9ad5b2d77a97f41a88300d241a3cdcf51b64b9712dbf7fd21c1326e9180af8c2af391779d9d7e06a2e336ce9df03b3f248156;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf6d682ccbc29211d71a6fe4d5e42529a9933b65a969120c08e5c8d770ce87cc451384d8728421895d7ed806f976d0843ef86c1297df253eb616a330f361c277569381f702d5df0a195641c796de59618ed430479a2721650444e175924cc08811db1ff1ae4aa6f546bbe652fbd264e594a8baaa0106573a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8af094f03cf7f0a2d7e5efd47028f9a40e0beca11ce1cc54b0b96adcb0f4009b4c554584331b372ce3f362f81fc51dcda27a1f90761c69eb8758386feedb525fa385ae27c48e26e393dbf2b31fba1adb51c64bc51a701953e25529f972656be6b2db69e61c456d1a8a5c083b3d6904bb41c30a1f7b36fc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6dc6bcad8ad16d69322aa70b74d67f0f33ae84ba8c48257008c85f597b66d8fdfe57cae0e6f46ec2555fca6a02859c3c62aa125c64595c87da3b03bea21ca8abf7025195ba74d4ade871acf86ab4b953d601b3301c99be64e98b216c4a826788970be5799d78ce27f8da3879d4126a04b790934056c6045e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df4fe70938cfe61ba7db868a9244552b2d13d6ec8cf70a50e1f5d77310e9d6fcadbab72ddba79ff94cd9f20625af3253a94db1cb44179a6f6d1f4ee41101b609a0839f0917ea0734effd130b1c1ec9434792b31eda69e7e1ebaec9317670822740d365ddd6f864c091acde0ee78c89a6f50f5b35c3420cfe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fb0059e950dded6dbe0043fa1581416e5ef09a8720a587c459db70b2d82ad22da397707316ce5efefe865dec8d29157b2b89bfdc95f4f5078b63877a7762b442de70fd98b33507eb977f29d254c0e2ae42e3cf22ff9cac7ce9e9ec1f3f1480213ffd97498ad9db0652657570420ed3b125593fae81d10e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb789cdcd60904b60b1cd755630b05e5ec23a84a2d92f7d50bc0dc6c5dc8c014540c3e82abbe5af93387301b4f7a8720662cc00605f6802c688ee0f10c46b9c10558b71e1a12d39e4d1d57c52463b500e85db9ea1f4da916be8703b2590995c3c82d7ff8ebf1a01114e76f63ff723ebcf96f9dedcadce1885;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b6b2343e21c1e3caeaa373768b299ca067d87ae1deb79069297427946b2a53e5f8c3fb3fa3b8ae1e936e0771dba3fd69582476a689bfbd5926ae4cfbd06cbab22a9be8a5f81190366234fbc57f76980170b0a5f1ea0b040bde2ec8ec9d76f895721b17861f9381237c2f064fe4ad8283ed719ed8fe35e35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dec59778bd4345bbdf424f8086fced3fe471cc94ca2b0c580d2dfae8440b046f1ce77703530459547adc116e72ce42d07dd6c55d22be65dedd9a6defa44dccd852b2cd05f6c25037ee55e781adb0d55ef6cd12c1a9c32b919d3510708de1751a4f09bacbd317d6e7406bdfa46fc4109191fb2412e795bf8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a6d7cbbc735b8e8a0d80218f278ee9cb772b689b3bb9fec17e436e435b073e21ac535254fac84a04a34852c03124e4a56d44f7fd5f9800db6fc30d9563d393b3876e2bc2e5f52c304ad45351b8428f5ff85886ee8b7227b209c2a8e5db4bc9535477dd9533ae77a11d4120c6e849ff68c7cb4a71bd2ba1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5014cf7b8f8f72074c915c7587fc387fe90262fd75667e194b473c2cf022eff70ef3682a36fa22098392395bcf772c5d565a7c61bfc75d3eb254ebb1b47bf757848d975ce5a06129eeecbefc291277b3296f6ab9ec4d8675978be955e2e4eee9e0cc526dd23a7085e7e23a0767bfaf31da148ca12838dc74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heec624e95422b9b8adfa89602c0ba25ff769c72ce7ce39d20619b938b93afc232eef2f2df540c5c48a6c8a31369233b1b6803e76bc8ee2f35e8bfec363106e4d6094face28489fc571908a43bf4ca3ceb2f075631d9c9bdcec2a4ed25e19df064f8613a88f6ee7e355627b31a84ba27c669a35460076f016;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194fa81a886959008b661b38fe0801cb76dde4703ca705eddf0f9d6a7d8725be93029dfe34f3c99dcf82cdcc0c199c36d487bf8e8413369716e6fb7bbc4e6c5ba06447c3659259b8e8cf35108a6cf475342f11c4617fc3692b2c2a8889d1ecf5acd2ab266619c5712e2ec58a627024d3b5bf161eeda8a7615;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd7aeca27511d51e9dab451fcc78306a26c9cc374d1a4113c59498059c9017a105634193d6ab673b8cfbdccdf9c8c43591bb3aeadedafad3b5436d3f9864a99e3bffbbeda20e14604c2c10ceb656495ef5c9daa80c916bd27114705a49c60f432b5440e76c93415cd58fe57ae7b94b66bbbc146e955abf98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c59e1d61a1c364e6cb0b9a78038af74e9f53e24318ec24ffd988cd6165b47bb1791bc5f7921241da4b49e8f76f7f0da58f54796786d14565063baac7c2042c1058c80044c2950c50ce513f972d1cb1e15b7dc31ad6de7a3f5f17204818d5f86d6462ddfb50773cbba4d5d59540d76ff1a8eb1ab74bc65ddf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf73b14a3abec6aa1b6e4d1e3f18c5dba77e9a8451755f2d421d720eaeac63a33465dcae26f9a87f5508bcbf4f93143072f2756541469298aff7fda935810dd7343401fc81c262a8ac80b02504051e618524fc700e1ad2919176a6b5bbd7027548b6b67ddd41b9efc322f84928a4cc9e1a067b1223fd60ee5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12dd9f7a80ef8e91cc063262a1ce20459f191b469b8de31b895c675068dcdeaaed5f121ca734d730056090ef362f803d5b494f05d3ba5f196c2d657eb14467a80b108216a82583aa538b72b23f777706a020646468e9efa798855322958aec481d29315e8a8b8add96d8a13d9756562d7e4f45f0d5b43daa4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h303d4a77a2920cccf726492caa9606e0fc4d6588bc0b6a495f9757032740cdb8552d7b63762ff78c6ea868ea0fa5f184b5c34c2f41fd36a22c6b393b838c8a6f8a4d146f8608afd012c6f41d16f70d0c3fbd62a6d5992057cf818a8764b574f3f6b2a90288449d253bdce5714b546214977d3b5c84f84322;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a52e01feeafe6fed818456f0578c0de48a8ac75952c6228a24554037409d1c24ae16be3ed703b7bb2029561be9066b93fcde0994f7afc3f76d5a0d03dda3116e895c438ffbbbb5cf78edc99e98fb5cd7580c96da33e8c5551dbcd4c2d4622a8fc69fa617c07ba233aad7035042afbf596713d377fdfd3bb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15648c847fee017f6edc070b053c1bb90a2bd95ee35b18549091fc6781a97c78b2882d1abff9547e53ad893579f5d96d3a3fb9f9eb2a1cb7a20e8ccd43bb5d084af434bfc5d43981ab3229ea7f3a17a0c6939d49372e2ddbdf29f19d5c307d482913843d3d39dc6889243251d019c3cd30e6b84f1eada3876;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d72374ee5fa184372d1031b37deb10a10fd8260783e0893f34dac80e54e9647897e5c37d00ed0f80f73d5519953885ce6fa525361fdae39930d1878ea72f6447eb9260450f9ebc193433683c5a65690f99c6b5587a424b28c266d5ac22d0c177df304b570250d9892a4cab925ed875aed5de4393691b9c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5869b3d61be28211ed593828ef046d64fbf706300e26f370d782bbc38d2f43fc9169ee3ae3d6bd06b5e8fabc06a3ba36c566a9272e7168f74bcb56bc19d91e08b4527c7693ccf6916facaef7e573f966cfece39e065a1f6983ca4f37eb9dbdbb59c71d1a13514af66c90bd7dce2bc84d39578b70425a385;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef71076644f5f940fe5ab3ff370cc0b73fca52d39738ed888df92fb69cddd93005b0f1f137ad7ebb4535b1a69b33612b411c158be88a341fda21a3cec333b066bc48e890c7c1eefd5136a3f33765dc03342771802d74b97f0d34b9edf8e9508ddbfeac13a48938cce355d3c1d10bdb7a9922fe8614c99995;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13be62268b72edfe0336fc22646713aab2bac7382313ef7e26b03e3dcf4a3b0d62658c9f1861e3972a2521ca9fd394df638c8a6561f4ae458bc6cef161879c177525a61dc80651cfb3d832555529a1523e74a2249cf645c9ae8f78c9913909754c1e54f835c69ca14d56bc822edc4e411c1991cbe0fbf3980;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf92809961a853245b76333764dbba8b6cfc962ac2f75bbe3369d659d2e33abfa2fa9ad19a45a69d1321d3857a85a89cbebb1a75803c874e5316fb9cc4b7f3bb9de822716d1fa7c501d5c6741e21e3b2e312f02e7867a829e78687abed140f5e7eecc0fa14d503ac4b2a45cd75a0bdf98a933b5dc1d67334;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d679af18db82d1f349c059f200a897e728e474532c987cabe6bbf76f434d2ae3a232729ca00c1bde88f2cf4be661a22ce6c111aa3de3faa1ec9b70bd7d9e31be69f89a0aa7d61282ba83dae1d3d48fecabec7399d292b1709cdd324238633bc27c2d151bfad7d1959e8e5446a0cf21d8fed87a815fd7b167;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e810bd42ef3f510639411a5404c749b1cbdba4cd6176100c3bbad818f2bbf9a7a67c5766bb51379f16e093c0cda0783012552c8deb2bad1ed28f93ded8be03d2348a04f85f41f68a92960e1ce5271e7e1e68a13f10a07a91d3ea146cb8ea16642c206dbfdc13bef0b245b5eec718fec6226676cfb7a0f11c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170c818dd2ecbc386f7b18c6935070537d283cacbda202ac398f50471075b5f9a8454d6eafc092a6edd5702d11262ae1113a2764461af26c982f7b6c3e2810aea7a4037cd615a50ad38dceccab921dde6615bd056b3d0c0fc5ebae5035fd748b85851b2839221e1975345523cce9a16a425daebc943adcb17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12255ffc16e4d2d8d12ff52884dcb352fd9e4e558a1f4873ccf30f9a4949d32611cfe15a63b371346f079f1fae34e2d62ce82049bc1c9c8c72b4ea6545f617e0cf4224b712bb9792cc92046225c692fa424f17f71b0bd17ed53f7f37ef6dd87fa58ec2f7b5c7f2e76c5dbd7b3cb15e4efbef8aec46f363970;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4880c766ddab8add0268d38549f979435c8fa2d4db9b242f5e5970f1b5fef36ac29dcd1a62e15339c5608817bed716d8c6ca960139ccc2783003c888896e1646b42adbc94e82bab9b17ff12deb75f5c009e0a206fe7359ae16bd763a107cc4654ba31724be4484b983014ae219d7d937c517c6a2076cabba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b15c06a20caaa38486ad7dfe418522d567b83158f392487d2058978d81ae3aa457835caddbe9c4e910bb3c350884a007620c364cd4aa69e581c2c885624fdcf864deb4c9c5ab6f0413af9ebe98ca091417d9b9d5b6b9a9336bdfd6cf503cb079b4be983806d0f06f05ea2c24c1b021bafdcce0f3ef1438e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71f6f64f1ba4d30286dc1da65383bde9d8b53cc522f18443e0f320f98174f1035b94ce6485c4a345c4e5d3492717af7c8ec1b3c82d80d533488b6cfcf1edeb84d13bf49c363fd1bd9931d350673273b5d65c5a2bddb6f94fcc60e469d22c2bb5df942626e1828d2c5173063ccb00aec812379873ebcba40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1deb0d424bbcdf36318043fc23557be0e0d70e381b7f75b6cf9edf78bf83a9b76cc274fc7e4bfc077a59b378e041fd2d7160d285684fa7dd9363701b5e4f7fb387ea131ab16fcc8a165f74d5c9d30848c36f00322ac55eabe3f08012e413c63f8325ce8eceb31a002921ddecc471a180ec1f7ee93d7d7cfe1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38d1fbd042685cf65c2f4b56d6d18a0b3b34c07b22df299c0952e56bed0244d1f498fdc9bfbeb7e77771ea6d6aa05828b9848b3cf97668e04fa755ce31f537352c55a3cdd8d5ae3cd09b29a9c1953f968bd71d8e99461cef6873ca3e6db7862dcb69fa1823464c462c2ee1b847316715fa6d6508e78f6140;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cdc57c90f00e080e42b7d8592f7dd48a06555a20a6ffc88627cc0edcbc3f6064c7a6c12d4b1c210bc36f55e65d38ad52e7fa70ace7873a3b441f8418054b57c9b3c4fda87eb8993dbd0617fa32d7c36ae2d85982ec07b4b79bbc641e36d6b1dc074fbd71b3aa1339848c42925c485291e1b1401b7e30042c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1231d17d5e9d2ed73f5829f8ae6a4a4f77e211c655488217de7ec40b3140b37ef2606652dfa2b9a48125ee02eb06586ac46c0f8aa48ea804a6f2dd7eacac8c47e07780b04fbbd24676bb837f2d39eb2a5096ee52da477581c511c286f44ee67700aa2d13c915daa79c20db66663d78266b475cd228ce7fbeb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b303446ac6b20c8bd397e4936ce2d29162d012a833853cad378e393a14ec7b86ed69335e01e905f587c3d3484b118a7f419e6dd86c1bccce0eb88fc083ebad10a88e1e153342d1a5a8cb38951a5be1bce38b8b799a26f5c2e26069607c622b9db0c82cacfc66539c0fcc9ae1ffeae300a3822c92e36cb3f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab0bd1cb6e8f431810ce0b4150b3d4c27d84918ffd762847445f2913e04c967fda3bab65fa2824e78e0ba8f6e2932e65fa645d50d36a10700b3a8b7931b54beb6fc2543a3a573bf52e0a7bd7b4cccb8c3ff2e75486f8845df8a5f340b08da7f809477526722e9db70cbb5f0d5e562a14e20e4ccbee238d1e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc772b47f7ef817e13df744564ccb51fae5bf15e6f55ea80dc46e77d5dc41e7c2e9376be35b47a84e7c227b887237b9baddb75f6c6088887d0901ea582214afd7ce83993b6712bc7d9aeffb10ff0feaf8809901d7c9f8123a13daa617ddf5c482ab9aed9960b60e2d209ded21c2fd4384391a87f8e6f55d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8735510e910e71ef6ab936a46d21370dff3edaa337ee51a0b8cf1235a3f5d448555df06888d0a2bfd130cd874a041dcc1326e9bc625e5c07b796d1aa61d06d95fda36ce6c23b96a4f3f72bfa6620235285ccabf111714fc60786102b212a69085422a5a860e8c247936f3ff04846a9641684fa51dbcce0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a39713affeebc41f98f512913de5630383c09f3290b41daa0fb85d99b849076080d57cb7b5f387f4a1eddc37de105bc16aaad2fce0615d2f0cb30b783370e5ada1363d94eeab50e4f758158e7f561705cb100217d901798bca2e75b0799744b41c3ce2d5d936d26496d6eedf9e8cb201fb211d36f70ca03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c510d92c05cef6061b8d964ed6a96303d3d4b13d6aa96001f6b28ad9007a4f6a9646997ed50b47e4d0e11ef42cb55e1af89c03ff8a5f402e0a7a7f30286f71a46f126a8e3969d0a81dd7d795db266df63a91a5d7a3517563d901b14e46a1abd938a9edb46c479189c2678a5c975be37f5f04ac426229ffb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f186bdb589c045f6ee567abc3a6d519eee5e2b1ee7cb7d646111063e01d29239d77dfde8f7bf19f81d6a4ce6e6f9cbbebeff242a57599f904e735f577310feaa78b73ba709f2e6c8f22b09b256328bf166b32a3c28269e0f2f68eb0d434afd71e29da3fca9e8f697ced2203cd025f4eee463d93e69ce4d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3a98dc0e124f43d78af7d649a9404f4e69122f3f1b0c1a3aa04edc05c3a4302c55be210f36ccdfac695c9533fab7f037c3ea99551c7f5b1068d5e2fb8423f57cc860bf984e41e6e982a56a012bef25f06e9b41cfd6658d4a3f6e36edc4a7751a91ae9c293f39c72da97c7d85b3e2bbea9deaefbcf94f2a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba1552ba41bdac01fce1fd33659aa77818a4aa98bcd89c43f4faa1a96319657a551bf971fc496496dffcd7732b726063cfbe303747dc870fea5a7615fdfc570c1b8a597fa16aeb3ec3bcc54bdf56c38d3a93d4c53b950527a3430a353ea50283060f1ae70dc45842e177acd8b2a91d7871ad9694c3b472c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1dac99ca66044eaff6945c464e7f6d02a0274b80ff286111a48eb760b3d6df6fb7fc4eaf66da029b487871d8117cb391d22460cd874355f29938260cc2777f74bd24a43078a75bc513ae14c7c998a2e42de393f2e08adea8ffa8d1bcd2e146e64412ca8f82e4b309cc9952f37279c09c6e785c28b5c328b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1843da3f6080da0bbaab31c018aff4992bfaa8c00a673ed852c5888b0462ff699cfacc456832c06f86ab49d1a4107c915ff7a5a301fbd8bb289ad4f6d70731db75428a2c4bdefffe555e285f37e1cd9048738278f6c774f45ace114eb0da7055a63949569898dc14623f27af45863cfba4ab9c0e56d34fa97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b17dadd4c1579b4907daee1ceb7ab79fd1341d95c43fa61c6887871f90f287b8aedc2cbecf16932db89a22e4a3593b1f4fb74e7e72f237a8e9efe70e1d7369cbf35d514b8a082f7f8c978e149a804ba8e230144bbf48765fc7e189535eca3a772e83c54ec3da1f64b27f996637569d9c633a82913fbb9cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d83559357a602a899f380ee875f55993266a5abf7997b6eae1c44c0c83ffdaefb55df1d5b1bdd47044488973c51364ce8ecc7adcd4af58ba8f8ae24f2fb3379f3b807df4e98ba28a39e95aa834c008faef621f280ffc481c4c6257cfd7064927a5d597e815271054d69ce02ced5f3dd621aea7b77599237;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28c21a45f69e78f39ad4d220204e4b4e7a677aa4df6356b4bb3dbcf7a1227e879f4513f767bd27784f01fe9756b489e017b0bf8c3f787c382d0b044aa5d25673ca65e7f927b898a4a4681af27021719c7f7050941d0a41feb69eebde3aac71d539469d7685abae2aad8232a1d5001ef37f2a4c5064ade0e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128f1fe358547b34ec0cb485322a7bda53dfa8ffccee7c9eb9b72d1c9fc68b9e3482c59b505cfc857da6f07d6536380fc18a2ca3d54388455bf86c2ba2ef4fb446833b031e53d60c36f2875f8856515ace149f6c1b73c83023216457ac6eefba4d09899a96921fde6213d33a3e0cbf5dd1d07a5015cb77b3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b500546696890f2900d88823129991245e1994daf76e3c9f0a2a43075d835854f39d131f63e98e61d063e47440323e96599d762fdbff92845f08497676119a366fe65da0d4a37ba364ccb9e8d444d0da4e213910fa7d6ad9187e25228ced6fac4d34f7b0d9179d708a3f92216fef6b6fa882b59895a1ccdf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4cc245b6046d505e4c46cc23a4794aa27b3f6162fe2f687e6af2f75406af5d896e598d3c568ca15d1f64cbe14f6041435988b8bc89c7d3ee311d36d9c8e4eb1eda6d7870f87ccec0891e6298f5dae8baa3c09ea5e6caadff04d6ab67fc5d3d9756f5b3a7ccf36723f31400d783a64f0eea13e03d7c6f8dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a844c96ac19beda3e7f5124d42b2ae07bff5b776292ebe2fca5dd78f4200f529b96c571e12df00b355df64a443d5ed7ff17ab1b0ab435067855255050a0ad5983aee1c93c7438a9865e7a83d49bc281b78892843d14df14f01a86ea6eb21230e615450b54ea05c010c0e4c2033182da8beebb95080dab13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dcdbc254c0e1bf635dab8200da5b03e2957186cdb652503086aba7886a7dddc6f0e1269696035df56ccc335c2612d6857b2e5ce8b88d2b327d7b5db64d2d744f74fdb0ee06d6f962230ad63a8ab891218db095189c3df3f70689b1b7da0edad6e75706214802760dd1e930090c8321b7c2110ae9b1fd233;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39002f8d61827346adaf4b89c0868cbe3b236d4479bdaf7cd06e33b6b3b382e52120b5fbefcde7214bc49550a437b849b5ae5e9fb7d3f43326830ea1df8bfdc26cfa22052a8757527b5cf8345da82c92c8df6f60a059ede8cf235e12bfa58bcba94f0bf6a8112d7f3b57ab93d32dbee763c70fa3ca106828;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d18a0b4e5d89c9ce2f12b32087168b6fc46fca9bc5a60451d1ed15bfba23059fb8ad7513377524f47c69a3e6f12792c655865099be329b8ac94b10f8fa778e2eadf645823514548af6fcc3452add7aa23d59039ddcc90dc605b8b06c7efc9dce24ba5b689b7e9a1af49e83d676dd322b263689ea7e4335f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cda99bd79a0051df2f3d453ad82f1b0662d270edb961dc71dabb4dcd4c23dfae66e6f3664998d76ceb38a4311e38c34f431a94353036118520b54f65961376d30bd8ca6e0202097fcb7680c31203d2308ae6d38ab6e730d8d5dcc683dc829157aa8bf7ad45e4f52ab891392c2016f0c2742ee57a2c0808f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191825bb87132d483cf729d6bdd47499121908d0c79969cc48a1913cf79d05da8ab67f7f5e64cadfaa5cc87835180506d48177b8e7ef372b05924dd1b8d7ab26a15533f7edbade7f2faaeea27d7d792707055203cf1e53eac7b0b0fc9519a9049fc33e7a9887544622bd338c1753d9b2a7e2d0aad910e7d03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc53cf11b294ca3767b4e85fcba650683e8fc5d3c06ad6d3efbe00faff44a810297657145e5300a1ee76b24032dddaa57e6f22bdd9b6d1c4b8c4c1c6adfcd2da10cd845134fb276d66fcc8e5fc466bdb05d6e026e23846a715039d51b4f75c4e2ea9a5a8c4a026e7d3552a100fd6a874818783ee0766088e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174748f9224dd43b286a41e173616f222dbc0ec8e281d886757b1ac55bad8c9519b306c676c040b9a352e9ad200f3eb5c90405e5bb7ef7a20723ef26acf5e89ac435e6f0d3715cf2c7e983fd6d4e4d9075313f6ff0c556a5eca4b98d9cbbc4036567de7dbe4b50b279c3674c7d840fa8130766621e3e632d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1317f4cda1942e15b0521cab667a6c9512e00cce865bc012b3b03f387ea620c28f980e4dfb3ebed3dd1080f003861b9acf61c4d8c1ddb1d74ce2804bccad12a11aff6f8acee36112e2b3908ccf607e6fbe6f2095bad873dba8806f8d8b96e16d0272a8faba86a814135bdaa4ec3f43c3eb273527b2ee3282a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f86d231243322987b50941eb6abe686d0c3ffbd5fc9395741f463e5dbeece4504966434d673972ebb23f56c5dcfb4c68e2e75458dc67b7bb0f16db79506c336fad363d5ef2077ef433fc9cb750235b154800b2c1b89b8ef95bcf810216ae44724ef42e9ffb0099d47ee7b22dff0abdcd0600b9772cd264f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h795e07a1423201b9ef076316610f904e6f3ddf516a65da9415b791b8da2f246b6aa63c923a879a6c19a6b88e3befd04827da6ab99556284c7089c5cb8a14f6bc5e348300bbb0402a33f59481e985467ca88f6eb93f5e3b52229c9e15a16c733870366b47749646f9195e2eb34a1e688bbab6a7c791b7075b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71a2538ac5013ea000df9927a3052d6053b6e89d74177c90622839e4f3fa3be7ad2c6039e0c06c31557ce1705ead7f259671914333df30fdbf850a8630b085f0ebac95e9e08c6cdcd6ea59cfa7769a8290f9fc1937e763ee87ba3e87677cdfecf55632f22edfd50dc97e593bc10bee635282baaad20a7219;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ebd378e3548d66e8eef29f4a35fba11e1ea16d79b5d35bec90ba96f47c5a1ee0e47024f6868f7b408b5fb9472181e8ae67c9774d150ca2375144d7fa2f7cd9903b449f53e297ba4d1d7226010c0e56bdb627558585053f81fa013a20298785290f5c2ee619c17d9d6926d7a79714f8e27d4678f499234dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36b51526a5470d71115f3e01ddbc110237f0eeea98fc28ff9bfafd327c28c2b03541c332423a43c9e6493aaf42a486bbf0b2d7ee9f4360fd2e20c5e910de61f7be195435ba9380478e7287f19ad9ae75f5688ae877da3ca30b0e5cd47f51d17249c1bdfa49487a7642ce5d8e9c6a890c77864ea79b2ba9ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43737b70cf403619bfa84c5abbd1c6e8213ee050d18479e8b010cbef2166e10713a53ac399ed4729e57db6ae052ea3a02d0ed3ae3a2961bd3f10d161bf1ba45c2f9d1e7728edee34ec7befcdaa4a9220bea87c42dc39b5890d831b825d9613b540b8f23230ad826700ffd48ffdc831a4194643619f03b6e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7299973304381f1b0708550a2fdc8ad7685f71ae02cc408bd688b49c507c688be96ab224319bd426c36561b70e9f3f24e68e05c41b4649560736b6328ffe3ebfeacf782f7ae9e5d514474d8eac005a3b251ea3e3de1751cc09b00098ad63abbc6c07d9b18cae1656d4e3db992d4e6f32c0947b29b148d6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d95f4cc7330664849e01afce001a95203d1b6261dbc3fe68b74bdc5dca975f22cefbd17ae213d5fbe88c1dc1020ce6aafec9380be6fe34fc51085730d3cc8ee7e04c2d0c839b07af75879b9b58370cd903f4a7c4c529cfc9d50bc86b2e01efd19fca40eb17dea33482e7d61d86d64c8c164427cb016612d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143243bbd986e7b723d6342f40ac655136c9357acbcdb32a4216dbb59dae6922c0488731d53adac836bd92f230011c5a0e29b783dbf8b624ba78e0628fc7906b4a1422d7f49b658a4ee23c964400db68c1fe7e371c8822f38f57e4fa397ff39dde195cced0abfb0ec4c22116fb3a91385d82e61e2c35c349a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1acf696fd77147e316c37c86a939376b2581521f09609e0bee8a18febd4f71d22f991d4cca9ba4b2f7db4f0b29e8a2b0542eaf0636e1957ba7b8bd38d65614f59a89be3df117cc429323a7084125b39a676b7f6299ddb44d2d8439ba1998636af8c15affc061d0c3527c540196f8e313f2226961ac06b3d5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16540eae800b8cd3fcf2c5e610e843acc9d5f7701a0ab63d91bffbbd54b4b85874664d5f5be0c92de322e9d063d9fd1f0c6762b6d432b5193a2f60fca297106cf1249b6002854694b63c6856cfb347ff1549884533b61e0724c7d886af054f9ebd1d213366db1731b08ddd9b96761cdaaef8d77b2c9c69692;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed942ee2032888c2072eadd7577e22c5b70d1bf06c605f031aae78ec2e0ff272dec58bcf77df433bc53083d9f51d165d562a187019579937bc3c24b6ab5e328ee135e6a9cc246d63fca2f69f9bdd9f41573ef11c4824df4034891df9ee462afaa4dd640c516d893420d12fa161ed1df397783d7d7749f477;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1355d6eb8e29c614de3e42e1ec0050f98649d6ccab5685e5619fe87a0edf1c0174e9d00734b0c0f3c62cb5d43f210306b1658acac0bc0c0f9ed308508c88e3da7421eb029afd89fd43ae355fb71a500f5f5118e2782bd1089e3a2c53c463fbf42ef08cbfde695a2cca6caf67178b8c62dc3f53780e41777f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1216e0f9fde73ce6f815d5f5163903545b8cb70da36c4d433b9d7e4e3026bc64ba8d8190a16b7d1e4959d86dcc4742a67fb964e7d8b860723f85c5b46c5389343b22d2554c206f00f56b33101b9fa4099323c554e998bf91829260ced942a107459ca589d1b3488f62e7b32111ed201527e6e0b44081d4470;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habba17685309ba38d099e546e80f8d85413730b1bead51505a5cb113581aecf319407d708d200ba4cbdaf62512b9f1d0af3593835abb1e6f49db35fec3fcf2fa5859b449c483514df0f58f67d4aebd41ea40879cec0aaf168a9193f83c4e3b62e0f7002ab8fc2564f0fd9839a8e9d643957986b84a87938e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13318b95422daddb1f661d999c995be0ba4e7fb78e4038b29fd7091a6e63b775bbafd74bd3e2372bad30d81ea15fd6d76b930930b64a5e8a4a6288d6c117583eed86655eb14f1a1437f328102ca6e3649bba34368a3c03c1adea005c8a1137879cf17cc1c5335ec7ab954bb106745f9001a9e81fe018c1024;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a07bd6952c2d483ef570d8a4187987122600510ba113ca8909cccc90c9a39c09be276012e377bc44424eb1a7b441673516b8ca989c4597cf194e15952ee01eed4c7a571b0c751cdc28a48729b14e1df3707e37401916198108783b4db816a0b3ddb34ba9a80c938a6f96cf616a9a7322fc173a91267c992;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c059ae2e059d00132489749ab7022b4b9dda8acb1bcf670b020bb01f0e8c1503833d67c468777263bd5860bb0a2d17e96b0b0735254a60004698d2459e564a1b1d4c54475910107ce8524b25d27bcd37a20c8f2765edd00b6aa70a040b5faaa99659cffea16eba3ac0b1a2ddd553561c63fc7406576bf2c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a0590c2b81a51b67463971d3a0100621eac2ee95c9799ede7f2ea6e7bfe02ba3ec2c1574f92d070d15eac7659571bf9736d0fbf0c32c338c336c4ecbc6db373468a0f245e8907abe0e29af083d85f282874caa686f4f5041535288f70b2383bab1a8b654b85007b4dd8abdd88776bb1f7c81f15041dda8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe67fde25d830046d6a87002d174769f8c5fd1f70a9f4c29b6dd479af2b0548bcdfb30a296c07931ce1a442680dd31baaf21903686eea90afa4a950f703d37b0b0a98e137da794c3baffed702266200b9ee9ea87f3fae502336f68b3b6d5ddf52b7122b162199440993c03e5e44ce46655b6fa44a83a53e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6797ed332f33e0d85859232a5761aeb319998b66f40a01f4b2b13a9a8181766d9b7694f32e56d492b3c78300cab5c83a8673c0cb98c0d6458ec09fa452a4f319cb14dcc3f2c6ea1165def0bd0239c66f906925a5a7661cddbca24fdb58decd17a0a3e8877d0033ff6469c5c3c72c084da3902d3287dceab8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149699fdeb42e3456cd65f5f5bfa5cb53435375f92ed2c771e8fce7facbd198d8974d2c862f6b9b88ad7f82346df1e84bf24ac89796d2eef3d5edffa8d04a40c75fe9b3bafdd595f71fd1554eab4c157d7ad5860ab1ee6695379a62d5bd2d456f0c36f1a14aacaa1cc1ecc19a5d53521e58d211ac01c604fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b07ca7c88281de25086cbff476cb4744a7caa305182ec6360f9f08201ad0f67451722495c7cf20770c7334f196e680be28c1b6c7b3d14a8282b37d45be28e39f845b55362d5ef56aacbfd03b71577bfdc94b4503efdb3cfcaeb00eb99108efcb79f55486d97c7e728005a15fc5b20578cd522529550c6d0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f977e8d8c37e90f39b908232d319881a9fe153be1d2bd46091efc3db98435049ad2e634cf54763afc35ef4e37cb8722c8f82011ac1a8c6496238641d7d29860fb61805d4fbccef5579c84b6ee6b1c5bff85bf114e71ef50116778a2697e82f0d4e44d08031238c2ab4b2fee9146143492bf24f4d3186501;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c3fb75db1fdafff70cb69c3fa5a787202be817461392511426e72ab8adb7d63d125640a4c6492cdc75e117dde86527745ed71ca0239cf260beefe40522347ebed4431fdd2ec58f058ae478afbba59f3c07c8a3e0fdba98a1c4dbcaaf4e270ec9e302694c503533e1c6c1e24c1a017a8516a9ecd8e8a1911;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1537ef3ebda0c6c1a0cd87f76230ee9320f5f77691490abde22b24b7658ff49fdd13532448942a63c1911972e902d0e6cebd672a0efbca97c4f801ed69b341e0dd966c53dfb0e823e8da14e592f1c0a77d4f37ab7ec6d01a292622bae188e20165e35fc801e5ff551a3d6949a93d64c1f83def62000b46236;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4bb07f8fb6256b3108048e314ba5f11f84881597c5f78d200afd138466edced345b700e0641adc19d533f0a9bfedd876e214c538c6c5ceaa9251c68d45c937a023823f020a32aff665987f8c6be9818f3ff9c3b6cd9abe7768d8ca4c37846c3a8cb7cf33f9c42b5a24ef1ae237bcc244b5f2a206cf05487;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b63384387ae9ae498079930a889b5f8d47bd2039f8e6190e6b51b4abf8c2207b82e79a5973c218482570204aac19710177edcdd6a3812780ef695bdabbeb94deec218f92927db776c2f7e89fa54baef222c9898057ab51dfadcc5b35c65367d775543aec3a46cc8b8ba6bbc85da0bfc3ed1937d7cee92c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefe377aab0014cff06094e687b6f392539c121c858c1b17ca9b32023655c64d1cacf2f3382f4ccbcaf0acbb8677570bc45bfb3e3aa33b596dd393099f62daa9914b0781b0a90a7444b807aa7a93995d55d5611bfaa65d6393adbd47d0e0dc50929b6f946ee29938e8fc83bc9c3ef57d24fd56433075c432d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e0ef61f8ee76b229ae0682debabf15f4877c00fd28026a5bc058b4a8af293dbd53f933b5ef4f75ab925a670c2215d7d073f40de84aee53794b8a28657b2854966c1a8d54fa11b7f909e5908575cc2d79030a65750ca542f3bd8b3793d8068a0d8f1fbc58c40c3e6ff5a507168b46e9cfd59a12744621c12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1928c3139140509bc1058e8b61affc6f9f1a41c395d923a95b09d37331e3185d7414d798826c0f11e10bb6b7c51b701bab5089ae73d49400d5fd43bf60fd3203a2595ddff76ea39d0da4344f903cc6c9bf8e19e62e99ef539873298f58c5d3100a17b228301aebf34f2ae8577d8bee93cbecf4caf7b63a4c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4bcad28f5c0fced1aa222b50235e214d225b995b3164e565906d9f1d753f7d5e41f84e9a1fec2c31eaf0a18780b8e22f1586294262cf46bf0f522ea8b70661304eea67e1f5694e6b755aed2a6f867f8c7d748ef13fb3eca1b15e11d4bb7347fe345c6f2b8bd78634ff0e04ace3ccd95903af937295715a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e833a5850ee3671fa9b578f7a907415bb02837c7ce9575f6a63c1144b726d13825bde329d63de860348354c55c0e15f3ac860445eb6c2c7efa97ea3f56a0fcfefce19e81c5db74f4c3b449fae3d0be80d74d80a46844a5e417e8ea0190f7be3f21da1d3eed3f68e6108e7d3b0206ba057267462d85987b57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd972601a7f02f59c7bfe37095cf191c32a8743502cf6606ad09b3b7d26f95e9b5240f8860b22815cf3db8568598596b7f6ec4af8c09a5cdfefb4e27a0ee7d6a1478397360e8b5e13d7f947ab85ca2abbe1fcd604428d541d352b4c4ce24844dc7597885028ad84292dfeaba2a2e1726f9a8cc5a2eeeb55e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44c6aa7fafc715119c07ce1b67b4ee13e0dd5cbe9afb10363b9dc9ae2ad0d9bd00b797ff3d1a14c2b2a29bc4dba905ce355f4b1bab57334219d2faeaa1a403eb61f226e1792c4c8662319671e092034da2cf21c3f891ebe7e94dfe691071f845092301712e2aa372a9684b0f6abadac1864ab132e4e2ca92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19eb05313eb4272518ee478e6ee2e2103ed9b1f1a73ffb1cf5a262713c227e37c04a46ddd53d97fe6f7801aa7f7d34e38a8144f2c5001e7b03bc7610f6b2487aa3564f3996bb0e75f5f83fe6f74e4b5555ce86a167acfc800c010f7c9d88c813e30bd0e3ac74f62ebe2e740963095aa112382e7fffc7badd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcdbfe83800ce78dcb24f0d1b3add57f53230d27d882cdbe39918820633a697c5f9bc52624f9dcd6a0c53843eed3c7f577a3e513be690712261f35df4930e3fc8650a72e266c5ab9a5390b1daf3698fe4f07ac6970efe39e42200e9f227d3fab47e7913acc08b40731c5c9f17fc8ca34a8d1e2868f2f7d126;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d47750fbcbd1646cd8b8bab5d00306284ea1e83bdbac5833a3bf978b6499d840525096083a85a712f17f80fc52d106d4cb203dd1ff3bdb510a9eb44d3601d083c692b1ed0e7d25c70a0ff3aa6f595896882a2166fe976430884346fc809887286070a8d264abc88417575e7b27eb93aeeea63f6d5a8f2813;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98bbabb6cd99e521faae24cecc0209a74a1120c0e5e7acc7c5ec2dfd062b4e6465e0265f4a6de3553e405be690febc66ce59881891e60621405f049774df13ac8fd4521a72ad63c0f3307fe5c6d02f69d74eb18b55e60f09bfd5f34270359a7d46db435c66a80268a91e90e3ca3dff16a40094b6c51946a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32d1bf1dc43c4dc16963cb6ed938b57fcc49100a8b67f3048d06ad6c3527bd44fa6cd5436129b60358b7d4b97568b5a1d33c3b78651e5ab3f18080a9fb24315d4c47ed6b30b480be43045e463db52304ffb711dcfd0b1a2dc6bb3fca2db12c9ae0e36c6888b23704a6357c021036df8627b94e032bdceef7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f2677c049b13cb8c7d3dd5ee6985ebf67ab9bf013ba0b28e56469d44510a395cbcb41b1b62d1e56c33dd06ea246d3d914575c3e47ac5983dbdf868444688e16e4b3e0e2b14f2209fdbf7a448763551bbee62bae2a1b23be012ffa0a4f29784a2cca29ebc31d179517db044efddfbdd0fce94cc3b902b52c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf5c4295aceea8fea484d12c3b8d45c9f5b0fe1b2a31e50d3bc1daf55479eee3a76fea989f5d8cc3cd8c6f01c093e7a720a6142277a3afee2f92d0286e628c3ef61d5fe7ce47e5ad391f5232c1a9a8791369b4ae36ce8d647005c4f1f012e81cfd661dd501aff82ed581dee7ae98eca520cca56fa7d11391;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da45cf34f4277424733a981854d4ccdc6a11cab12883191115f8785b2ac9f7f75db65ff994e5eb6bf3fa8385c12f1d15af454c7a52f5fa712ae18b355f5046269fdf66362f4e4761ad423edf8b9afb3efc5a964278643c13014ff6c2e1322c1f9b70862ef1f74832a507703b5e065863f62e6319f1c8b0b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196ad4aa136955e9f3732ac9ff4bc8bc9df700f78834cb27bc193d49a794de2ad7588f1595951c33686a5f5777ca8fe2c3589225912548bb6ce89caddb712c894d8c0d2ca841eda4ceca38e74f37631933d6ed00295dee20cd6c09e8cb9b069c9c6ee334b17c596ebb7675b07fe5e5a4e11cf3f89e7ec745e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf07f6ac6e4585aaacc1a2ba4d87e35b625de11dafaf3bb770492ee97dbe9c4761a9ca0aef7fc192ee5e16679d38dda3295908fccfe3683dd56dac34dcc8f3e3502e1ceb798e2ffa9c06c351dd05af85b189b9760b18e9d52c47bf7f674ded85a1bcf2b06b4fa0cfa75231eaedc9e53edb8b799337cf64b58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e01b30b254a6a8d13f0250091bcb4da98c061538f61efca792be7493a388e050973f5eae6f581de2e962ccb05c137b3c1c35f94dd7cdea5d74c25db13c59e02b537bfd41e23f380bc5c4c2b3076c27c56f1b993b605c157006a5eef84f74a826f781cfd323d987cbd8c4114d53e63a7a59f08a2584103e3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192f7e058bce65d9ed6ce2e387b4f8f57bc4d28113e52a1729e699c2a3c2221a9b29b81bcc93cdd77b6eefef7690328fce39f36c4e2c21ae538cfeeabde8049b944819beb23042d1deec44af284a8917b2b532f4b62facc51bbce1ed86f244b455de5e4109230fe22d5da49c6ce7acbaa4c5d1718c0312834;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae2705552927310c80eb576206bfb7dacfdeb14b25d89ff0b347afa4a240aa69a7d068c752a9bc030a24605a88908b360ffe85e716aa238d29542af4933cad1174274899704633a123272239224ba3b6735330ec5b5b6fff07767b797780e2457eb3ea6a0743f6d2424659653625aff4b914c65968dc07ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4b608e82f39879321a0505595c55a3066ede4fcefd901bc2ca85a3f14fa09e4a4c8b3e70ae6757f4309802995e8be2b0e1ca4251a9855a618750f88081c1dbc1c27114fc97bf2086a560d5eb17af9f4c1e9f9c6bae1e2e0396d7cca3e81bb74fe61881a84cda84674c5263f7cb51cc9b53b1d01cc212f10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e0017d528b8c34cf9281ca2966b28d476074a9769db409ea55ba00a91d0e7ff5a3232a32bd7d2382beb8076a6dc52f9005109a2ee2e84f07a1d1fc0104cd130d0ef1312e03803063497f0f48d15473863d8f5e381dfe147b5ac0c3ac38bf1de02ff55e82bacba8ea3322aa80a5a58715d18eb7cf3a6f568;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e3310574e195a505a6e16a4b349a0b3eeab2128df0b76054dac0bad616f3c45ecef2777373d2b79a55f8238c46499445ebb8f15a4a72d359fad810ffab251260ac67ab2704c2b9b2ad8dd954aa4661a3dfb787178caf7d569c05970e22a0803d5de466bb37155f3852de604ebdc7fd075bed8deb3c385d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc61e9876564569d909442cf33ab75c2d1243da54d47928f19b83ddaca9b3a19c0e5f8fee40c8ccdeee0f220f9c0470d75da529a1cb5d9861b759be83ebf3f25e82fed213d5bd4dbfabd7e67931d9b4b963107e9e6b06a4ba7a040c377f71bff0bf9a0c36b518fa2bc5e33c3659431acd29b6b1d625686513;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefadc82cfc01fa52270e8cb79f49520ee769a048fd09d2d26fb4032d0633f8ad6cd075bd65cdd19b011bdbf17253d3016b1cee22a3ee7273d7169266c6738303656574445bb9ec259c77f2c2ff5ca938332975946196b56757e5334096112f11f31d75692c38ea27cba32f56ed3f0cd2601aaecce10fb0ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142d87326738114e17c8f671f64d2bea43ebd963d225fffa3664d52f546add22f66c954a23d9dea42d9024db14342b0722e89d3ba73bb87d082d06f000c56bddf3f44733a5db3e5cfa272717523cc1ef52e27106bb90530da67a992fd5c71ba65e9591c775d0b704d1c1cecc76120358872aaefbbc7e15302;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1675f593ec4f6e6e16d6bb419274fd44e6114400e1f7921cc18aea0cfbf0f8ec639458d7c987f1a9af7db411aefb0f8cf4be34f1796afe0f0cc787d00ba783b6022c00b76f861c40d3af365b1603631dce0fb86b5af405244528fafc26115da3bfb06719be79cd7d61ec4dba1ef91b1271ef23404d26dc8b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f7b0bde5f81c8f9110e3be46bc2dcee2cdca9356aca4e625c1dba6b2cd66dfda0fa7b9436cc17777fe3cde2312392830f10c54ecb10883d71b612156b5ad3c257198e229c712bee4f986c298120af51924fc18dbdc5c49bf927102da2602d0ae30698639b0dd156c648a4eeb6254dde0b28ab203e6b96d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab64bd446f2d6ec1f8a415ee089d0675fcef8b899bb0a8cc8f686054d15da8e9a3bf5c2d53db9454bd6484002eb9378cd352922bd8965b67ee58a958a7f801719d65c9f8db30731c89ace105921b4942ad213bdf8b62b5efd1dc890fad259a1366adf1afa311bbe729938060b7b7157c530258736548ba0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113f5d7e14996a823b9b70ca2fdcd0744e502ed61d0602d6a44bdda47cc9fd83efcfecc38d37d4d785bc2270a55e7c6a2a3ddc0962deff6bc777697b50bf48aa20be8c8ded65911d8582d18c9475ddd67ad84f82f87473c5e7735c503df3483a4d2a61fe16e1f5bd9c1023510abcd9d79fa94814f59a6deff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162cf9e50b77a74991a5b6bed96bd63248454dce8391b93618418fe5490f18b2a8069f577b22dcf5c8e95686f72b3e2156f2d3248aad39bcdc85ee21f5745db03e566c3a313bc49bad4c353f706faf10255c2a619b09495823fa71580fd1f732cfd2e39ca241eba40951137b06ebed026bfea27bde17b682f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106be7e7ab1426ee7643ee987ea7984be505a137b3143776a6472bea47c8aaef52e723d2045733d334c155bf9ad43c082ed35ffcd8d133f32b1687e700ca16d463970265ac928c3b484487839b69dccb56bd6a30e49a2ea2b85c8e759f6584ebb257e98bb452fc96aed49e832780ab6c20b7a0ed0be74c21d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5cb23b1774863c862a101ea934ae4f6619bd0c8e4002e79319cadd14f9a4e9617b7bf08c251e9f0395a5a16e31f1a73a286a72a6e0a666302b85022591b5549af24180058f17bf1f32aae13b3c150af0031de1a51892a38a0415d043ec463589c3a680fe1a4a243b9f33ccc37f686e7c3429504300e91b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104b80f4ede0d8a8cbbd17cde838c955ef13e097b7cf3f089fbc282f7ddddbebfc6bfd5ec190143c2f7836072d2a96bd1321f149c015b03975bb54ec30fc78cd4c97ce6fa15c6a33909c83c58fa8682d5993a29673f86fe5281e79186599499c0ef82334d090b78d34b8e71dc0de3cc063fef7d1cec59405f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34b19ab7ac7d3aed00bfb424c3784b8ef33249b8df54cbe29b7aeb232c6053fae45bdacc78dff0b38af5ff14d7c87bc87488ff6c12e2dce63481807b0325ce0915601d79d0185954961ea70f3cffd3b6fe1a29ea18328e8e0c34750d9b75d3ca31683c7adaaba71132df207d6a69bc2b707dfc578eb5705b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fae0333bebb71a46dd41ee865fc70395d514ce30158c03acdeccfeead351204bb4244cfadcd90ac134f33b9b6b823f1d7b2502dcf32f1dd329ae70e9cd2f17490eaf082970163fb410e9595dca44db1d2efa2290fd361a41fbe17d012157fb49070701eb0c2ec1430e13dc3675d5e93a0898835e5e551b33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47de66a176725298b167cafe5c7a2993a550ed0efd781c863c289ddceb8566f7c80322c7c61e8ebca723101ca25b323b296fa467a9d90e9d40a64bd37ec626c72fea35e9e2d3d6fb20db8c5477d562cc5dcc8ce1edb00e156dae9e96339c9eadd2e6d011825328c4778550464482a843cd6e40c667b32b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc599e253c05a205650679633994ee6b2b1ed1a5cc9370e4d0c6a5f97dca47a762ee0bd00a769e3b9622768e8cc3df1e69cadd27695dc90ab5c267d899034281847134892912a3d70d1969b6a43eab280c0e28ce4977b3ce1c937e300ea51f0b16e8a37e9cf52712129c9e23d3def8a25f17775586eeaa80;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67e6ff06459d3e4df41cbf6a750ab75764a93ada0b0a7b9f8a2cf22508a41b42ada82d280a86a2ff30bbedb93f862099c267083cfea721f48b94dbee38b123794712a1af524f9bee74281a4ce323b0129a94620947486e53c9e0ca29f4fb70e7544f84e00f0197ddb25445b4b9d5a2f485df6a25c41edbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c6aca1a7742268621d1348c026612fd000492b1e28b83547694f315f608baddd26b550a40be60a40829ec775e1f1c28e645325dea07bceb24b415fbc02f672a858456bba7830c6a40f02dfad719f6a656d00947726280c81f757fa1bdaaac57a9487fa237dceb5a97c9ecdeedd8a1641a5fd275bfb547fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9254439a52930217a1e8aea0db66d06a0bebc289207a7fca253b43bc94305b95dab5ca8f682644c367f84f643eca55d1f2c8644b23feb5c9dfd43b51ee41b8f4cc4768da8cf3288d1c96231b12aaf266e80e28404cae8e45446d841fd34cbbad2279a7bf990cfa437b9859e27ff2b12c9871e944bfe2b40e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc34ab1b1d7781859fb511a576f8f13ffd4278d3858f73fc8e844c8a8637116056e12b68ed33ae627bd773cae8046f4eb6072f6bcf5e3af629a67c9b420c81b0f0ae12a6c1fbfc16ac240778416ad0b4f862f747bdfeb0bfe197714ad0643f7de598d902bcb173d217f8dd1e6cec7b93236deb715256140e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fc75360e0d449cd6ae87ed63c19deb60468bee76a43398bff086b6a5e2a22769dd955d22584bbe0c5c883b852ac9c8a6522f9b2bf4417326a27b2731cc7778b2047b6a0612f5428a71fd2d30ec2c0d763dd42a52a002649945accc7f50bf4561865896726422f0a0b9edee63c391c69ef0bb9ebc5a7412e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136b1d09cce1cfdadf49a7959cd1cf748ccaeca468f737e473cb5ca164fb00b5d7b2b506e52622d5672a143ed4601d485013e3c4c9b23abd0324d98284d6fe110e34714e1e445dfc4437488b1776261f8fd2ed1fc98d77c2c3534ae7538bb4391774c5c748f172b36cc6f05468478ca189c677963cf448f3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1147befdf4ac48505914bde1e7afa4b9aff1094918f86b1fe8454cf6c6659fd4e483b5f230cbc27afc6269033f2447df0a5b6a96772feda657e3a5709bb1dafeb18a81f88900ab510cc6ca2a73d40be65a227aa20c466d6d7d30e773b110d2757ebef5aa9fdf454838e5e7a607d91c7b8ed0c1aa106f7de56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha853606ead2aa393aba5a6a77df2b336e165e626c1e08db5fbbab1650cc0d3f72971d268a114f2c2c3ad05c2ce0c60e93806e12c339568417ae3a5f13efb02bf9e6445499863e2973a99bcf360328cf98261bafd34cc0ff9a04c5830d0b84b4193b79fd42bbf9f5e989f392a24c5f0d71dde98f851f6bc8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1574f2a2b023a74e953f50de95f73bb127729ebd1a1bb58ead5bc6b2f9c4e50012aa9efdaa3f9276fb594c03cd7270acf92b5f59ea74e63dc6261ed4d1f70d48c6a3a06a39b88fd78ebdf92e65c59355ac17f67b436398d20e9a37688fb599458247a6daef99e3de540defcd07ff5292bc61ce9e21c3b66d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc284521950ba51fa6794b9526148c1e78eeec915585b8a6b1c0f12466fdd939c19ce83655aa197dd4a31b090c9ed7c3236d0321a3f19fb433ee29aed8289fa852644f246af81ed835054bd21707757847b46a5f788e19a2a6088261c0914452ddd0d48aca61c35abaf149b311d63057c6aa38ce3312cee97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9621a9d39bcd7dcacebfbf3179fe02aba54d044ee06a70dd62900c4a9ed2ed751fce10fcce8426584581ad674b48c9551260503890babd91ccb65366b36ea783d24876eaa2d745941adfa4cf6606f2ed1f83f693d91ebee496e71bda8816b40be12deb4c25a0e33c05906f6f75fd7f829f579894ea114cd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf665807f8f4eccdee63c690b294dca1d6272365f37b8bf5cee88dcd233de68e812606c9d9f4b6867cb7a10c5c365ba5e5f13406284c4a2d68490b84f9ddd14a35e029462f3265086ddd0e01cf97aff4bb0a9c5bfd2db5958b8eb85466f88eb12bd371882136139d4fa1f4c0a98c5ece169bce24052eb2ff9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf646850dc36d4f2342d92d27a35cd7b1ed01c2490c7d4b955cb16babb10fa9341e778d0b90b3c32ac6f6feb657f63ea5e35169626885e09c7a59cc13f1013d9f6954e6d38bdd451b13f3654b1bb13792b6c0699cd5d99c6c6a4b5703a86314074376ee83769b46bfb6467f9e26b50f8d7db5b87333043ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf04682a3066cb8e098e31d4fb43d82cb4c04bd12390f51ca40bd98f3fc7edb222f825fd96777f0e7825c355e2d55e90e55682a2dd87de93338529af0ace54add3342eff001cb0c73eb987e05877deca3ca4fe0abfcc9faf9a2491f2d2cf619f1a382cb6b2f6698df39f56aefbbd4af4783adada15be1f69b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143ea14de9e7bc9bd7f4b07d5b15098e25a2e09c55d85341e709df73cddbcf6803b05591a8f19a9a208311ec1234aee5f446a8b330fa61dad6be74d586deb65aa442b6bcba82db288b34fc821a8b7ea72c2d94a9a2a99d89a040720b34f3baf1229363583c5aea62459ff9d9e85897d2b5f1e1899542639f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14edb9c99c2f1a336c6ea711af36aa62866f8f680c7e530da9d82c4e5f7ec0f5d73c75d30a9038c4d33734346d118436cc6dad32651ba256d0c5188117105af888d3a18c6562cc29152fcb1aa41ae89fc7798e7bf667b52ffe879468eb585b6430a785489419ab6fa4880afdc0ca0a39a4865ae0e04383f53;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6479ecaf07f804f10617391ca972318ed575e5f2d77298a0032c49cfc5468954423b2bc708550ef443e7fe577beb70ff02df5a688208408e28fd91baa27c2de169abaa4951f0e4a73c9b30b4486da03cdfd41119a7e13968bc3087bf1fb5dabce28323107aa85655a0920d047c42249d8a218286f2b494;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd79f7bbc6e58686044fd939836d37295f1698f6470ad6511bbe7324a209bad6bfff96ad9b3c9d361765b54de5279929eada14bc745cedcac06972dbb0a7925071056a686e535f74246da1b4e2ae046033f7b82c3674a2bc46b0fe90b91e811f4d4fa3baa603386d8ada5ed4910bda04ce14c8fa1972c614;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a233cec257cef520e610cf9d37a4350482ad8de1c0a531e785f75159c96d712fb4b728b01b032ff9e5ebb110625fe3346c228740946960b381ef32e9888f0eb3624e6feece2ac817523b2b7b5abc36c23d3db93aee076adabf751f22e4c0118894d2e4591635d798abcda4fe22d694e5d45b79ade6a96fd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a390e305a41af0f21d1fe39f7a036ab90a2a66c3b04f6245215d0cb6ac3ee801b8ba447e1de3e02a09d6e811b4bbfaa09637b29921c2b077b07f65010cf840e216e54347d35d355b135a498912f27cb450a42c56357deaa104192a864eec9e306de33a2eddb598be39ae319e48f15d44cc0531584391becf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104cc3890f63d651641fe377744c53a64c0847ad51b99977ca80007c4e45c98134a64dd4cb84b10e5db9516412691b23194d63ed9f0a88cd3d8788e5156dda84d9a9ec71c51bbd903a6a10d3b89ffbe12ed195773ed7de229d4e2b5d1bdd9b28fb98f6fdc4e129f0670e975ade593085688a8b21c243c3d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77188db9c552511e2b574295d32fd0bbf248174507bc5bab470a831827ad73717e89a3e53dfc022710615e65f52ec1694e8ab20eda4f4d17dd83d951b75cfa1a95a7b8195618e98feb0d9ddc343a9a9d39a3fc38a3ebd257378ee855af28aac9d1abe4b9c98283848b7cac310672f2cfd649884f7573c732;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b43d5c637f1dfb0a1064c285c7a665544863173da2be2a17e29685091406d87f3a4695b8bdfd6cdfe8f2f0a63e0c5258977836cbf3f1783f44637637931e1d73cd4a7c82de06a9309ff475e956a860cec0d3d35f08dd248a377480f851cdb836442dd869117bbc7c03e969c4f6dca8779d3c06fe4495fa57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9385cb38ff8bd16bc02dae59f30a9cfbab7624f49b8e5a800214f24ad6ca6836bd535dc069aa9c917aaae28a2d43e4f3a2d74311c4e395bfea57756f6c2bbab406e7277ab018a4733e27a495645d59f318e6fde1e46fc2f17bf30cf221fad2909d1d8e815100e94de018916cc6217c3e4507f6b1a6f1af07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c12b1fb2260a8fc0109cfb5a68ce077aed3a4915907102fc68c1883e4418dfeb0ecc681694243d1c418018f5b48a440d18b3b2917af94b5092d0d686137ca3d5c5215ec808a4d6d734815f51effbbecdc80d4ae0d5f95c51a01d020c9edebf56994db503f06e6e7397fc2682770adc2a3182313b7792d1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bee478205c797328ef5d90e3d4913fb66e2c47c3b3c37968b9d69b88e6dde2c20ecacbafae828ad8162c338b6999cc6a86ee7afb780191bad0726ca8a59d7cd8334a2fa7eee48fbed2e213e581ff13df7014d16ae5c4b8955f486d0de692251543e16e7a0ea92ac19f75cb9e6b501eda0932433a0a7500d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0380dedf5714bde102130145ed639531f42bcd5ba079f1ccb4da9f698a145d32ec79195b90f4ca2d6776e91884660c52c91657d4fd8f9aeada4787bce06563419cbb4a0903caaae42a3db8025650dfc8a3fba6a6da89e682bf2bb00a9e04489b0cef3a9e62512217c22e021338afa35d48f8aaa829b2443;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f105876d2c6b73a96226fa0f9b0c19c547b4d8914d8398eb82139d9208ff891bcadc4c6f55da1fa001960c715cd9b58dc151d12bd591bd9e1a41a2a09e49ffc0ec2a0b0d25e8ef8314f3dc5710535c72b3cbc18b588f7ce0213a1feec009aeefe64addd0f5aa43b388e78f01e5f50cd183cf70ae74914a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170666d036056cb08b0de073d044506c751a9802f827a8dfc4a9d678516982fc28021b0c644520a4f7b36b3d24a7aa0f26b2c4af4408567e84a80a169927103004afc9c0016ba52acef0bb1c000f870ce0dfa1411b4b89c3518b24ea8d62dca15d4637e973782afa3dbe601767f4a521d9acba46c38a80107;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f7e38eedc275e0659c5c175f4f9267d4f60ddb61e8543e4dc74b54fe5d1bfe48c0642acb4dccf1e69ee0920df403968817cc2a3f0307178f642712b7471a677401dc63bf8ac75b3e2b3ca84df740f9fc9a9e26907e69fb2278f4d2f78d9c48d2f0f69814a8d6fb4c5dd1303eba7fbcb0813fc21c2661f43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h710c2f5c6e3af982cedada2c4675413d9c3b037626af3b7ee6234363d4f1bec9e2db97d29e334bdbb29a63ad2d5fc680490d33a6cfcb60c72723e7e746c7bcd4ca2f947007890a9115cb004143ef382915d90ef2d202abc239870049ce0cdaeebb701ccc43085d60b74e1c9a064ab0f26bbc2f69ff0cff8a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da888ccfe6a6b16c0332ec8cd78c5b7904dc62a5f6d042997514eeec46d5f2f59039489f305f74acd7638e48dc90bda817a00c29e77515e77aeb175622bf719c08fb3f9fb3c86d05a8ce756785e3b1b04b619a9913fccb94f80b68df33182a8fa2b8b970e4359b3b4a2d42bc2b19ab33b12fa2b27acef2d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62661af77cbf7950a04ed918d9c8a398ffd5d4f9911e9b6a8145063cc46bb83111671ad8b85c8fb8f2633b6a8f4406bff07a97eaf9c9e7fa5f907fae42a9cb3a962f0b0363d9539882a9c22b8687451c7a3f80d985bb66bef0c5e9dac0cdede875d6193986fa190c3b6acdb7ec3bcbd48dd195b9a2ba3f5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189b22d4dc0c757f817ce10ccbda38e9ba481f4e2583d8807abdd4ec7cfe6dfdb02c9d102220eda5f8941156cc642d66d071b88b7862595d4fbdd0a2ffa223976ae38777dc85303b7df5ededb4748637a28877cf069669ee6fec5e98556d9084a84c9f9c0169c2c0f4192fa4342c33e289dec0f13981b4611;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1132f83ce6f078a3ae7cecb008e67ad77ad9471a484973b87157793d5ef3ecf48c611781a3233a32368843b09a175eecd6953e8ffec970d762b31b2a84cb25b42d0ff4d9a67688bb48eead926e1c430db7f714ba9e6eb5a106dbe01698234ec4e131040505aa9172dc3b61698d4d37e4061134f6ff08ea933;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d2a355251094ab7523825cdc81262552ce18085bb0679c5553457455cf544576159871ec098a3fedf0534b86177b0dc1fea27292758e971c35073ff749a9d8e5c74ebd091ad11bfc8aa6b2e152d04a3269ac82326d85e83a58d95b5e4fc3969bb3a5ae146717646b46f7a82f2a74b7ec7cbf9a7adcd7495;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13053406993757c12ca257e59d50cb074b5fb2222ff20cbf5fbcc164b38fe2622fa26b156d41f515a9c412b21e43b8c78f3d03188b9a012faaa7695e9adf9926e3e1e79961a873c17cc9c94d3c7235dd79a811af298bd7ff4c40d9bd5155fcbd9b853c74f217329048eed7c7b2f8563b18d50f28ee937da55;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a344111c2ecbf038427e2c6deb27a89a740a6cd4c088a5a462d123d7f54cf263a19840554dc2e6c3140582f0b919c1be8d993fd3cdc36114fe0b7aea2820731a6c3cf784c65d6d54b16df2abef31560e0bf18697b17357dce320ff54b09a91a81a0f7ef7e0ae68872c06649d5e3d4f8b24eb64e30c173b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dc180a65577b9c32d31e93086923ff3954e6c2f70b06cdfb734d6064963c6cbc4e65b822c5cb2a97fcd6410180b1d4245c6d375b857ede7c40c8af997a6cfc25d227126903ad46ebd030b676384a95e2c23763946fb32d94f2ba08d269d15e46dee900087a8be5193aaeb50f2c46cfe817f7a0c215aa247;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72ef8b32899a508e57adde4a63b6ca62bc1c9fb743d01abb9682157457efe8f592ec590b14b2fd4833a85f8846cc73671e68f5d2a575dd72c4491b5756f9963c4efdcefd8dbb7c40e43117197fa1df97bfc2f9d70d78e620634ce129abc2dca99c7f699823e8cc28542a83c94d4f97eb3640011f3ffc3e69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2a3e2362f7e8990a3325a94a0278ec36fd9f7aa72e892a85aa6db8d96820c5518368c3febe21b9a9247955bd51934b52b3c838837f2ed96917f67311bb0d89d930806ba471f4c47930312e624b5e37c2f9d5f15fdcf16925827d75370aa23271e6ae1785c5cacfa0dc71b8254d396cec8030a1f22db350e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0c843a8aff51746cd167dd603b926ee9fa89c09452ec5f42daa9b1994d5bf70d87cf454c6c320888840354b23e7f0eec6b894ba6ed24b754de060107d7ffb15197a7307f7958d5a1b85f938e11bbffead497fc097e8d7e5f4a7d774ebb584e08d440427ec594444c7490800f5a24c4d4b04a9d817284bd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61f83c6749f0d9bddb047d967269a0e81e825f9c814be0d46c503451d4a472f21d955e845190340561198ae7376a7e9c30d0d6de656c31cba52381df4d92c32877154ea4e5a64cb1efce40854ec6b586a25860337bdd0039c826099f0355fd265a8c9608ded21c075d1d9ae7d5222d42680d3994a783d1e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e372368c580211e100104c526f9b23b37ae050038182b03803f1e08eddfd35cd83b0e9ff6fd9edb604136223dc4ed1532ba0e0df97975c15b0eb44b8f34d1984a46d2df0017e65a0599632a9babb13dbffd130cb7992d7b34434e5c39e38713e3d16684d407cf412d038bda3ea17eccb5c96b57f2728043;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h967de53d329de245b9d816dd4fbd387b76e2b32f5230e5b638e3018f1cb431ceedd16b3d922a3f1048a6f150bfe84512a90056db65d99fc9a8940012a1f35736edb87d5173b3674cb64657132eb37f4c2b9b8003c306209a8cf849908333316d6ea6ceb8cab9deeae3b4af6ff30968ad3a884828a500e5c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf101210b3ce5dc4dfa0908b6bfe39bfb3c657f5d17817df6c4a1b5922e6fc07b412b77ddd83bc00b1567573068e3104b1f95fd184b32e0327c800bf24fb692cb21669ac6f743cb3c4aa64c147ace0048253edf5c66a6fefba44c819471e04f876c6f32f8603ed01e15bf21b87742d8adcd6f69fbcff5356;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc584e769d0b3951142db5351240a3a25c5480341669f7c6f26bfe47ae5f25a5fb50ef78b2a978c9f580bbe4eebd320cd1b97d6c10eb00d0de4a2b4656d11ca543b16c53c563f85d5c41b8ab7e1982bee92db6fb79d9cc15b338fa33e6645b2daa8d4a3c34267146866bc15c7c28b3faad777d2546173d83d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19dea6b61f9199dc525ee8109fe34909289c215ae817867b5c943813081593642a4e88742b00f7f3569cf181376f6291315b93d68264b28862871fd845e17ed85f9de00ae8f486d170051140670bc682589f52a5918be10c97ce8e608bb570f2cf4801665a50e79862585266c76334b04c3ee96e78af2a78a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aab6814800cd9fd12a94affbbdbc468a35050a4c44c8a2d14604ad6e8faddfb7f709f58a034b0107d8ca56597a0fc3f6ac75c9f297c4754b75a3c8aecb5f9ee21c04a8f8b7315b15b613d114188a5429d4ef3ef9da704ee13f7c48bf6e48c06102a1d7977a3f21665a12b631739f730a0e48304027a29f0b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128da8712e13f6253ba3e4fd295e3df65e216102a2b3b4e510c0cae56bc9a8ff262308687f5d24199fb2aa93d2d5db4038428a8c1f9a5b50e9431e8250086dc5f36a1f4fd6973deb309592ceafcbce4fc62bc543d88ae5c8ed3abcdd4e293e1b4ba0ab69435f2453eff478eadd5f7536c3fdc67d9d42bb17e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebbb08ea5b21ed5544de78db3be74853adf546069a51ad509bb6cbdf84ac4154cbe17b46830c88bd18223d105aa1185746643a04c43601c59d080a9bb9fd289071968c91a0ce84d0b9ccbec612e20e2a84dacaf824ed7f1e7ee36a3957a52233a84bb42fdf18f50d96342199d816557a4d34f3d110a3d2e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15201d003f34ccaa30bf518faba53de55f443a496a3a408e3c012de68eebcd43b2d85dd4afe9ee32f333cbc7dcfc35fe50cc1f4618149bd48443474f294a264817e61cfe6ab9db436f71d2e498cca738659e9c1e3388a90bfd63ccdabdc4fda2432cee6580c2be5126bfca373c907256d5567fa7ee9927231;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h914b44aff471fc9577a1383529dea08d1c58ce52fd64d725fda498485c8bc04f1de5f0f6751c272d51c5a922370c7d7fe97c0c920aa5666c1b83faff0b989c3e5b938cd5793aea7f467603738cd41e1abee3b83b249abee4545ade32ecf4ae9b803b53077be69dd43cae618b0f4b2f14851574861f8cb13a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf47eed8c7e51386f44f1a57dee195d162191b04f7cde8109a10c855e8c7fc2cee2c6ada44bd38f30785dba324449026b4090130fe1c01ad4b96b2ff647a66327bf7730597d4c64b23eafe3bf8448b2da705b367777214e2a451fd8912ed0b0f36371f68c57899c3c406dee3bcd18e781c9087ad57163883d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50178640c1757d9dc53e3fc6be47bf362051bf2677e4fcf7b7699c3ab17cf7df0ecf118022df2e13b56e37abe4248738742ac2374ae7e87058a3aafc63724e7a22444679c156fbcc3d97c04ac190743ed17f50dfb5f76619d97f0de29536d62309e5c232ccae74504d96b32c08752f1fb720fb95059baf4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a2c5f1203ba22d97f181d16b73b8310c0b1cf8236700b206478ea62535a38523737c71eeebde94471d59020fc8fb03a22712c9d33fa42ce904082c980b06b8955c02ce979923bd912d5b8d27f046086e38761f7611991ca89fe83cc65fae721e6c05102022cb5d2555373bc0736d18cb4f6bae069bf40e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13725b223d8d4b5cd1f52cf44c3b8bcc4c492d4a1b47f26ddb3ebad8f116fdfada47792275de2b2307f92a13d2b1d7645dbcba1c75fb40876681e06e1a9b229c6b6f531799c0d1a88e3db90b5974cdc1c271373a5b2d410146c51779e843a5e329741518d4c25cdef86cf67fdb1e243b959d0de4b2d221172;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165c09f1edcb5a5d2ad361a407bdb03e03eb29395feef0e6fa119c511b9fe1181e2e278eac943d2a296555afa342573a0f695f721ea2b9e080d899238bf3e584fecbe8d1709ba071b3e02d92499913e68054b2438e707c02924d3e5f42bceda689b4ebf5578dfc85cd48f08db71d8aa0f0586b1e5b5bc57cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c551fa745400b5274c577f7a3515d3bbad8bbbb14b6c26269023675b324cc44db4efefc71537fb79da4ab20be443418bc75e81239070041dba8fd6472ff3da83f58beb7d61096457575f5410543e3d0e03802c864dd5a3bd5f81a0ece4a46971e1587954c541c048544aaeb1f7f99c53248d11d232c4253c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb927b852c9ebbbfb2eaa924f8e3a52d5d262c6002598c5b7c654b84362685d3ec716e11ac6b172dcbf06c1173970907e5b694ca7a201010c796205fd6bcf199de0896bda55a320799d97382610eaa06b143a077509283e7b4d03381305311c3bd5b113bc388edf1f05aac676dbd1f000ff602a5811136950;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f33aff02da5fb7cc6b2f7c3ce73e457d5da0c10307481f196ccb07638bccd5ca36338e248a1b1616d7aed92024c898309f9ca3b8b2d40a7427b37cb3efb4302395c73ee4e66a3e95de5a487ce1896c5d59a3e89b3c0f23309801882dbf0d421747592bd51a7fe91f0a3ad96332cae0a1441127ad0519f365;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e02fb51a65d5fb0def7aa498d2314f0188cb71c60891e39e4f5258d83aebf805d381f0caa5c6e5afc267a4a242646f0540cf91fa88167b07447f20abb73dff0a1ac63471190b45fcb3a9dc02fc4a629a6afb51eafe618879d3284a55849cb2ab09b111674195fc8aa86fac2f6ae10fe3c8577ba234288c40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h237b4ad8934022736f0fc1c2e606267cd2d8b726870340dc167bfde233efa81ea8f3ba9b3bd59911b7898285e568af8d8932a618a51cd92a6e198c618db7c808864f193110afc89771db33b57e0ec57c7b835b2c7f90cdbb83755429fd201f5747b25f50fa55900a9b313c64bbb52b65cd032410e7af02f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hffbee7ebebf0a78646d6071ca4f6b7eb166716de70219dc4047c3c95d266a9e9a9be2374d6dbd582632373a4535d2c5a8b34e9f58b1e4b6b9ed07b926f73ffa6bdfccf1dc4a87b0e5cb007efc757d3d1831028df8ba157db9e701f7284ae4fdee0e732c18d0e2519c1980fc527636949b703869c610c4313;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3dbc4e7341bde5436886db30f7885efb19881b0b90f8054c91193838efcc081267e052d2f3b5d2f6f4a0805c5c9f62bf95192aa4b92b50d906c3f94f75f5c00b1a6c12941dd6e243079c605000122bddf25b934f83c557c16759f71278d358f652a04c73eea53a0621b93dbeea55ad62e1067c3acf4cfae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc7ce90f3c5a6bb9cd614785a490bf667f2612d429a49c4afc395e1ebc2b3dd0f5c3e97f6931efe4270281cfdc3589bd8bb7d092573d705fa33da65055cdc2819fe916e08b8f590acb00fc849e7e14175c26ae131e8e8aa36080d17c8336352cb7630e7866d645e7c911f6f1da81aa75d97f305c9309957f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce57160e7bc7a6f26688bd42c39b5bd791e0111bc87384dd7c57124b5f4a4fbd9ec8d1e9a62733876645e84bc81fe65be61c0e3992efe175b170d6eaa5929e165d5e4a4d3a747c69207b1730eec01f20259c872ca45d65bca336937c4fba9d2fd904aae23a3b3be60907496830ca5a680399206c29aa1475;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1397a585e0406431f57c9db1f83f105b763c16869e131a5798ee6a38a3c778b02650e801d1c37ffb0ec7104774188c97d7348fde6bbd66a88a4be4b048a62e85b15644906e93f70def1178391366673c86cb9d9047133c304c58df892336ef8f151cea5178d26ab8553f02b72ed6de24ebdb59b9dcff45bbf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1807853eed541ba6e87cb3d98842957d8bad3af3d3575efe9edd335396ec68e98a4860097e7aa269d3a742517c7a02f68f191d6b51b4550dcee27c20dab803300b01724baa926e5b6e3aa44a40c4746632c6f0d26b0f3b6417af3d143822f8da2b2466234959861dacaecf7a810cc9b736f782a2638a1b4a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2169ba5d2d17880425d149e04b5e293a31ca14d08ec5e92d10a859f608a4c5f74327b315aad39f687a1305fa3757f91447a5d19583f122c70d6f666b43767c703e7d4ef442a68a5ae87e87936e4380c7d55a055c82465b35335895091e0a616367eb8d48c607cbbc5f2a17e156bd1525ed8e24984267bc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128c4e4d581c1ffb1f206887c1f8642fd57ce8992d031cd355d712477930482127449dfd15b8b9a617fb84f48847b66856111073627b9eb5dbcb1f0902e2931bc014c19c978d6767647f139610d521094ed8f79b67363dd71175960933ae2348c1903afb02deb68964f88e3d3a59700fcca65d1db6009d997;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9e4d483faa00a409624c3a58ad5eaf2c873ba8f23b554ccbf684cf7fd52481388181be8b86f2f34973232fb1c1dd0e7bb5653b10d3fe7d3c04d5f9a6a8f5e4f4b93c8380da740346e95131045e53be4e8c28faf7d1b21ce4d2413de42d03fa6e9e598b2d8e9d5b70342997d0504b3de3cfbb36a14062033;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6b208da6a0092fa9c5848f28b61101996e610ae9cdaa0116f553b091f61050a1ddaf2a68c59c1e45daa0e6e7e99bd1697269662bf2c77ec584af672203492e1eaf9f42b6c4535b8c87bb31f49719dc59abe78ab3d1c1fef7cf2936416a5412aabc01613f6102d236f134dd4cb9a131b803d2fc8033507dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9cdea0d6a18aa20630a6e83f4774ac2921e885ff19223bdcd1601341d8f36cc2301c2512f14e42f6e4f9e98913e2c7d70bad597bb1466ae0fbbc76a75c5e82e35b2e7702b241fad3d30679a0c445dec8659e81d9b20e9d70b4f14504ce80d2749295797c208fdd5951d977dd2d90186e254867350afb9ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb387f89788669dcabe42226f19667da8b0c9cb92157adbf946c784510801e22fe4af67680dc5a9ec988570b1a002c1115c9b12fa55f090580065c2e97068a81b691894e2fef5acb5596d5f08d0a03ef5e413990c102299a99f118d501c59c9879a71d98e51fb732330f736a45bc2240724af71ca8bdbebe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b83f9e47499a2de5e876c7c726a55256f2cd6cf9f287db15e032649014b51ee6774ac464761fecd45ab0e69bd50c96e1f8359519bfba13254db459d19d37d395b0dc3b9624111c44b66f28b95dd145c1c4c8fc4c144f744989a7dbf636c9e8ab727af36a4a5f544b8e3de7086129c2e6d7f57baaad50d0e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1661c46436dae39c6313ddca4a17b501263a5e03fa2117737a7619b3e336ddb5ed500193825be04c012f10658f9eb4708416523d7ddc0bc370d083e61dcbae5d98b5196516e8bc66ec3fb6b78bc6f39a8e2ab21bf66d1bdab6b2635eb053d8b5118037136759e6b19e973dc90bb2a3622367c9170ff83a7f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4137b432f2dcb95ed61562f306b4ff3649e2690781645203a060cbdda1c02a5233cb6b8147db936609f5a952e2356ec7d47d9724fbecfc7826af34e321860be393b37873bfb45d9488c0a6f56e80d223ddcd6e42532589acce72136976e25197a4b3112481ac81998e65b4ae867f64259b63d817a82eec6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33d78d2da9eae2c993a16d56cdfa680295e2ca756bd926425343f16b6f7b76dbe6bc01a1c1b5aa8a19ca2b6e28029bfe8f3e149910ed0c078dccd8bf1553a4a0179192c95b11a1c85636b5729c859aff9fd9fadb9bcb5044dadc3be5a21a629ecb6a96d370e4ea754ffb41251775ba5723003c5265bd42e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c6bc5fd57ce69ad06fa8a091aea0e6ae49ae5b5a783dcaf1a4a97afcd6fd91987d278f3448d4294e29e6a24d2be1fcdc74276994fbf0d3a9daef1ff918238256aeee2109d50e10ef48f71a0dea517071f63c4bdc2d795d68ef8809c7b77b8d66e664a0a60de8d1331254149fe72b2829a63723aae44c1eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50c66de5b6b212a483bf6829103e2816b64c2f501a115efd09fb34c2ba24c7eb7842db8c32bce9e2bf14eaa3daf171619260b9f8699fbfe2c2d84c84d5edee8f81f36f3119196e18e64110334052beba23b5a34f781a0ed9a95dbf8f449e955b5a72abf2200f160c2a9611dedb712e50e927e057bff46db7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d5c20cbed84e2c8509842921316d2b4aca6386370ebcb3b5ce6a8119a5f0f8c9dc4c126e8456cee790f6fc085d5f1ca1a05bc0c2a851a9724418929fc0e1bc70593bc317c1bc3b3ddec6513fa2068372212f4b1b0897145a69b3663b6f7596e722971a33be65ec6e8400cf049ebc247740dd0f38277257f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dab787e9e1f368011e9ce604008f1fa55302ffc7b9676ad1bfa72eb709aa2711f80af0672e3ec66e24f05b83c783c323cd21983a26b433cbe5528057f74d304d2707c7d805bd9a68091ee5b8d58a0e5c804baf18542968b16b52cbcb43937f268b084365f8c49ca746ad311b7859c28d418a91eb4980e89b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11eb301d225afad9ce23682fc380f9a459b56bcbbc29440649d65c810bef1625e3f02b7c4f6cbd4f5638fa12abee30478331270d59f13c99ca5eb97da350ccf284c8c90cc1292f8f9a3aa2b5503659685d28fb2d9d3e1bf655eef8f04691c464419c4a2e861eb96d0a8679b73521620c008c26919ce795424;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd43ee945b838ae97c4ba6e2a13120a0b8dcab88d3270d88e1e28449c6d218d5c35a3d737a13d4779f693270f87c47d323a0c8907249931e9e6afb97c440ceaf0a8c350b7e0c170fa334c718700e6d81fb73386b9016c9a12c622af4173d9acdd5dc907ba422123cd50480475e512e928414df13aea53545;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e705f1d2993449c14eccfc7e38f844b55026fe3b0fbf5defeb106d72bcddd5328a91bcd13982d447a64e67355e3bdd3ee3fe7f37c48f31bf2ff8bc71403a80943b64dffa1aee9726f5d522cebc628cc58a450d6cf7a8343518c7acae46e86a203c199af3d54596ac56129a4b3fb73a292cf2231fa4bfeef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bb788a595eaa4a2c7d4c31461d920ccf186d93fd56e3670013de774c609dc373d0f789fadef5729c944a7cde627f272f0daf50fe2f61ad1a6e8e14414ee54329371de356629e363cfe62d1dc18406c4d339ba53679bcf96ce9f3d5dc65e19de437af0282a7693eef2030c2adfa57a014c5a417d0b5e4dfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf86644d9d37aefac17b9acc3f8cebe3c925b3c6ff2fd2f33fe558c3f6c4c1d99b91611520b9bc4bf114f08a348b9eb47fd27900f164b2b6f23b773caee1173cd200ba1224d3f9e03f8a4f2d25f033a5a2a519581c143003a3f765241334b4a4893a79c53760a1576deaf864727a071fe017277a5b7bad3af;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afcae024e2df2d39725ea1a183154c60c775dc037ffa9018e13c1905a5acdfaaefba2809f352997c32b472c19d8980b8099b8398ad0032f7e002946f579684f322b030bb1c53197869eaf171fba266d623f71ff676bb3959174de9eb721431c4bd45bcb38036d6956b2c0bb9236791cb681b0d553451fa89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf896c5988908c77ca6c0d5a0055314524a0614043b0d3e378a57e614ddd1106d36ca823fded8be1106af95659cdca9d9b5633866dabe9081aeccc8dbd6e7ffc756440ba022ac94482ff509efd9423ad475d05c2e46b8d411c89b6050629ff8f88016d1883940bf84481c8c0d3b60ec83fe945793271d7db8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h300e8457492e796fa87b907152aa93f7505ea1e4948940e501b85c8611cc96e4fe169648cb9c6ef187d5ee14860048b23fb8ccbdf400f526c5603281c68a2a22be749c0ea4a324eb87cfb1aaaf63b98ccc69e8b36746b2519f5f04b1baddffa37f467d310fb76dd23e1c0e8a9b9984b08c1bb48e2f95b06f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137187d7b6d236f736a6d8d8c1e6e002946ad3cf40e5bca9514421be21696d6cd38ec88a70fad66aa10d6c5cb1056496609c533e9acf377e078315c1eec54d1ae3dbf535b7eb5cab79ec1dfaa4edd90c38ffd8db69228d94b50ca8c1146f3e889ae51943388dbda4422a7b8f495c62ce418b26560af82529e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c691b272c50a15265c3a252b3bd7991b9ae93695726d25e8f91ee9e0d48dca9ca3d91fa1b595b9673bc5673ac6ccf44cb4dde537bcdbdc8dcc2b96db600744dfa829cfe617bf67684be072c9483d2374e7607af7ec7f024e0fb64fd335160d495d48b0350d6a71f9fd495efce46e306abbb0bc7421077a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1373d41efb7504ee69a9537272440a6f9b1f5796a9c3ab1d63750e36cb8a00b770538c9a2cbb87c60a8b9aea71a8910cc3b23a74320f126d29b09c1c618742c947b49a43ec8ef16780bfb0802cee37ac95eb0042c834399f8d5cc2bee1ec1ca1cbf05fd6a6542ca233de419f62d57ca07b0f429b7a1d4c926;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d1320ed81de11b7acb737151b051300e6f21e2e90c1182dd99f2d5659877f971a0e73f74aea7d62ef2b6e45afc4f04ca733ea5b701495411c78dc94eead22716379afc2f5f04c6642f4a3fdfc0b0a26ee8faccc06bdf18bf5bedbfddfc1a910df3fd1e3474ac666eb26a11953c051f307ff6b9de0fea115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5ac62edb80ef3a2759810ef383cf32d4c353c9ffd2cfd235b5a75eaaaba361a44639ca2e35578e4e8e31b7de5e9fc6dc66bbebb08bd48ad3a080f984e2a5549424ab39ff72aab718311a3814c5736060cd7e80775ee51e179a1c26772890f422f41cd038d5e818a1d252496368a727f371986289d5ab422b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e65aa8a97c24afe16d37dfed6ac2eb26064784f4d8b5e7ab9893d450dba9812f04e21792508cf97c2dd62922d937fbc1188ad65da9565e62c83ad716f2eec38eb8d497486ded1451a04c89b4e8a09c925ab3ccb32d5eedcc81d08f37c029b5c8eef565678fcf8e076f463baf5b92cafbc0991c331161935d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h457eb284b62816efba53acbaed1a527f7a9646ff4090d8cdd3c7ffbce717d963a2c747646834095ea4163d6735f9afaf97057597f4531cb485d316ddcb9a1d6f4c58ac9873e767455558f773ff9d4c9027d72a22f03d1c09abb74f0088855794572a408d7b62e80e6eba50085346c1d653157931ee431d38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8cea58a05dd46da65e513a0fa5eca44589f69398575d03a7cb6b7dabb301f4c0fd56fd1f7b2720f0f62d4c089a5490700bf7247a7f58efab5967b14620107547fcc2b18b2f60b3622cec5e9f4f28a6e47713579e1cb70a907d85b96e1bc1e1a79e4bfcf33c0452462f71bd5dc500dafd9339d1806e96580;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0a7cdbc1f1c46807bfc042718a61f5a54d6e75452f902c8425d22678a2ce6086764a97fe59c3b31c4fc0829b7fdf002751689d12ba8bd3583bf8f3fda7bb4b1472d9e7176275fd03e6e24880128e98c511a25d96e63a88a48773f317241d2774b32b5463bc5db126bacf9db55d6e91226da16f651c28516;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2f76f3ed5e37238bb8bad8ec8d8b781c105fe1a8c58c111240edb861dd231d7271632438f6e09abc37aaaf603ec198235c92f8a7e99ee0fcbf353c66a316b1fa22b7ff7d085ac22266cc7640fb7953f75ec47a3d1a01426ca240864b5e5bde04b976b7ae60996c70517bb044dc63f931e9e4aad05825b67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71e7623c46e0309d7f9f4356b50c713b06c4019051b6367b18b390b80b85b6cfafd69a13c3bfaa1c02ba999064ca188dbcf5289f26bbdc0bcbce9bef832e137db38b8c12c10afc75fcf8a51ace684dac93e12a58bd921e593be4f492bd3c2eee6630832bb226eacaae6e0bda05fa82576138584ec6bf5ed3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h657fd776795f08e23958bcc9aa89f209394d92be66cfe22f679b68fc4ad650a26c3d77f3c013dacb9688a96024221d3d87d3a437ccedb973733d44518cd5105e2797a1d71fb6285a272ea4013c4520d612886bb7d64be8902bc189014cf49120b637619cde4d6510e4e347c4394c794b8ddd00d139bba82c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h660e78d72aadec580da5dda49d10ff328fd157bbe758899fc5a96374ad6ae8394b202a81d3e41d561ed7ece051432cbcfe6f846a5c57e5039fccabf0605582ea9822abb16d781f5dbb71c730d338c79b4c19f3d31882e135d8eb2c20a9fa3d3912b021b949da9a6eddecd1c0966ada88e30d531ee027cc0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130104f9abd4f59a5521d7d22eaea0ec783e2409fbbb47ae19ccf1166936603e9dc0d8db97b2cc4f6bd5fe11c7973f76df7c43ff7893a6828cf0b0021daeb2c103aeafd69a6d3cda33d5fbe450b3bef32d8a3341cc1d189e1c2c3712af2868625c570f6aa862042624fcdf5e18ce9d95ae8c177ca6a7d8949;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f2c864218b0a9ebf65fe45ed6195bf4aae8f886cf5c23693ab6a5f05e881cfeee3e1183d3729bad89ee5ab5cbead974c08e74415d3e61e5718b9f669db5b9b4b378f8b680fa9fe93d398e2c72b648c7ea12d790b80a2ecf06902bc4da278b467e5011246baeb5821f49da70665915351ac666db322bfb31;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha538445e4f9423378cc95a966f607470b8d413c091901bff68729343946f71fec06591d43568eb9235c2a9405096090397b6e4031114134febcc69ed95a7d5aea6b90f4e7d5d183675f7ee0953ce9c890e61741de588210d07ff0b37d152df24994e3c4c2cd5c9278c33f743f58861ffcc1f2db0a2076e01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h755c8bc0a7712d092709a2b9f3e537308dde1c0ef937c64ddd3b6cbdfd10c9e29d30863f1de4572e4c32e9e8540faa4ba333eb9b466e4011bdbbed0f60a52391bbd9d9d6c278db9c5b96ca9c591f6e27e0b4d8cf9a933d12572f8d120861c696cdea4785c3c42817583f81be1989278728a0c45964da7a2b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d063e4d4573f06a4afb500e4e721fbec643bcb19d58e5ec9d8b0596f2e71c03d885a0f12d7c4d711deb53c6d6d4e41a92a032efa9051d7fd775237c059a9c24dfaf17636b7ce8ec70f16126cf337561611b73825033ab5943267a778d45967cbb8478974e994a7f9387a04a15ddf3951ecd83b1966720e9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca132855e3737f056968f87c19a7c9e87ff6c77d0362a5e8c2a10246f1d3dbd0e243a8cb04b2098708fb3a5613fdcdb0b411da9e4e0b23d1d1b1637d7145d9664a5147cec6af7e52e2ab998a65cebdd7e26fcee1c842969e36ad36cded75ee7e4f6f0eeb9403392fcf6e62da94b14f13010a4447c1b72b97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2f7d13a1dff9dfa17a6ce63b7d192d9cd36122756c42dbb1f678db07b296a38ef8f3a0566e28bf82bed84d02cc383829a2e5138a942826d48b34e65454053e9202b5ed113acabc8219f6e887206143febfed66c6d8fa6acc88f3b06366e39324c9f86edecea5a4a9a563ae8e70669ae50d804617985058b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cc55074c4e4044fb4a0f84d774731d8266f8912639dc953213f2a5f2670daabdae85d98eac4599a7fa5cbfe3dc80693410abb98609cca666a244b4dc58ab7622250ee4045dd37f303dcbed7c408e73ecc1133841717406f1c487d1771aca341390dc86044ea37287a718000ef9edb13a6252c6716061bb7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b45e5b8fef83fac8ec1a36cb96e52706484c234f6d24a694ae1b432ae070fa92854f9a4543416fb6bc8f38842729407895828cfa0926f6e248118c85b36799f5d6b023883424c3e2bca9696408bca59c25dd3d4fc0ac8fe0318067fc7abd8a0f29766b8bfaf01b548af964a3d9987faa598725acec90084;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f7ce4a1d6984c5356fec1b78ed51a6801b75b2db177864f816651a087759628764751f688d5e4d9fdcd2c36ade324d879509e43ac1f3c195dd36de6ad092dc163266fe230c53c7c77fdbed7723b0aee971de1b33d1ad5f93376657ba58c352283807c02165fd643c9399bb09f955fef638a5ad311a2e9b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1baccf69a20ab04a53aa926311e8efcc93dd70bea938c1415953bc98db31d70fb695042d04bb95fcc1680f2ba465810923403e85731b3b63f87e04fd62f63fbe5185be9253340e8a07ea439afa9bf0e53693b2059ed8520536328c581f0a263e99a16e409913a58908f4a0bb8c4a2ffc49ca0a96e69cdd5ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h675f6f47400726f87ffe5aed25fb928a5e897a01a9278c47003b2d1f51aa898896f6c86520e8dc66f40c92469151068bb6b2c870bc1e85bf021f80e9cf0ff697ea4146fc01a4f3bdef2582f7cae48ec651a3f825c02169e6a7ff1e75ed32aa1450047fdb03f8f54106fedc0f0917cab76d73a4b64b56a307;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc87777f3693c067246c62f014825ce811dc192c70a894070fa204f5669d23836762ddcdf497a933ccc4d162d36da7baead7da5eef3d2b9b448ef7aba589d9139602471306b1cbbe95d788dc1f320cdc3aaa95eb4c9468bac7620fc16fbdea01c5c4d6b01adcb5b6115687b64bb688ec320e370d52ead763;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c2ec27d73c90e6a21951c4b5ba19b9f435033d3f8950e529d4ffdf1683b395fab793f3d5e7b0c26d0cff0f4bdea83d93645c44fa7a9c30a75ae30f057b5f855219f0386359dd699f52e285bae137c4f135c0bda1156768e65763e1c60733818e8a25fd1dae21bf0d2646e2c0eef6aed9fbf92c35070cf8f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fabba49f98d04931934490ce302c85c6a637dbe1e182294340d80b31de71234a193926098d35c1bb110c898310f5b04fa9dd9a5b729ca0804f3fe0fe7dfeddb2e2bee9ebdab2e4706637e7f65e4e90835411a521666a8acab71deb86d33c2879377ec95e31291195942edee4ce733d80ca641b6872ccc23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1847f459903922af779d546b54beb40f8e9d556f421fa2cd19dc8fe1302cce380e89a38bd5e1ac8e58589f5a835fe3e44a485672f7470c78964b1157cdba2ee223e3fd8ece4fca55e8d0b8f66c46dc0383274dcc16578fb98686647935667356764970d10f93f9ddbb28d1fb9b0280d71e55200ab4efebf85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b446b2a36ee373cf2f83b9c2b5cd2a9e3143eace55b61947f50ada9121b20a9d7b197e6b7716cc18f61747356a9aa16212d9a3d303d260a72914e0c7e3f73363d7266fc5167c036c23ac17daffdb826ddba26cce3fe706108d5c6b7e2f7ce5618568c11081248690612e779ec35e432fc235de9b600c6f4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbe4a8592c065055d484737ce6fb711016a87db9c7f003d09244975657469efebfde08d42c9bd38ee1acd3c9b7ec45b954242dac3ae261988c88f85f8869022e7c64c2a2d8a76d70f6938f95e2ede36c910319fbaf70b92b61bed53c776ae4385e8fe704ba395c660bc935d86acaf7e0befcd03f5e1da4d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143a3345e536f752642a1ae14c3a0d99556bf6fa882be206ed42ed93096c086dc22b13043d61e9686eb530361e8d3e665f472b5c88b334c2283948fa10b2cb3dc28dfa633cb62ab680f492e7d0708b39d66be0c00ea55876e3250c084c9c33cc80e8dd5c7a1b796792d4cde9a14a21b9a343256f2419371e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e5b356cbc6a93bb030163afe0b2be797ba0bec61d4b8b1d889a3cc296920abc77d1c81927d1b95c776a9cb2eb8c5f68454869800e0cfc72c8c28859534748993c7782053052bfbebbffcf93b3f0d75acc209fdb136da580e8fcaaa0cf866dc421ba8c4b91f1bd7a048f49f426655cca30f265c792a9dacb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165263827ea4e54624d80ff5ad36361733acd4783c22c05a1f69bfb0eb97f7a55c780473ecba355d6600960372f65c17b23b931428d16a14024cb076708035c373d58442bed7085b177109c1a4222c4c7cdb9f4e81f1001264191b15c34b36846b528b772aeda236fee0be70fbad2d207fc46b2de57b02d97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1308dd599dd38817e44dbf3d3f739eb15a38e96a4286306633c32af9c09de48e8732d9df0d2198151b6f9e965554bc1fd40396a1e8f0578738610f239f06d2b852d3c85380ac896a000df8afdd7980653f390e208524e5e998a9c05fe3da491cf6408115477c9f463dbd01f3cae5b2f020dc3c4fa6ab5412a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10176632529f0c64de5d13e8905fe44fc02da58b20a86deb05edba7af356d8d68e6f30198312eb26d4681f530998f22f7183025d26d1ac85ba6dbcaa9da459017fb5b4c5ac51cf651d3d7e96217dd8b5594e22c626b12c199bc85a2148df2573222b4ac1883555c2a347d23bbf4ef42d136126bc41f29735f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1768650d27e285a4b09abc1d49bf9ed9aff76794de98b23181a2c6916288e1569a15682237f49e1f8bbd6d4b49220be4eca7e6b7f6954f387dee545d56fac1324da99556782a687059860598c38eb005e41d9e4ca73be985db5ab129282a7ed2b30a71106b3f5277171d969fbda5051fb52eaca6cd48129be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154178d5af68a03f897d26432273e5c655cb8bafe123f509c2dd7e12fbff7c46727c02917a05d559c4a83b8200d8f2ca7c13a749502b06bed028fb9ea5f9a7cfbb93ece13de94df843ff35247471af7f73ebaa370a17240aae17b8528e0a0c8e8ffbf62c57c45112d2d70ea80393a13eccc27b0e178e89fc5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h834fa2b615938a705c42b34df0f7ea32eacbfcc61a9589f6c3ce748357b3c8c962f85a7615769bf6e5a57447b124d9eaf2e62d93f6a6bfb59a56b10fd4a1c5bfb6eba0a1572ca3eef4577df4aaca6c0e23f1d05742845bcf3c2c3a516664e5e2b5c289370b77889edc01dab454285f30a8485bb01b93380f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb508840ffd1e0f29b6f6d358e04627a86a7a369af5349801efff17d4c8d4f2d627d5c8ad654afde6c71e6bbbefaf81bf136799a6d4ea6c2e3cd5ec86ac22cbd2cc33ca1a665c3185625179c113884998caec7a6aaf995ff1cc34db25d823b33c256d8288b88340d9f7d3b2cb5e004066eec48d0e3fe585a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff0ba6e99442f692f9101de937bb3462249769bccaa8ecea9ef5145c141d41e48cd15b1281586b8fe3eb9c0045e170f8073871f6be0e0b8dbb07ebd424f5b72d2ff1473f7469e46dad4d9ee5d17df8a16b343b8bb1abc5c3e4a7b07a6eb7ac6ff641f632bb35730258d07dcd31188b9b8e3c4249cc8ac727;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef80a1d3f36799eebfb5c8bdd466a621ddf38fb63fc151d67ce09fb26162c59644536afc8470980a33572e2af3ef304074202828d3d51030e466fee7f9c6d24b35c0c1176fb97fc35ed2afe744c042aa51c4175c4a4ac9e2ff0bcafeb5d5e9409a0918006f1b9d3db7955dbe543c7de5e3fad753b212585;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f542e76f136cf88d40b42aa3f1f2c8af00d981dab4f74431f485cdad54c520e8a2d1f4a94eb3116e5a109a8bebb24dbdc6044df6050c0a5d089e13358366faeec1bd375b6c137e0468f5f3acb51f97547798ba5b03a2004e94114261ed37c3de1811f538b589821ffb94b004ba493255b2e52ac367f7b68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1acf554904e198adbb7a27e8c588d7dbaec8c39d61a01f20abdb43ba5001b1ffc6a68488cd4e336049f3d9cfde8001acd5089ff80b2420b3597043177473111e0b6c5ffccb3b7dcdb709aa980780ce160643cfd7e13f4efe8bf8647c0b2a403f01da3edffb8ca712c505995ff1ef65bc251ed870fdea6b71b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd72b6e9d50d51b56f54022dcc014b50aae1fce1d4188d766f0b8ffc6c8d6e8a6aeaea8c354e8b585ced8d3a991bee958faec59a77256d1ac5bde46958a175fe64f312caf84d3f09fa4c96d71534752715af03033ba8c5cd53d2b60c4e82ac049d99cd0d6b58e2ce646ed4aa5c3e1ac2081c6efdeb1862c8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11aa8cb181417bcc91440994a0348e0145750fd6421e7c9509f482a87639c7318b7b3890c8a590d86424f90ff645da13405ee64f2919ecfb3a36bfa7f39b2f8fe8ecb7573244cb85f36dbb5029ab5dc349056bb86c95beb6c8dc6ef4d6de1e3d89de49d12fe122fe2a3cba6488dc0f5b6291dcef92a6925a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a398d067a4d38e44d8d2aec148121dd9d4b1e9ab6c4c100c0f85b97611a0117616224c28aa3582ff8ce7dcf4eb28be90d3adffbfad7dd7ab6722ca4926435654a9a5cd0fb13ef259208780b4802cf2d17bc9bb486a77710adebfe9647611cb66e4c549cd246283da25d9a7fb7cd4b167e2a1268588a88b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f3035b3b089bbdc386fbe4c98e00eba73b307f48a8050eb6f15ce349a02b60423007d020e1d6d768aaf18854da9b106e868d57ab3733e721d11b96d5e32cbe887c1a612aa63c4a856a43c040fdaf260cc893651d486183645ced5ba9f998301d4a3f4bf3616b701915793d40bdd9e17cffcec57a5648b89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a97ad98b4d2d88f1eeb97b5fb9bf650cd3ac552c13100962790a73d2f4325b892d55017f31c99f09cf1157a4e34acc9ce572adf74e451b6518dedf3c83674b3e51b6852591d411597bc1343cad4636dcbbfa7112ecd2d7b67890c5456f06d4b218d47f91c3ee6b09e70e01f0e1d1acf2fc538755c288fe0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82718cd26caeae2e88d4c5ab2192518e45dd4cac7eaabf4db991db2e77ec92b6ede2cae0b8e24826b6ac7950638e51ff24134b1f461983265fa8c93a04b602d8926f4d442115e998d98d2fb63f06726827d7a44ade7b01ac5755281a37c52077ccd32425395cc869b8e2de2218d08a7a7abcced2369185cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ad091eb2885446eed0aa81eee9fe2db37bb038a97279b796ff493703a0590d1a109843ffbeb5323101e234fc8a88952a4a5fcb1df40dd288d4a4c07fadffc522f659a684ca30ed1ce252aae93b30f8c37f2b5aa52874d6575fa2813b6025551a35d2db5df75c34e93c1af85a45a76f845241d97c8b23f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5858e26983b2d5f14d7a87267df05d5cb3d524b3b943e2de89d62af2c8ba49ce9ed59d44b3262f7dbfcdc7bff8d9edc67a3aed123afef442cce018178c1ea16fdf405298727f33b654f3c172666b5db505e958c56e2d0ce3a0b18328ad04bb72eb4a7a3fad65ab632a93e3e4d01820b8e94df88391bc2704;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc7b4f8ad69b77338010e86b5a88b4cd24892f647a8873c181fd21aee7fd8035d8ef29d493d58b2f62f9b04edeafc2675d9eb4de8e33079e2cc5e53bbcb9c4a198fa5f3d7f5b04644b6ae26acc55e422963b29d6a73b74dd0e1face3d8825c024417d93e0fbdd9339554f73ebed953ca5e1e7f7d647d611e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h494b626c8aed779d98c46ba6786c6396275b247b8948d86537047dc93c72aa917ca407da7a08fe7aaac008d4fc1bfba637c4b928268af05a0efde135055721713686faca077d16a0e7fe2c0133d098cf8c40412b4abda48bed260e6d9ee191542306dd6350165ab25cefed7c9dc4d35adf311d674ffa2e4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bc27eaa9f0f195f26cde0a6a5ab0eac6142a35de7207caa588706c72f43526ebcf4a7c4951a7e92b2a70a4b791199319a47964ffc5561c1e5fd3f5583bdfc68fc8fa32de26302780010eda65a9ccc8a724c767eb09827b467dd5e3df995eaac782351999b24f478576aa30a6e6f01451cad7ef0e4d17142;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he82893a5f0e862dbcc69485232da50e820ce9e6afbc083a1e3628e18316e2f0dc238c558e4bbdacc29a1533d139626d64e3b320ac84ecc49f7d2a1f6c50095695040d115fcfd20882916688812e86ccf630dd23789680b40c87563ec4e2713df4229566473fc65d3e7273da2d9c6900db7af2e514dbec35b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15555d6b95bd3ce915f5b7fa33a1c41c72ffa557fcc208c04cd29ba50377e5b7e0403dcc8a2de933c1400c7ec8c076271211b9f19f3513149bf81015afaf8f8d6e5c7de7def4be4c95ba54f09891ab89a81161d25b0f7e9a2170b3b1519ac80cdabebabac8ae2d6632b2602c299d829c33b6ec19c7294adb1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h305eb32498210e74d2e7b9617ddb377b3b4f4b4f02b912a67c6f315c4b0c853a1299d04610f40f77fd3dfb51bb8430a080b347619ecd83b4cc8c01af738178f39e120b9d9ffef49ce1de6418d8b34bfa83a040516444005897c6c3bc725c0fe2013b82aff2f5832fca13bb77f7e827aaa9bdad1da32a530f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfd4d735b83a7ceaa66d6ff102e1c7b5f1b3dc04ef513aa883ae97afb5628f2670fce7b0be419eeb5196c8a57c9851667c74752f5c368ba37a6781e5d131fd23b81b24497d043f3c6524e7d71bb0ea9f5697638ea01d077eb3f96d23bc209b4acb5b740cf430aea19e32c5ceec3aa47601fd425377a62308;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1848b977e177539269365e7e8b487ca2b1ef895c95f55f82cc2d599cb2cd6e725275e43a326122abe4a397ea0d3bca6d5b46932c003e35fc0962c2f0cc868c3c1a9790b7672fcca6dd90efaff45ff31d844514881813a1c092635d145f0a049c6356be765c6f59b531b54e6b898229086476f99a83a79fd7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb1edc8b5c895adaae955148c632534e039da23e4f552c2d306989075ce803e61986d3449347ec1309559749fd2414f14c4eaa8b5fa3d8d57e5c1dcbc5a99bf509aef9ded04f8fdd15abe3bfa788a599bc527649844aa204777ff9ef4b90177089cbf0417abf3919c3c152adff314bdfff61f7d4a77e66ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca4ee0730cd469c8b6c08edf256fcf2b0077f655c8ead2b9b952c454787686a5dbdd77818be048123214a2c19e0dac458c66d3275a964e5bcba93d812faeefbbfc96a3aec78a9507ea3fb0d789a372e0641b4415f499d7fbd6bbad04331e820703b7be2a93f84c09c1690ddc06e1f651ada9ceb2b2ebf95a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c7d8a297b4378740d9552697657832c78035b7345c8fdea65ae1b3596cdb7c33762e3e29ab6277c59a57c4b2449b7e3b089db4550f6041e81d82a43628c445a14d339b44a3fe6577917da6e27a9aaf9cbb23c7cbcaeb41b403e120569ea029e7eeaa8efbaa94493ecc5e77228d2c4362cca06c03d52aa54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc509e7dfd17e3e70815497be979b1fa8312b2248f63aee1851e8a88809eaf7c884d211a20263d8478172e0d1b4c5c0025f8337f1e027a8e2a29fa3afa3846a655811551793debf5bfc84925bb31fb627922ecc75b4d03c3fa8d814481801acf8dbf7a5f53c8a8a070c9c9ab4eda4f011417fdd32b1472556;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15882ca775d4c6c4484afdedad2af0128c00eb54e157ed146e84f776c3d5f698b72f39d322398902f2fd489a6be3b1913636b5de5003bc6a71d9bb27b8e3b0403dfe3b3dc0f42694b806c5de43d613dc83ef5c644d33684ef6fa0f70f3de0589b7f99a612b3041b005ecbeece3a5248613be0836d47e30c73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d6c50bb06df8abb3968c2e2e477fb4ecdbab70be06665a6f55c50dae9423df169d469a882bd1bd155ce19bf1be9113436782d08ed87fd415dea27eb8a1fa05e02c17aacecf0ea3b6895e0c7e9de29ab1c7fea6695aec9c42969c8aa637724d19ee816c00294fb51cac919458f8fe990568c1e89f0d9c4d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2908d8783303697a49a78da72002ee9a4d31eeac0e9102b88a833bbd54b78afacf19d5d0992c20a4331f97de87b3aff1062d2d7221dfbb9becc9e56729b54daa78c92eff439c7aa9099b5e3b19197abc5abda6c4621218bd724b3cf5a30112722931ef4f88d1e76c6f77dcdc87de166516d6f8f3af5592fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197595714e6c14fde3428652fe52574870edea2fc589462f623cdddf21c14a202b23554cb49d860e2dff0b0683747b12f560d61cfa4128ec57f02f1ffb96ccd7b1176bfc43111f7c1ba99e4b3f537811929fa4576bae862ed8286c6bcddf77130fb6da47021e2ec479276436e04d32ef6a1854a41745141d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b41595211c4ba44122b96302b0b0eb5e2cab21416b627c77fb87bc13edbeafe6989d32f77cad12fa3d0443ba058e537316550d0907837ad64a5f742350ace3dc91dcae3361676459efd4d4859f56284c18dc56945a3511ee88696e6551511a2a8eb7d0f4e53b4c21ac668065bf827cce7638ab65cbf0a281;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b99ef2fefecb98de3a08b27be3768bfc9aa1340606844de7f250d590302976664a1a4e2fc111e3d2b1245dae1d45a502f327f27286c949c61d6f293a6b2a3f15cd75d202e57c9b25291e6a8e919ca693bee87a32cebdfaa7b129fd80a3629586775e7a768743c72dd18bc4add51ec447510f751604297d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0b085a5f750ffff13c1f032017010e70b2c7e69326bf666f0a0222d611e9ea98826995210a1df3b0961418ccde8e71e81b6efc6361baf929a9da73abe629ea5a7624e15fdf2dc09d7ffd7bdf84f84b2c677a61c17b79ae74b6b2e228cc1bf7de7d9dbc2d9037d561f208804b787e062f1dbf6cfdef46bc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94d2af1704a5f1bf86997abfe1831adca6f4a88f9f1497a4b8aab68368f6cd31f4463919841bc8ef5b7fe65e9710f8e5732cffe39e8aaf016361ccb39440ed4fb9a2f3cad1c267486ef30408a56e4b7b4a19649b9c8b3eaca5717959a642520f4fe46dfafb855eaadad97d3c094d00dfd37cf40dbcc38fd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbba6aeb7de99a574658ba6a5fc5b0b2841cff23baf212e60a3e66eacb8b3074deb1a8c9cdab18aae31ea87d0b7efff5b0aceb391c4556aa743de3295c2dcdcf6e40bc9175b909b456b83c394982aacd8d17f10ac0a46d23c18d22333bffc9efb5e488ab0eb628f838f0944acf6a81f6d7ed632abe897441;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ad0818f4ec494273dd0f32ac3af51d788ace55437bc27e6c283ee852ccff0f600dabf06e1a025c7d83bafa8bbfe9dc284de0216961912c6d2782702bd83425ecbe799d2a26fdcf2784c45b9ef9e8fea4b72c2ffa3a14fc310836427fdd22ca2f8874a5d077f21a05f9d3949ee509ea90b65d23842c48db9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13cf0150660208ea4a2f13e15612e0defe6acae6ff4f6b1cb7a8c80c1124d53a99b6c8b892385d3412eac4c9f9bcde934a51fc0b468129649f7322e67fcb8ab4c183d7cb3795f9a2b98e384c4dadf687730b0cf1b2e5d9a93ab8f560e6d3775c24f4cb814be29441fb68f416dab0532a39a6ab2a5c2a8a2f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4d2243b288bf77e2ad0002fca6ee8aa6d5b2f21da4dc98814afccd750e30d676ef9183de758fa55d0c416e0a62718d6b7e75fc6416d5682aa25583996c3d58290d7c3d8af66e342e1d22282d61c2be296737d4fbbce525cf32e050b145bf568bacb929d4f5c3bd64a9a2abf7192b179408f78c30bdd4032;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e0d1d579fb5f7077901ca1a56fe6db0cd2fc5a88e82cd2d8bab904d03d19bbfd13119a535f96b5be17033cab409c7c23808395a069caf2611508e575495d058dc90be128058de75a98421b6937dd24bc7f6367bb5a7b8be3ff2077c4d7421678707bd2a6af15b82f8a33e200d596698a551790d4d6f0f0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c04e51f06a13ccf64b5002bbe7ba9061c75d8023b7af1b88f856a5f53542779c894a9d95bb144d32c6ef9e6cbafdd287adfb18bc4aee7d8b73c9efd4f770689ffd1a3c62e1551a0542a037ce4997d0812db25be8cc83fcbd9e39d5cfb37b3b2b7d78c757ccbaff6c05ce60c55b0e9046d4b553e6c63c886a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a019b767bdaaa02c7189265815fb8b21c889335bfd11d2b15bbb94c105dfe18c2b44448dd42b3a40ac094d5d05d67647b467129ad115e14bc5479d5101ded932f7392f59aaba01fdcb7e7fbe2e122b751ea1c567b0fddc3ca20adaa39882b52b1e290394c880ce6205647e82c6e325bec5409a4273c145a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35bc7caf8342907231db32a928254ea25d4f5e19a4b0c6376d00c8c08e5f4be5bc9874a5e85bd3e1efdd36e12f72e22378d601c139cb89ab6c800f5577203f5d3b3fb49ac0899fc0620ccbf511f3602e17fa25f6400322c1246ec52db60a706238ac84647253d861b6afc9a78fcf066c2156e5928e030bde;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c73d236cb62157f0e98cfb32c913f6b133f1976575b8d4142d057f00607ea8fcac6b8a6a3d1b997c19c208703f926c1297f7b50c30940af5f9809c68e4ef0f271cfe3f394a9edfabec742ec0e23dd925aa11c0974cbaf70630ddc6df66a843abb1b282cea8353579d0cf3dc29f2585d62a074e6c161013;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a15a94b813aa1532c5b21b4d723a669cf39603be7da551cd68a54c4236c1bf21437c8167f17fdfa4968354c34aec26213386073b51b686ea0d9eca98076910b5f84fe575015ca57063fe405aa3e02155ce0d2d18b6b567aa394090e9fccbb669627dbde700c31b6470cd77bcb9d636fa657541f2da3db18a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h826e82c88d7db57375e5f949a7de18d75f7f4fccc482fbd035e7d08b5ca1ef0ad2e35ea27fef3363dac8073bc5084261d2314c1be71eb5e131f619f4f59bc9d12bac6137681267d6dd7495125258b490e263f6bd60fd2c7c3244f68d79f102f72e30e0bd68057d9478950f7048872de26764dff18d2c7f68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18819f004a44eaed2be312efbbfb763510639b9f3810a87df6d2025cede982315c9bb5cde4eca3d1608cc2dfc6c4772cc9f55650ef7db876d394ac08eac67b40fb218c7565f2302e90ceae0d9b1ff365295a90b3dd4bde47e1718fa48b7346c560673b59cc8e6b431e222512505884f745ab6f74ebac71231;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132573e039fe81f3b0478fc2e1d8e522f09a92baf5f73635d2f3fb9f311ab7d6fd091429b0713f01f0094e8f2791f328bf4f426df2a737f0aa926e04339fbcc467233525035e1d1ef4f96f4ce78543e820d3f902f389c7035d82aaf9276f7f226a7c6651761f3ec24d87f1a6061bc16db5a22fe7153cc38d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9e36ce149984a82ccd9646ce32e503cf11d88a6991bd472b5ca99be55a800a6804d21bbdb5914cd172d5299a73ec07f6e2fc88cb1aa29719844c7cbbb1fbfb2ea2184c8949065f1598cd34af85bb17e9e2cc896a5e2542791fc0adaf0621e2cde7f7b366b5bdcd304a1ef7f1ac1cb852153810dcdf30ce0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h554c607f9de9a8b328549f15e9b7633bed6cf9a95d01a786a089ef6934c7a21f5248b549bf7c31ce8788d32949a4673fd0866ea321e8d2d608c444a7157af3f945b9aab5377b4adec14172adf1b315ba71d05e93c526bd18819d921483015badaed5342ac4424fe59fbf403b4e8f1a87abdf253dcd2b15a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2991a49824b55193582fd59f3f29bddbaf72d22b1eed26e256feea2c12faf719e24ab9bc53ec1659774f86f68cb809fc7f2f7b4e8bec17cf285188a0a4d8b67137f434094d8cc3bebcd6e721291a2c0181543dea4c185809237e2cf687337de0c5b93fd0e81321dc2e807cc6edff6038c7a98d33f0be5723;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1757a70e2abca9ecf1ce5b65d01abb74a10abd7c8f4c33b48d3927e62d93889ab0978cb914512916c4666f82d915d44f8f4fdcbafba17f83ee79fec6237884c306abfd03271acb42524a33de27f8c08067c49d8d78adbad5b3b3122d6c79e4ac5d33698a2eb4c2356d6ee9ae718c4d59bb16fe288f84633d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf342b52029e68cadca0aa44830b1940db9cd09b80671b2f9be7a54d5607022876d6121808ca411c9fe5dda89c6d33fd3706cd0ec7d7fefde39c4de97e49ac5090b72b23b9ee6ce599cd6a8fe2a0e9ef33015d1e5d173063469d9243853b0f138df09a09f089ad6c8f528dc89f62c849994cac19e9de82114;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bdc08fcd1b12a57a877fecd376d91cb6137569ad0d0e64f354dcefcb26d7ea3aa4356a0d78e6d580ec209d452a9748dbd786c5ad5ddfa29d70a110e230e5324e86c1059c07067fce0c6b3381385611fea466a4da7396758700a2e820322e2279cad2a9993ab85e03fca5d3d024997483ee136600684f0b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfc3a18eeea04c3542863e93f212e3ba86f536589166148aedd51b821c6b7595b4faf47207ca0a1798a322265f0904fdfa238d481e6e545a834cc331d3faf27500476aa266ac41a30c5d09f66d85de1da9e947dadc4e178ebd4744fa2cf1be7f18f06f1490a893646569ad67c55b3c795c260a999ebe2fd1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185583597253c184bc1549172e3dee3884e5758cf9f22bc6d1d90967c7b187af7a756626beb68acd91d04583a2eba6c529246495d49945dd3bde740912dfa28ba8ef9544fc741682a2caf6805f5115e017c84e618ef01eaea82e29f892ff878ee61ea6730687ffd8cc3fc2dcc35b99541063b8a9cbe93ba58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50b695175182953944704496b836df90ac22095d087dc2a0382dcf52a375391aa15242f37cc41a2b9f6dae8a9984efd092d69c3eff28dccdad331167df916a96ca39115e4dca2643d5044538a14bc7020ceeb12d2f904f7599818500a90d62a1fbccb0d94035040642d6a2ecb61f31641cdec84a47c06eb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1bbddc709ff5de3ad3110cadc48ab2ce2a32a5f8f8d2410dc8b26fb40c253e1957ed555187f50f5ff510669500190f1bed35a6b767edc414bfc2211917de60840cb012eb7955dd46a5540c177f566b8dd3f961463e6af91b0f750f5080a5d75b5b4d7df082d12bce85cb9920caf5ea2a611923d2d73b185;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5004b3df9c9f786401a5d837402ed6d27fc8c76095bbe1fe221393f799869d85ed2e3ce07ee0ed4cc6a29c56d451d8e7f756e699c33b43bb5eea8b8f62e96ad6bcbb37987c08e1f0e324aadbb138a7babc6b34208bd3a8aa18721402f3e105d0a46ab471a6cac8ec648bbd7c42c96a730015a9aa404361c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38e190864abb90c4566c49175b99b846ced8dd446f0476ab33a5c33736377dfcc1c36ff9e3cf9fb783af25f246e5e2a48deb7e2dccd291f0427070258e24f73663f86a03d4568d612880636cc3e0a83628eab78a39f1f74bc8dc912d7dc4a7d6acd4248fe2db1736c02ea91e14e7c0b720f2d03c6c965745;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9853297e660d8419c1c591fcddc91a25e909ae5cf0f3ef0acfd22965acf7aee39a46ce2b94f75c8be8574ddd38bc76de9ba98e5ef48ab732df160f0bfca077b2ce338a5961edbdff4bd692942960eb41b5c2c6356ddca1c2647501606befbb02ec738b0ccc80b1aba698f6da9857e2d192b4d28ced83e2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2d8de560e80f2a17b269cb05baf89b8bc80ebf5ab6568200d25a242d678bab94d9e694249723fefa4f0b3184d9bfdb554ee4503edc5cc796189c58a80fdd8d3c9e772d33bdae2f91cb9d7044c13aab256b24f69ce15e00ad58eddd4ad1b62c23d566a81ba1c540f51cd9d0c500530e9f7598813b9fe6804;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha130e8634a1810b6896eaed7a33e8687df679c7196ff6c16423409b1219ae36fa6e7db4245ff1b1e6847edfaaa37c907b890eddcb013a6528b8d286dcc5de480f030b0b25183c132a202509528c6a0c02391c830002bc8f12be337fbae9244eadc81142ee7acb5394ff8b5d9089ee0f0fd5f9c1d31b0168b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2cb06eb6e57eb118bb54f14aa319bde3381c13867878ab4212acfc66079becb361ab12b87ae57f783bd22b642b11e1709637fcbb8d4fc86093b4e970081f5b39662eba55cc5c6260fb2ee0f4487a676471f23ea2de1cbdc771d2235df59e208436970f0e24a8ed6c67a46cef33601158998e3b7d234ac3e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h800354b575295c3cd3a1f879876f32ec746837c97231f7e1ba6456db65daa99bff77ff14baaca35d784849cc06f0704c8a1530087d15de97f847b5573a0a1c5610d8bf59d8b5636f9c17ef727196d663411c9f927c61bd3d3d6c7793f2bb2fc8a27b2fedaed9cf38218ac7a711b144a1eda05e5bf3646a49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14507c0c2858b86c2f858dc66ba2648c16688d485e069aff65e486082b88df32f475cf2a1c4bcc1d66ba6c78834e9adb85bbce322f57147d8b8d88541e460f250039f4ffe52ec1fa1b27890396dd86d7cdea33ce9bcb8a959b228baeb825d2dd80987eca4754bcfc2f104403d6c15ebb641576fbd76674a77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12671b356ff240a0cca0b8397ae151a5d20dca9fe92481e69eb350a22547ccb528c93ab546acbbaf1ff8eefe04b28fc5dba37d08987ad3a2e9a78836bddedeab397888f2123724a81867d3af65144d05f0925f324cfad4a5ed3974199b06b4c64e1312abc5c1c7edcfc8ce8ec00372b8b7efcb07b0af306e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c218b0242366bdb96c1a267ac38315bffd21a4929bc1c18d4c84b13f20cc71308e40fb577879b4effeb8cd365001b14945389b1e72aabee60dfcf857d9cfc4aa9e2202b2641d650b86290dea58b4753e2fa6efe49bfe0900a50655ec38314c07f462391620a6b37aec18a3b0a0404b61c0b879ec661bfe43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b30aa9005bab939730e0a6693444b403d7ade30f2ddc5ef8c6be6695a050ac27337e5bacea1e5e4b64ea51a736a85d33d38b84f9105c44eb545dfc3a8b4a69fcf4ac7e9fc4e9f5359a43c8ffa2294f318b343a14c559bb25dc87a1d804d7a22c811558dc89d10a8591c8a208a86891e3816aa721d7ca2c8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6fa68de4d52cb237b660a84b0f9fb6f0c0ff0d18d4fcf1e7cd15cfabdb048c64661b2f6fe51aa1f461675b19be15ec2c2d051cc752874f3c7179d50331bce9e1959fad1f939f8db66c81163ab23c39faa34940169fc323cfde58ccd79bea46df4f5e0536958ff09ddad1600051526e4c5115777c903d863;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2dff3cf1761cf7e5c77f70e61254d8c67987ff91ba86491927cfd7bc4dea1ab1dc317e527a99a922b166759865cfa9be88c3cd2c94ada486c27fa138bb51cd52298633eaa7ffe9e09aefb392b40c7f94df7a00f85f0059f760c4d441d956c549764654d5fe8b12050cbf40180dd59881756d39dde3c2e36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b095b0948c72a9c3008b9f758997fceb75b37fe91f99a2e509983300df06312be3a35fd08b9753a225178bd6e942b977eaf7714316d0db2f7253cc9ad88fc4d17e0bd50e214e50cde3ff451f8a1456059f6ce88cbb4e4d6461ac285ab5c93e64e4271cd9668a5a0bead67e1da8186994bf9b4e68a38babd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f466e0bc04c13fec6eec278d06742df70904fa90f2d675ef04c33412ca9da0a67ec7cd69a2278e9d30f9927d0cb9acaa472e01ce41e5d8c323d3f3cb4ef804802431f6ed62f25564f1030d15ca786fc654fb818787a7d7ed96e5422dff8e881a08301af475f17651cb9c5a1e85ee2d51dd715d1280cf5ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34ad7a494bb3f0294b85556eb474a1287724f9b928413fb012e6210c4d7d55df1a55a6fadd9eab2040421ff73f7127c51584eb27cfe9a763c0477e3144b03c0fbf38f46f4c0fdb1a2f11751f365ae6c6db4b9a6d1fa2f35ba4541ed304b30cba985bb60cbae03a0a6123ceddf470bb53ba07d4d8304855b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f3c01608d52c0a77356a74a87faf028b57502229e30543d2f8cc28d4e6ca3c61e4f9798ec50a611fceacda67da6c1ed32aa8b4800eb4b1e3b9686f00128a7ca26d39bab3e110ccadaa2d0f273e75447e73f29f6bea123ff5f8ef13dfc63ee4af4593f8dc232782e5b8f6a75d1930d92426f64f5cb5445c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105c10cef2096396f6f4d7df70b4cd87adf55c94bfe112e7f94e4c7c4e49ead1a178b16c3771335b90b04f6f43c693abc709679739581f8e841c995cb4eb9742adeb9f0c469417887f89657ab014d83acf1b77398bd97a29a52545019e68603b34615fb8d06a43b8ecbfc3df29a4fb18ffe13db2a90ba27ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h528085ffa57e71300ad165c81292ab42d2f8336e920fbff5db7d6d7e49803867542c7d905f5816906e847b8f193c4225e8098ebe1a4b7ffbe873bb98c245083c7e7e697dffa1880b02b605025fa69c6aa5f1b9a8b0ae921597f0379f230ffa4c134f21798e387be8233816ccc31ed4d681a92321735b75ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h977d43179218a608e5c4fe79c9b8c054bda86b1b4133c7d3dd0ac6b5260f0f7256ab2cb2dd3fcbc9703d9278bf8ed8771c83de32f549df7a332dd33a3466974b7871eb7e0e0687f01f929e3812805eb9d341b420793e264edf4c2eb25dbe1497a4c4cdd2579bf8e9373660fe2a8468cfb9504c1dde7faae6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e84896152e4b512bf5f54215fb1d9a6e1df710b0eab57ab200973c01b5600f81b34d51995689f293a4be6d229f6942fc36c67066bb9065d3cbb67acd128656b5d9a3b25ea951787f76184ce85b7789d35bc467a8e528c4e205b4f8191814d40f4c91725de2547b1584b6166da16e5eb55b2a49c676283db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae28be3e6af6bc2c9335c29b03527f8544fdb4b35700459e31d0f41cd4949493ee6e6d0fb126e9e54f39428ce82a39f3b4098c33069f4d2c2f570e2064029c4652cb2199dadfddbea068e3a4f1a83eef11ed0c61271759bd3cebdd35f2d97e9b3b6eeca7a29663100affd1eb2c2a37fe80f83e110a99c594;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150c8fedbced1c1928b95515fea420ffa1a7fae8490694d1d5fdd098787a79f836975fa39c34e90a1ae1b7e3e9cc18c55a2d976ee89b6bfa9e5108e40b3486c4477db8eafad541cb89723ba17dc50e3ccb683dabd602990bc202b65065a96cce1f89d14fc0aa506e9aadd837f22f64cd627ab2f7d12a2533a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c0fe74a37be94865f6cfe48bc3254a2f8e7386225530f0c90a3de44c8573e396f018eda5d116730a7bf7f84f3c8dbb7c12d1bcbb265dc2ad5dcdca72b786158222b80e3b83d3004d6ffa8ff53ad59d4a319db0c605e139a93de2e4188db6fcaf982cde682e95bb69259a2b76aa19ce37d976c53f2b7a215;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b8b3014a0bf1d75247f2421e7ddb4a08dbb5235c55b8fcd929c55db17869a31069503b1cc7c61d44fbf3dc60bab4006ce38a441b39a470484bbf427b4ede9c1f1d4eb3cdd26d5d48b8dea5fa0df02b3cb5540407d1fc27edb85fc04daa1df19b9c76cfa19c81d26dd70bbcd9a503b5759cdee1baa94770e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h549abfc6b834ee72d0064d848b3daeff0ba56a5290d9f933ec3b9b99a4fb91f9867dc6a71ec21a0db9be56f8ebf8de8bcca0a7720bbb110febf912c2ae209d5dc3e2383103aa6c6ebef7ee6a78eee0aac3d6129d5a986cc97b73511351da06002d76c54b5b5de4acf3f43206b349804e90a1b8b385d3f9d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c9cb2943b0d30f687af34c4ddedd9a817c37cb68bf016fa748adfbf440a50f074fa0396fdbebae8e74e605c0536dbbb63d3fb3cbd7cf874d27a4bcb9a78baabd0b1b20e6a1dda641998a08b89974c8d9b755b2b0093bc2bff78a3ea2228d4b0f9e8a8a302284b1fcfdcf1d684240e492218e7f80fa5910;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cab24ca9b7f9cd7a6c180982d31639780515d30b61e3b2890bfb68684c2d1c65fdc9e7320eac5681ea524c221195bed0cfd2e45ad8e575f2f99eb4a07ca8e43c4930b3338076e087aa83f448e73479ae56330fbfcbc34ab6e7b47b44aee060af117ba470b9f755b87dc4d03506407a2db68afaac4846e2d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4749f6a69b2382d99f7f6aeabab91ebd1215992623af648b585e96c5fc363f23498cd3a4dd8dc66a479a25e965be9a6e5ff427a78f35a0efaa09a8b772fd0d0d548835f8829b3a98cd496f81dabd7cc31d77ca2907daa0ec630e07f8391d697543fefd496d7b4579ffecf856766b74e4b1755139a3420706;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haaa1fc74735f31b0752954336192ed7baad03da46111b27bd52f026938b49aecef9205fe477a5bda4efa6a1640206a6fbad1cf24ffe866a8874943b61c8bb1a29095ff495362c88e2567aba2ed905e1b71e28f6df37ec4260be5ff94566a69d839d8131ba1ee2371e872bdae4173617afc7048337d826756;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a08df0360e78a9d27419aadf2334dd422eba16a256ff106164a0a414911fc4a59256a99db48aeb4da147c0a7e45d9c1dc87f1a258831383593b5895004c887234955b00aa2e0dab7e16f766ef8ab914b43998c8fc9ecd6d4cbae3975a013c9154c0e4df246e9d9b54174a7f99c5499ea29e9efb08efa545;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d71a871bc84384105986d5684fa2969a79af76b6fc1745dabf939078298d2f5f91334b3fde14be42f925c6a3312249520b99591a6d16b49dc210186782632298fe6ccae2b4276621995e36cc494595143514ffa35bb789add7479f27e8b08a45af569a73f39f08a43ad81c2b8e6fbaa8a382de327b11c5f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1b523e47459f876e736af6b65c11132c12b66d6f00c9814b5f2610479df641a1a19883e38535b8f804da6217796127fe4db6bc5370a93f2003a33769fcc014a0bebe6266af9aeb585cfb9d2f1c8b564729e8e4f19052ca0ffa34d4c20f36b150cad14634a25564c72c92c434826b2ab13d1b4948fca2f76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175687d020319342aac46592e2940b80d59a11b4b601187bbec1dbee7b51b71c456844b9080119fa8258ee5c7a7a55d52b746b3e020b2936adeb275dffea6ff2e257505af3c303a5ee2f9015cd6c5e7f5e3e7004ef33f9f7e64a5ef697a9947d3b1d8e5c9de3af858ffe9045517f293f08db474d7915f5f3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139413927498bffe85b9385fc32d7409801e8a2fbf9e3b4f63b27f5db17accb954aca8946881841cfbbf8229fbbe97de0177efb5edae2aa44b700651d534f54426888ddfe8cd1a3d6fc78a312ee47e955f6eb85833f3ed09bb98751112559ee593843f5fd2c1c32716630f2bd850d15b480629f71532e3574;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163334d120c76a8994f578fdd3653ddbc4e8590d997d1c7401d5312ef0691ca468dc784e844b6cd76cf4457a7d3655f8d8ba79c7a335232e15ab6f0003e57fb7772fe38cd5031a79edd9185cf49ad4332c88050ea7ae5aaeeda9dde3d45bd43ab4ebec0b7c8593ac2336343f16cf345a1a405e5a5e74f63cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8aa0109aba5ddb82002052e95733d979ddff094b11ea222db99e7f03afbd4cccbc59f512c630ac800aaca9125fd59059a917e0035e8e372ceb18a390972c50f4202e541098e304d5bac433af0bb61db7626be67cafc70d66814b8e0f2e125ee5d01ccd881f249844b2659dae027c628f6c6becf63c5ec97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd192b9b96b19516bb7898ded2eae1f07942257616795d32e5b40afc7b505e0117943e40d04110ae47aecbc7194599ccf2c2654d9fefb843f401fa1c719a98a754d8957d7a672b26574187f53b7757412da521cf1685f0aebff587e69c6672b49e36aff05a4f5461a28476bb4797771041c22439d19983ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0ef906c44c63416b50b875950af7b4e34c8994c55eeb4d7a03ff5c04184e4c0f065660a137f9b6d428247241a0c20242c40559797d9e308dfe18f6888d23ea262a301d28bedce99a374b1919357773a88c81b57c672dca77c6b1ae4493df27d496b1547fdb175c8b0b6904794270059952444be9b179443;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d84383328dc4d32ded96d05c28d3515a5ff19baf0ecc0715e95b129d49b858e4f359daac15876892cd1fd675d37bdf37806689e92882d61c88964cd0084db0a3fad3b6fa66132ca03ea3a1f956e14cd773d2a394067df9f64dd09dace14f183754a576dccaa4709e7e70045fa2f5a76b73d820415cdbb256;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2dfff1de0b9e91143ad0791f51d76fc2af74c60e4d891ba043f856997bf5bbb4b1cb9b8a1b8555ef22154e23a6761c20a1212d903acfa441dc41a0c5119adbc625268bd8403cef4b023f618812a577a15405ee43e415819a3989a26bb8329fa23f8722529970ece29abf5df01c039c57c9f1c5d3f6e7dcb6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h981c7f560fccfcf0e962b1a4d94da322de5edacf91825078489ffbacd68b9fa1268263e0ca47b09947853c59d4c8830a6649d69e13b8139be5a62cfe66b5d62b1c6b61ad9a1f59b776acbf9f671129b9b4e761c7a90de772a0448cda117af6af4c91e2d0a576190c79df273040c8da24c5c605d718404a1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128acc935dbaccadd06fbcaae72d486788da98046ccda58b0db1cea9a134e3344ecff7810ec737248d09435993a477b4b478ebe4a73a89d07599c4ae46429df419b10f3137a603b4151dff18cb18a30c2de6e910f8c7a4b2dfdd52065214b56ea144a789511a0c564ba5970e857cd9960c1d1042ca7579e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbea4009d0880730838995f0969d515580fcc372649dd6e031ef5abf1855b95ef8bf8885cb185e1c6a378ef97ff57bac7e19298b5aea96a3170eb0464a6447352876aa02feeb998b21ff95b750295f77ad27227273c8705c9a3fb48dca1eead39a65062ab67b9dfc78e6f66e596120427af9948280649e31c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbcb65ba871f25413977c11897c5264cc749623c1f335f0567dd1ff054a6f383f7dcacb8190fc158ca429a26eaa4ae9aa4182d6e1613ede9faf0a26e9ebce4f6c20ed225f997e0ce6811d4f42ccb122f1f044b3e9f9ed7f27de63ad8406dcccfa5742a0894c13d17946c94e6282e095ef6b7a5b7340bacc6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a92072d7618159ba244a712c19911658e68a71e968c50ee888f060c73dec34ca297a0d543f46ac271110dceaa8e84b5dd2a7cce9a7209e9a68990f48eda428138324e974795f10baf01f8141a304f47c3c9bf41411c965b5f7d730053245ab59adf2add2e7b7b262cfc9a8b9e1d0187a65d60d4d4f0d7196;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60696b215489b67c89c0a268640ee5e428bf9d3d1b661f3cd834698826ee45a289e00cc770d6ef3f9bcf64e13b7c4d3e41c945c5514d6b244f9127cf6bf639a82eb469be528978259874abc485d512b5e7e5c17dc3a911efa3b5083c790f38991083d20f8c23dba2b748d71b42a8f0c0c7fdd89875dda4c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1103f8490a43a0549d8a27862aff965acaabe1ff74289b1fe22dd81bfc6b480858a894e7638c9c4ece32944b626ae79c0bbe44647957546bf01f4657b6335367f6b4da0c721be066e432bcc1344b9a47d860ca4941c723f204e7c05727410e966f26adf5c7b45a651c738e30e4ea7d7d5ccb2e4dfd8af3fbc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10427bf30252457cd56670f42f2ece93f07089198393639175b50665d8516f10e8ab0ad03eb3325d14ced7bd0de270cc350884ccf52f00201f991e33d3f931c0ce68c6fd6595f77ac87758f9ba4ba25a30075f839ef4739691f0412ca393d45fdcb1397e75fc5ec76fde5eb03bb26f0ec3108d29beff7ec83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19543615b67401ecf42939696bc91357d7812fad35cc36fd37fa122bd014bb26b142ad9b8ef676236e85db621f1091146998a3cfbb5d4a01de3f4aec4e55dcc70a0bc95979685f891cca83e66a8060066014d9abbb230d1c57b32cb168421541710eba8b2498fe5f1fd31c52d7c5cbb39a88c0aa1edfd0e07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54b9340e2145a486c50392912a5a023459203f89691beb48cd5797c2fcecdf94f88b5116c0987ae4a9ad136a34be4f8d46682a5f4e02b390f2b6c984c01c9789f5c346062700e6f7502b077161f8946cf1e25cd3426a0d2c40ff82b251289b90dec73001a90f0fb02feaabfaf623ff4063fe9f56b313716f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b226e84721f91d2a6122f685bf2d242d71b902ac49c4d7b68c8a7de2d0cd73fa3c18fbc0d4337f26b949927c678c40c9aea9cebf16e884d74c4b5202ee1aa5392edfcc887fe6330066fc8dcddf60d4d8a94b401c5330b3d4a6b1fd977db714cb0faebd8f5126e2243334ed996b5d4799ce6f5d9e41912559;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15edd907699d2268e3fb525abd6d6d75560168ceb5b1336318735fb25f6995286638b2bacfc2ea883086bb1f753f9e3b87037dc9bf6ba3d5aa21183b72a76aceb6c1a8dcc8092a6aa3d44fbb52567ab8a1dfd8fad35c7468896bdfce51dc3e4424b3a20bba81e178e72ac89e787d2bd2aac2aee007e73ddcc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ef19f4cfbc327936936f641fb45329ff05b43ab46e2a5acdd17893731a3320904742d8cf189134aa153ecc013fd4da4704b0ec9bc2221b261a946a25f8ce86e0eaf2e5559c1b03d20d2da2b7d013e7af69143d2098d8dac865a9047223a8eab8c07d538098050669113145f22b3522aaf5bc2fdcc2927bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c3790f4fe275f87533d11067f00de9c9209246a3c5058f37ed7708e79fc0b945dfc8651f0ef16afaeb4e8b5855473e897ee31357f77fbd5d1c11511d97c4fb6a1e0f84f8b28aeb4c15e3d269deeed3c11ad8db2ef992f5ee06f136cf03082141d827db2d708e2c694b97b486a4ca56352bdec0b7158616e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6e5697a39315617ab93b4740018c7342bd0e0554282d4199869455af4d9380214e5d8b8e554881e4b53a2f0d1691ba87edf3784832a8aa1e57ef4c7cf1d96ab7af6204860f3dd68129c9cb0e4f8462630bdc2adc4c0981d1ce90ef7996002bf23d3c57f5e8d3f92dc6bbc865b55a233bf5bcf255ad3556e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3fd2609d3000cd65c9f371a5c0b2ebf96a8e5030503e37dec0918523fa901e545fa2b6b60ef2860b9233e814ead14f91ab16b6909ed2daca1718286889522037b09efd5e33c04e5f8293fda344513afe758f23379ce911d7118d1f0e680b8884f697721495935d1540a318ebf7cc7e55fdbd551a14705e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h960bb94f8176125f42e57fe7b15b7acdaa6ec3a01a707c708d29e8293c49fd0a19d995a1003ecaf31e017405c0ce638d16a9969ef9945d3ad5440edde674aee52a3b620fb34de0619d5e0dc508bc3a514cedd202345e1d7e854931d96f8b8a0250725ea83917afd7b15b484eadc29ae08e06b64882487081;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47285da432f481de1a44b9fafb9bb9db602beafbc92d9c4dda23fd157998bdf3f101ccff4f48bb46d335c1b2904dfb9a9e224550cc7207b34b68a5d938512bd2f0c36ef325d55a65853c610f4d60b3180055ae6dce1cea77c1fd474b36a91a72540fb99dffcb3294e1e6623eb882ba6937d554859d057120;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f17fe329e4aea5d11b8c67a6ec28944fda3980e137f31d9aed070584688c60ded2db997463cb7bec91338112a8e2d5aad476858dddd62bc49c895395ee1f1f0e6b1674e551cfd719c3e19bee7a74a607472f32699de022fd9404d5a696cad49f19a8b6ff1f5d893a7e3fae1bf16189e8928d55dc477977c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9333ecffa85c1144615f580a62ef89a3e012a557242843bf33517faf19d6f3380241df1a8517c6005f160b85514ba4b31b3680a50b23ac47dfde8d5b9b112424737faf7e24eaa1a521c1d7c3eb788afa90673c9f0a9d656988ad307084297aea9cc86ede9a7929b73ee7d8f59448f449f974c8354454c2d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d6f150fc967bb59b48fc730e5dd0d40cd0ee4fe108d37e04db7185403115477d0e9eb1059f91f1f510c473442e9cacaa47c3936a608f1f0d79c2ed556520d44c3c43728af3b8fc88032de07ac72fc80913120cd136fe74aa80c112e8de1af7ccc0e34fdc78e02aa24007ebfa6e069c639fdd8e05717ec7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3de4808f2568e505b185593fb67351a3b985330002ae097928671a44b58a3647a75db21959526ca97ea0e7670c7822b6581491581e01183fea2f7a03ad920906cc4cb3c2fbbc2bd88cb2a1697ceb5cbda572e27f006cdd1ec7f66c54f4650adbfd92743b089c3db5a81b736c14d722667805698087272271;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cbbe7c0e2a0135bb054529e1ad823fa02a9cd74cd656aadb88a4731aca306b5a9cffac18b3bf1c810356c76059b0ce758d7b69c09361485963116a1f369bc39c429a288a9f2f55426f08f7f8692476afef4399019287481dce0f0e03f6efb25919dccba7d26e3465e87c3e4418a0848769c4a67414d147;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4f942ded612b56a4f1484cd2cab98b1f58f9fb1b4c5c5418d5e6d478901029046f6a508194e4d706b58deeb55471049842167826f8337c765a62b6bba1dd3d8888754294115cb6aad570993a777c200a0c3d7f4b8f275d261be17bc8202d625ed9c4e11f6e39be12c139dfd3310f41f2d0647911e76a6de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca4898d16c013ece09168f8793844be6c987cbbd100fd7ee3fc70cf74784318bcf86b60378201515722d161cfeb1790e4295e79653cd8ddfa6d34521d83748313b01d5f73ca5bf9d060c13c9a865ea08177b5c511814c7df33e91d2b8ecf0014894845fbc34f78d2f09a040f4b143c95134958d69aa1a362;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h670e9a764ea7b80f33d312bd2ea9b44625d4aa9739fed005d464e93c932a27f320ac09dcba033c50bb7f942a77055565db411f9f31e7d69e11a68d049ff0932608b049d23b90cd9a5bfc99e0f44d69f633c307b10cfa20ceefbbd89679ab3be2308c8fef49ba3bd86d0ef6157af5f025a65f78a65a4a6774;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc0c4b19b6b981890f4558ec8628b58830bcd18be3edfe9dfa41a8639da2d0fc720553787bee8a62a90237c8dcceb778a7295e15290c5f8e98337a2ee4b8c3a922db3a06a1d7a036aaab070967bb154f90d8c000e100539c66cbc81358e72fbbdd313635081dad04b9acaf68ce0e3a1652a8020066cdabc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h753fa9b3ca7b01cb9f6bf7109b49cd901ccf8e84ccf7003dada1efcbb8578562cd41f5ef3f38dd6a91ded620c4691347a5c0640f730d73254be5f324c073764f2574e333ceb1724345858476f03acafa4d183747a8a763a41a7354328a4614606e62409dbdc155f61eebfaabb7ed44f0f40ce6411980da21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7fe042c45ac5c08047b82105d71f2d4819b80cfc433754e671f09b49d384766ea7893f13ccc2efbf4eb576b2ae46fb11a85eb3e4b64022f09130b0dd3d6b7523550c8e924b916d417abfb100e6e9e3cc7424d5212ced8f86717a6c51712236f62d01839f9f0f489689afae23dd9b0d763dfbc1f606a298fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1759f98e54795a3aa9cc8404b933a6697c21d93e5786516e5eefecaaa7c2bc646195f538d93306b02c9c00a2bc2b0f80cc77b55e400dedccaa481d49ffada35c9a497576dd15a575322c0a454808a9938d2ce47521ddc8fc8a5adb3b473692efd69f70c311c2651bf7bb96c79ee3310ea16a624b074ba994b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c981dbb7b3dcdb61500a4746faafe2d5d011a0c43776c8a160e58ac88b81a8002958f1ef806a01bb992edb620afc121c34622525755000f8bd47482a9204e6532aea0589631b817cbcb71ff1a6f86b8587332e35b8cc99919a616e281a08b6964e147cde3d93bfa90daed86b8e5c7cf1f41c7c4c7841143;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h829de4d196735dd1a3c9ce4735e5641d9f5f82d9b70b3b834bb57b4f3e409c7721c41ee0e30b95b37b7a8a1cce04fbfb077dee62164f3fb7348ed60b9afec416bee4382c88b710a5b473997f42ced694205d7a9f51be1e7d34cbe8156db8ffa88bcc0002345f850d44f5183a67fe3470e1d939cf96da52a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e1cbda69b3f924615f20bf97bfb496221ca250dd487b162fc862f84387af0534676ef205c854420a3b3423ff9ed7dd51faa849bf69135ac70e581632933035e7a86fec1f9d0d064b80181a81f86cdefe7b2752d895c032be34fb9afb3413076d77778500e8e0ef95d35cdec53b0e601508542a683b1427;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f0db847a18bf5a05b7cac5db63738dd6f53f2405a9e9f548d2efa6d64547a0457230af80113a194bb8b45a2f34808e9d93d00fbd85ea558884d731050215c8db15ef52ed274701911af0f7b40e94b8c1a1f343fd899b106d5e6d6ceda9e41601446550118823c48e1b8d24dcedae7e9478f6ac6bf57d277;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h380ed040b059e3be456dd11cdbbc0e3b684d0ab8305dc04bbb08a212aa8c76ef44ecd5bdb62f058358e21f16b6e25472315b40bb34615c86f94a3d0b62779bdf5815445b9f78a08373765d8a2db809a283cbf1f3bc565eb56eddbf7419245f1cec7bd25b2dff9450d92b5bbbdec5e9803b2771e09537d2cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4781e458b79db61c4765795e1639c81aa5b559617d355479dee54dafe3ac098341971fe62618c701ad01b618ca89c5c172bd0a7065a72092458f267c48c73905108347fc5275f8ae0149a8177b7de8a18e88a43a8b877d3a9671b9efd8d96573fc6679927b4448b24e14119d14f8094f81a9b6cf3ebd5b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee41c79b7f5974945493446165db85ed5a8ccf6acf5fa3b4db8f43243736b603d7ca38c01a12e7d014f5e9e1aa972cdfa44a5ae1f48cfddca3a3035fff9608d0f392e6d9a78a5b8668d9b985d189062e5399aba825b9c2aa16bb240c94b51ea88863ff2090f49ce7cd21b3efab6e7f9e9f1aaa9579d2d2bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11105ef992d07769476530b5432e2c7182c505aec144ed6b123171eef389617dee5907b6de49f0a3608f2fb4f5de16bf1fb95af456a93dfe690f16275d391b7f3a920dac52b7b7e7be452cbbc46426f650877e38774989e47f5554cb470ec2a951584b3d65a81b7835bcd1c9ffe14712cbc81e5abe9b5815f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123bdc36312cd9ddcd29e24e6a71af0a8d7e82bb1a987103fa5a2379269c5b4ee2a0ddd0c9ef1b8e0572124e415a344f9285f406baa369f978721a2e041eb219108da475f56f543e6d00ac1e0a427cf867599b4563513653c0302c23f64b7af1bddee753bbbf6ebb9c2f14e618d2a1bd0f2ec834e561ffd1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h289f9d8afdf20b66aea1c5baf36d7baec002bc1461517f5746b64bcc3f2c5a19c76ad524cf747ad9e6d40f0c95a2a745d9f091678f2f3af7033f2dc8311576be373bb4cb615f6f5fc15af08f3a83b76d2671711a69586942f8ef43bcfa11540d5c98cea4dd2b1773478ad9c058f6902e2067ed3a7d4e641b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1c3bc4f58cd082b69ced73aeb2af2485bd043173266f1557d6935f0ffdcca691ddc2a12b2aee20db09f90398d791597a0fa5a45e93013af09b81b19a0564f9fe402757a249414b21b006abd222ba34cf0200ad60965ac5edc6197ac985c11bb49f0b8065988e9b0abe62431325d0d38abba61be829538aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9d1148527ddff6f2ee4a51bf40d0a0c25a4602feb3685cc44a144b247fd4300e2e13bb916a1fff4696f73e2a9cfe62b2da7e2c7b4cb11784a7d9de18afcf842e657302db3bd149c2c22eea41e839b4f145b48c33108721b6f859bb055c79748b3855612c0e4717d760cc3a2287055f0578eba910038a84f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d8a346b06417aea311d2631c540c9705f6ae2820a79c8a422e80d8fb03f34abfa49663566b2e48ad87e9fd12ec04d83e85b94d10a91a166027cb854aea21a0e097960583fc0e4cad2ccf393e8b70387ea45aa070f24a83fb2c158684e76a053e4575c2b9711361f41411e953cd3a759aa31f408c985e772;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136c4bc57a20d3e8eb112ae7594dd070448f47d6db5f66dc5bd4146cc9afb28878e34521b159052701685c0d57338d208790527a4b463ba0d6e5267ed9b5244d8bdab53b5b593427dfe3b01de015ea482b009baef30d13a8a24dfdddf561f6507a4c0f177e0c0f28268fb30470e1b3694414c5c94318f2703;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ed86d71ebb606f7b4038d92d51cca5ea2ea92a86edfc3a058a10231b0d492634f0cdaea2eadd0f2b940f0b13ac6253a4cf096625b8083ce57417268968187f2648445a6caf71d548be94da48289fa2801b240579c487555f3573d095a0d7f3f722ba1c33237f00885c4f058608a11056bf43ff7554cc9d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19935399e1d7bd0af88e9760f8bbd49bb35f5ca15402229309d39df067bed24e416565c60fe9d395ccd248680a8612ce00ea33a470a46d4b7ae19c4ea0f55768730f8213339b300bfc7ec8408f3f7505de9bbb088ccb4a80a095ee826232a277a34c1c24f73f9d5618884a3ff5ffecf0b048c850d2c39dbe7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d7d06fa36f4e86ea472805eea777ea96fe6687b62923a36e59b076f5aedcda9d92450a3db08205bcefaea9897df6f1217bffc5d131b8ddb01285ccbcbf393b252e64b43bab3db6a02ad0ded81e539083c1ada5a30e6b7a0eae4a4d94544a65ae09c61b8d9e7b0587f56dcf78b7d9d4d7fc115c395d39b17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7306fe46f0641ca40983df1be90d4b8bbb42867aba9fe488a2169069078a773502cf4a15c782531c8bfac5efab9a417e930221a1af452c1ecb15f015bb3136d3227f267fafe8bd6e187255dc2924988047d3346864ad29d73ba59f3afa85512674278095b1f89e454fef297bb0266822b1c77f4d276949b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2dd3b19eb5b078d9bec8829bdfbdd6b45338938a78fbd62380beba23794ef8a4065d36d7c77fc03eff7ff5435e1220829aad0de5c5f82a794c6b6687f32d205606a547e0ae98741febc1fddb9d8739b328a575dda22b2222a8d502b2512d257e24efc8637024cdc759f3c5961cf8ff97646bf5ac2da8a6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h450cec516c9bd6a40e068fa099f996a6eeb370e09877018aaa8ca3c51bff61a5452a7894946eebe3f5b51eb9dafc8bc93d4e1185de064fc0f741dcd76dafa21182aad09e4bbbede85ee6bdbb2c6c49c25bad56f662abf69bc7bb456f736fed2df4a7c061de6415cab62391e462b165e280c59e385d245f14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12edac2e50b0be087365f8f314a4259bb89b7bddbedacb71702d8883e2d309b857f9bcce1d497af720dd6bce83fcdbe176789bd251993050bc9798e290135ed2c91af7e329cede1b1e9ef10d39867035aa6bb479c2660f03982a47cfc1e4fae3f7a37d8363e722d309111d89018798417cdb4e008dd842e90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h217c13e109feb30dafccc4c1c17e194d4378023dbde4079b39fb5b72f0a3f0fbea310243cb58d85858bfe2f58e3c591262be5754f33f11ae81ffad4f3d76b484324fa11469245a038d0cd6091493a62f4002f42eb08b67ec28b3c14d88e6c28e3ec09bfb6d33f735bef38fe5ede67ac69bfad7899dab5f03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111a75cca5f662a94d671cda8f89f27928d754095767cc7e397e1740706dedbb01476eaaeec808c2a98075ac1d692adcbf54db5a78ee0653ba6014fba9e0b2d6d7385093ae3fb924b727992270f2828bd542c62aca0b98d0ef7fb326d27cb20424eb2d70a7e861658d6534273a673ca690efc97d4ee4dc688;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b1104d189fb219c657e8697aa99182952ad3d4a42ea9045660742ef45f58e52b88ae8800245dfc809ebab5113f414acd425fd36851d0bcf00f5446019afcdbde82327f755ffc801f443d933ac9574e4e1785b8d353bf0dd58f99807277d1e6dc83ef1a32e190a6ab85409901672ed3b915244add9c73ec1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha11eb8d463d3197abca0b42f203810650c6dde9a80552cb474577a2b53ec2aedb4bef5aba5779149ac14cb92bc394c90dacd1ad8f645a9a8a3bf4ead3d75e36e7c04e12befeb4a59473ec9c6dfe50f29261dd5bf7075f4d587941030328d2b9a53c671859dd3483d63560049d739eaa3b7e770ecb49a1211;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e153429fbf3332d8bfee8452730d437f98d8a168c138a18d05e8e7164391c5408b6c96af0f73567b5546ed1aaef10a3dd5551959b1f47dbbe7e6d883fba49f2195d8472ea444010ad3793a11135e6bb332e2999c67759b64d58e7c972e031641b4df5543fa79b35bebe74aec84379fd7004fa83ffa5daca1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf66c721bd6cf7b22867ada13e04f88f872545605500ca0da00a56d46c79b0f6961210d5d64399771378d41653adfc51c9fe5d312091dc5957da620fb824ac8af2e56c9dc814288d478bb5ac6ab9a371e294d0c01fdb7b93ebceab1732b185371c4cfd87202098c41d3cf0abaaab433128f66b0095971cd7a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1026915cbcbd668e672c773606cc2a47d32972562b5b973ddde2e664ee49fb364a2b9621de86fe2ea5315bbc19376ecb36a5c9ea24aa6de6bea04456a4a0d5467402d8fc16205be5ee48c5476bc066b16298333c3a74dc42a47fa9f10bf70c5bf9849595160118e99df760da2d7e982a41946171838b90b5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c14dd9fc5b1c6d10f23651b42394f70da2c8883ee0c3b2b27fcd15a31dc595284e2be39ff9e629bf05e3200290dd3641080f057fe8c30b2f806bb392f93ff708f4c3a09ce21017fa9899054977e694696950093403d73a3c15415b642eed3eb5d29e56329ccac3bb6116724210772a0455641c6cf576c3bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1288be3efcec6749bb642d2729a519247c994705ea84c83edd37587d325ab536b8c176cabf1108baed91092d3c77ff3e22a418cb7f7dde8759a888cc8703d7db5dc7f9d62b9db52980fa494de433f08cf0b131dd8eedc05f580ca8fbd985480703366b2a80dd5a27dd27dcf608d6c37a403e70b4e265cc1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5454fa2d8e30dfa3636a9dec8b904087fd215dd266b577d3f5830889e2d14463eac608035cd5867d4a36093bc1ab042e724471f556f545213d4552598a44282f6e2d0028e1f92da3bd7a5a9803ee7e22606b1b1314dc25155f8b5d5e07dc87898374643a67f437f34080a02e1ccc798ebce8a93b180daa9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h522922a93235c9b35921ccdf0014bd4b6a9a7db5c26d4f9f1d6a96c8efa4f795f4490fba8fb63e04d1612e5e9a45ccefe11861acb432cfc0c124cd344d2835285b24728c6e21097bc7d1ba204ca58240823a158ce81f79ec68fb136f65c6f19f1b94969888deab4a6ed7205819e934f22eb6d06b9c114194;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15817dbd4c2cb9f126bc0690da254b92f97475c673509915296781633713f8e872660c02befc80659daaf168c1daa3a3633ca5bd61074f441cce8f586750e6f5c1c27010187ccf537ab3c8eaa5b36a2701465e14a17a8fe6c99e1779b0f8c171de3f89698e51199e627a5ccec6f959bc8bf961019caaadc7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1991929bccbd60c8a5b120102c32b1d71009db694a33a342f674f8769f784a8d1ef6c1d1aa9988cf3d167437bae32132e1dee823d7a4da719ec390b7843bcd6af87ac68fa6a9c6acfe50ec0256049d4af7289cf1c5fbd1c09dfdd8cef5cd9e4516f3ddffa3027f004a0fc672cb0b279867353c83fc2db33b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebf898cca5bfc38b1f58cbd64e3a367fdd376fd0e2959486a3eda80b295246c0c8ac74fb8f2a035a4f29f7170245f21a4860c2f90ce1f888247cb1cbf66d4399a2b7661f34c0beb101b95d6ea297aa2178d30d0ba4fe4922fc195abaad8a91a4e68bde1155ea215246dbfed8f992d5a927d349bcfac901a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11370b0eb85ad32d4ea9cbf139112ebdec964a0307b7ec8b6ecb97980574ddaca4ce0445ae42fb6f6eda0c4b564c4285006aacfae56564893dc807ded8c4ea8327e168c6c159cbf74e4930c6b4dce808dcfe3ba6d1690d2311d7ff001eb5885a69c24f5b748d6dfb289859fdb998f009577d1a904ad8fba53;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf551911edb1c7a9e4312524f4362a21756bf13fdaa2e539ed6f322668a28c5b083df6f5232733d7eb3c96c6ca5eac722fcda7f6f9c9256d9aeb44aa64143d19dbc682ccc1d8eac62be6751cbf7a046fc7328634c110bbd16b856654c14ca58e945ea8e70c06f076a65f9b888c64ee97b70b2fff79855333;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5a749bfb44f64f756c2a07eddad1fc9faeff3a10093ce6750ae2759673e70d3ceb28b388acb30b13f35213cfa109ca69da9091138b48fd500e55b7a27a5c8da470eab51468dc0f03112558b8f6c82c7fec1b1b9eaf71c46ee12160bea8145771bb0485fb037a92ce21f24f3dba4c75cb018f856a73e8835;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6612e8d0cccc9264a67ea6a127bc224ec75c71e22462569c974de166a78a5282922b84947cc125db2169f9a11e3fe732f898c1c2106ea5112026a4d36ec7470f4c3cd59ae7c56237cebee3023a67c5ba5352ce7436e8ecb3535dedaebeea9a18073d2a7d578d0196302f75ec6a86a26e6048e6839f46137;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132c27ad7b94832b7e6e06b3f11a0333e8e99efc15108810adf28000a3e2359bb63bb8fb4a19457a1663d3b58d2a5bcc2c95945528340632639221601fa6ea84f16a2d20a25b19ee36ff4e0f50ef16b4f36d34bdb391095bf90d8a150420b20e9e836d32922408a56064defea3e64386a9e19abc6caab8c81;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1608d71458d90f0435472364ba376faa1ea98bebcab0802685909505099bedc8bdaa51a747b8b5547a0a09e83b39b02b7c6fa13bc97ff7090e64e2703a3386091eacafd46ba17cc740cee375f901d9adc48290cf505383f2b66087dfe0aa6e1ec12c1100dd6939a40600194a88232571e1512748a793cdf1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194df8f38ef06cec5132a586baf5ab68defad7418551a126f04ccee67577498a3c17644c06ce983910b825e7fdce2e1b7e6221fe837a135429cb66a1aa800fdd5ccef91e3c2b467fc377d9c46de5e01c9324dc94b0b18835f4a9ef08466a8df2d7b8fb4c3c7d522dc4558d7a7d98c5ac523bce62cdf92d0d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c4c4a62d1389308e63be115836dd1033b6167ab0861810108ff8f1f4566ca98ebe49dc472b58926bed73e6de9edbcd24875086349154ad6b298b66f1f1c9dc3cb2dfe3aa6f5352e015e7d5429066d45a8e08dbf7da0b5364062a50af32c47bfeaf7650ac7425037ca5bb1c7358bcf13883b3a7637ecbba2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cad090b62febf3954e1984b22afdde194d1343eac2b42046a5893bf790955421495a46086bec0e0fc87a869c10c37e828e983065e63cc10b58915b84f75470605c57fc839c373571aa5041fc7f77a8c117163a597e72413bc469274e28e226fbf5023daecbfea4ca72e84e990a5b6519a90786b736ac15b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b281b3c21a1c9a899bddba05d17fd4765daaea5b1a47697fe8cb8acbb3f88ad9c688eb78c9e82c1eaeb94fa2134c9cebbebb6bcc85ef6a6c46edc1dc58602718dca3a3f49b47e4538d62482df6c575dec122de9242506679227f26ad0955a72776c8e27657ddd2ea1b291a07de53b87717de6fc74b007b22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147d13c774baf4d19bdf99b038ba6578b61cc06a2346f4da65e6b96329a459746211fc79e0570afc55c38386dcf492d92aa36dccbf1db4cd54b60dbc8d8ab449624760c7a98fa40dbcdb4435e5a63313f22c4a6e45f5f7d7d6823f682d5470d9d8497ff583729b00d75e16cf88330ffddf418498190606832;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7111e45726285b9cfdc2e3a3091dab509bdfee64b4d5a74b4b743428589613fa290312e856aa0e088bc8789c2b8e88a5116cdfa69b134e58d836ee799dc2b35d5a44af328d86b0ac4fe07778968aee60e3b869a9b9d5b5e4859b1719d8a283b714a85d46b9387f895a16c3e4f89541c97f413108334ef83f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65c546a3a4608ee3513561597e037ab468a1019a9cb75680fbe0d3d72aeca20d740fec6a3427881c7fbdb53413fc640902941a1f6523ce7b7b3fcd26e8d217330b62f05619f2eb50cce9f3738d47bf0b20d6c35a1245fc615d20e36cabe6bbf386db8878976c47b9586bba28c575a242c8b14018c8f9d291;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a887359fc2403a9c74d682cc48e5665b310af5a4b2784955c46ceeb585cfeab9b4d804d02e624ae405ddff1585844862f681bd3858c9015786f5d9e0ff8f9cb58d57a1ed3d1a8cba7c7f0eb54c0d85a878f2fad109bec0d7ce4113673d8c8a4bd1089279762b467d91d128748bb8d9fdb89f3a8073a4727;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e94881753c8a8bff7951c4238483b887ff7722a6265136f35cba1d429d132e07ed4361792e9a8e0fc1d78e7cbf8507c340ab898ac1e6a02e222afd5bbc43b58f4ed8c7c16fde8a3bf1001b7651dd7237a48425700b0619e9f28c45d5ccacdb393b0f15f9f92a4fd8193b6be51fa72f52ef6dcb14ddcf3c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda24c821464e79d9179871233125e07d5c440434589cc64027e0e38a0013db7debe9c41a7bc9964873be8cefedbaa24cc8642619b4d5dd3d8146601711692f9aa3042baf6bc9a76a0661bd11ab84decf8aada1b04d7e35ec5b122b04bf47eb5935993b41f7384b85f23bac6bddcf78bf13e4ed8cb90ce921;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cecbb7dd040785a859f99aec378fbf8bdeb865d75846634b1c077346a81722dfaee1345ffb31593d3600bccfbff3743bce795c93ac61d3de0c009ed64757bce59068d05e1e5171b23893e5c74ae31aa983ef92396fc388704cb199fc60d6f134acddf4b0f3cb0f8250055038f79b29cb15a91b001ed6237;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he11c7461e2b22810f0bf88cd33ad326db9f905778effdefc0f9f462e818f329de25e62bf2a3b9faa2457c4f8188168319cace991245fc1c8ff00628bfc24839f717fb4841f883d7a33a0bd45c8022e89e1a1923400bf7f29a8bd8eb70e7364c7797c37ad6fab03ec21171ecd57c386f842f68a65ed3f26d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be873cb703d266f050e906d60c17ccc3d1ad4af1773e313b38b21798d64476b2582319b00446939c5c021bcba109ffcbb102b8246c12c281cfcd308a95b0aa957349068af3b51cbc4b63ce87ce49e7d19aa226a607318e36ed93429d224652868a4f3914daf5996893902637c44557069ab691bb151243e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d93ba932709c09ddfd4146ddf385b4b8af71bf8acac15a95dd31cc3d2bacd539ce6643fb8400e6a8610ed2bc2f5416a963072bbd2c589528282ac0fb75c39ea68b1851e1d85f42b505819c9b12e838ef6cd669c7ab7a78de555751639da49bc064ff4a509a9829da08849abd26573f07dc6969881aabb5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd61d0b9e9eb6a2dac6ace391f193502053c023f56519431f739bf6c4a41325618d4841f96d1615c946bd0f94954b30775ee5fc93eecacc63da1519c9c09e08d0378ccf80bfc8caa959649fbc921afd5229ab83edf90734808ed6438f44082f8c1947be017a442c22db75d6b68e235ccf84b8827b1410625;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h522725fedd9ae8c9059229b108055580cb1236f0518369c781ed1acea2d9c6bb9e32386d2ca63bcfaf937b884278c82c56c1399fb4a7f75b6d0ec05cdc59972697ecabfa1b2b0ef05663da9f5d15ff1907a551bc1a4ec7764f1a01795187db922f2ab450ac08dafb5d41dc05bf2ff4bfd5c73fa10b034e3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24d2baccfd962be9cbe32dc40e139e987ce91347a9b27661521c05c69232f70269e0329b8bdb9ec80255a279ad2dbe1eb5f1ac9a5712642519d14105d9ce0e4ccc121dc50dd7557db37204dce3af91e76ae07b5e94dd0fb221ffbeec9b67edde36c6f9539272374b14bbecc7fcd5f613fc82808ea31fc522;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a601f9e9f93df0efd98a8402000693372068bad56ce90a56c052412a02e48b49052002a429a6d7e00be483a6b51d34f4389445b624bca6fca7b77245cc8e0846c6c7d8c683db2d7fbaab1aae59b01fb75383968db3a294c49601ec45cde45ce550194f3bef491df009ae29b2227d2c9983809f255d7850a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1476af0fd1f413febd5c4c1e1eeaf3aaabfa8a3da1862027c8b4bc982109c38aa8c4dbcb7a8b4f2cf8083e13bd27d5109d44a44fb94e7fedb5368b3e6d3d0d74d3dc6d1454c2d4455a92ba912768c22efd9d1c0f527b13a721d062e35c65e130d0270f4aec63544d8197fc48c2063224b7ad5f335154c9c5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4f3e481afce64fe0a50d795cb2aa745d9aafb2e86aee07c4591209d90a15f8c0d8997b7c35904d20e36da0b42d957f3e6991232cbcfb480b3cae083980b57ab11a5303d088a50c51f2af1f8957e7db7fea10e35090e431aa9eb092d3241fedcdec2cc7e755fad79163154f59ed317dac33f060bdb7b05b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2296f51b9746350e1e12abcf7ad4b3305c3dcc59629525c2385a0ac305923d123cb58ce93544f49b5291c0f61a78b5144eaa10271cfb43063bdb704fa2f93913589df17eb1a0fdc291034d21add438bde0932346bd1cefeb7dfe058ac24aa5e15ff39a6a5da4cf679f7ede262d1da33fa814c0246e322f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3d2f9c41248cc573e12cf530e6f4977380d4fe25f07215079fc5ac465da2ad44be6f8690a16f0324d9ff813033d3a04afcb7d16651f51a8629adc0341634991aab7fa7c4532eafc0b908c6c39ad493293ce2bb844ac61a6a74f3e14b6fc86b36dfcd23d4bd8739703c62a69def17d82c2bc14a8a9f3880c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h759a3c1151aaca943d668b200cf29062ce51a03b570514ccad6d2f33b2cd500e330594acb58da20256ed512bdb47c66de33432e22960fb61e10682adf99c8e994cd3aeeceabd2f00446eb14c4e861d60daedc9b10c07215ba535f676c643c8e49e7fff6a39018fd4d25d26e9f56b3ace9eb0c30a4d300bc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcad499989aedbc7ea65e19334716a5f0bf2491a2d21c90e51f7524833a81584d7205d8ccbccb9758d12548fb15d7ef883abe9eabab8879b8a932eb6bb2dde28dacefd3bf1830ce73743b68b3fcefbffe4ef2f44edf6fc0b48106bd2a75627cf08c401f89a13d0520b8098ca71f536acc398b6095a1d37e3c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda22303fe8c24d472371ffb48a657d4ebfb9f98d599be45a3936bd237641e124670340ebe40b95a629ddfeb4c66e516749c585a25618dfeb8da0aa77403185a655df34f5c3d38a0e94f40af1e4c3d773dba3339b1d6bf84da02a91fd70ce2b9371b52eeaa69cee58cd53c62bb52769410716abea8b6e04c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ccfedd849dbe604a7d4379aabccb027d1bcd956ffeadd6570147995b7c23682011970fac048a41342983116d979f71526e9b4b860e2546346775ad1737d47abd60e480d49faa91ca66ba94adbde1ab80de5717cf05447e2822d7eb4e2f85d7ba02e5bdb1996040a6c4069924f2fefbb06219b8274b85071;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5854e35e3173e4d4b29ff5d19d843e6bcef15eab079f72c9a26f88b313f6936fedd835ad6381b5688206939fc06ff174aa1c2a97afac8a25397d2e9c1e8515963c8ffa879f790ef45da94ec4f2a321e013f94ef5015527052dbe9101d5bbc693396fb446d678b176c2fc2b0825e4cf56413c9eee28b95e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c6c950fa964f052dd86f539e6e1d5ee283be27d708ae9420cc6b5b4fb6cdc4a27f878cd52c4d927477560fa1f5a3cd6b4d1012d557d057a0114bc5908a688b1dd6b7165c6f18370cdc385e5f730da1df71724ca92f2329948715e5737c481117bde6a6996c2121b1904f77c413c4a980a9191764beef38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecc02f093f1c51dd0ec670c844f9fccdad8daa60a9d7029a8e160afa04c8eb5472304b17b8d4b78741cb224fd85a8636ec468dfb3ea40876bc6da2e4e0afafe8089aeb4b4748c3ebd61b868ae023e9a4333185a06ff9be99c04a5dc64c85c4a9f71d16b0004695fb58911c97a8f67234e63a82392c0096de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e55f20dc4882264aaf802976f4ffbfa7e5fbfc8a049ca9ede08cd71906b55304958fc7440a59410c3f3dd5bae9735b2ef71e1c5a1c27954760bea6d2c758940e49d3bb658be27749e0309f840eaf27d94034f44937697e79e205b2dc7bc678be5612d420b347b605a539907cfb9964c500f29e11a6172eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h625c4ea879162aa227f4d1533c760ea39625474561df6db85d158162239baf7b5bde115ab0e731964b01707e0fe79ac93d63981ab7a1c0ecc8a8a32c7e39d9e01db9bca65a0ce46b17889b5a1c7a33385bf3a5cf6f3ac8716fb24577ac2f5485dbc1d80ae11e92e90003905ee71d8581b5136103470475e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefd169dd4078d6855c6b2678d8fe9340849eacca6c53676833f3fa4f59ce65031a974cac934b23666ff41b6f22714e2baeabd30915d9ab704df3ba5e54c53b3133876e3b666c9223c5cd7a979b01020d39fc48517c4e14bb9f6035053d6db155b75b107387bdd65ae3f5e30cca63ce0b5b1c8fd4411a6e2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fb3c8d433ae4b7956a0efdc4b8035299e275dedf5e336bdc782de03b6c791799c3da256794b33646ad9407d6cbdf21c67b26c9ce345375ace80055bffa5d69eb0fb1ce3f23999f3310efdabdac0a74cad03a8716eabc4ae0862e3871b94f89098971d5ba4bc49a08a80a0aa9529465f5b91df3ff6b9bd9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6c546bcb159184e5eb62f02022defd409352ebfaa1b655958132d1b4e17f14af80194f722f538b13b67828d3ff30d0e5706fe02b414dc7461b92e8d61bb32d3f40616f1a2756c693dbef88ef0ff1c37916514c7c0f84429101b6e0b14e904154431ab33e27ccccbe7e39f80b32d6b2eb9d5c767c9d7d22b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f0257d56615ed11a75e80bd5e32b21f25278657ccc68185661a8f962ecafa86925e16f322bc21aef9f457ff66eead7cc2cff183bd427342256df9838fe12795f2d5a31cbb5284a90c89c7dff9dc8c914e648a2a368878176f443124f80ffd7d2c2e561b474839db8aa99eb0dde90266907edc0482fea4d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb644b504f4c4a2b9481b715a8fd3cec79618b2933d720d67f22778132525c449e212ab422b43749628d4e5708b9dd017046d289c2d3884810261dad630c015318d1fa1b19c87b057eede38f298419644f6fcc5ae0a9ddaac66cdfdae2f97537de27876dadd81eb18788ae3fcc99cc9e25e8c8c23c1859f9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h240b7bb893e6313676501ce5b13db9739427b5502fa871accc1a83991750fe7a5ebbd3700411630aed2a1199d7507b2f849484d7d493b9e24d7e0c183b9710d8f713ef32544a408b6fc5e508ef42bfbdef17cde6a1a403c9bd3c912386ad990489b57ea4a57ef473bd3eeb12d6b199c2ec5e2277d3973ecc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b6469472ea8831a5b534ded8dee15ca167a6e085858cdfe93c937ebd148b026aacb61d2bfdb2174de89bd024c933a9a2e257dd6d379a9935377319487d393f2295f4f4ff1b37b6e7c81da3ac1402c1681f5aa34a4b0a2167a59ca0ca8c9fd5db15bdc8c4a4743a655c253ef73f9276d72a006a0646cde00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b73fb329c33c74e8f09d6ab8e782133bc01f7a70b8ba4a83195647f8fdb7f27ff47c9e314e85db1c82908125e014221880460797b5ad24fd74846412b64e85fcccb410d91ceacbb99ea240fe66feeee402525d6ab955a0bdc3f9af2cfa20c64e6bd0d91a2557ad2172d3c9fea24f1c126cb7bd2b1374377;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c83203356e8c157109258014f10d410683578677daec628ba3ca408a1f82d103860b6dc128765ba43ab7fc24f5c80e5ed0793aba163cd41ab9950e8ced017bcfdb9200f3133c85259e35bfeeb07f3721337b4a8d712cf00558aa2309a9cc476ab544fef34dc05f5468e66977bb317976668a23107cf66825;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfaadf258ca7e70ba910e4078085242a79f9a246eac8e797162efe32e7df7c8c3279f606cb7f145b9b93d3c2145c558fd349087178e8c5d7f376b93a8da45864b5d4aa3123c1074594000a7624d1a099d20eb292921aa32462d3ecb098e2ae3569cb063bce63df3e75dcb751f1bb7bd1ffb0442cee7ff5bac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h112ab11cd5f5a88887cbafe6806e0eff1e0a4fb4b73a57b2be7d3a5116540b551e230412b447fe7b255aaf636768ef15c2e5731682e1264accc0afba9860f7a7f8f8c99910814369343c9da0f4935b41072dd0fb73f62b3d4c4630f32d0b7deac3101c0789d8a64bd54d13da382c399cbf6689174e94856e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e3dbae9bae8e3fedf77561add71091844ebbc73c1eacccab4f192c80e29b3c3598b88c229f4bbf039e2b2ea1efeef4ed4fe36be6774a24348c87799362e782159b7ce13e66c553c9cbf00556a1f4089e220765dba68ca020414d0c04f21a724867e22b185089c814c7c8c44d53af1ec393bd3cbb4b069da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcec643576124819c571c3c0552ea3d605e47d7dffad963cb6e7661c5542847ca893007d605b1ea3aa0cabfd0d7985a19884f5a6767711d3d395b428e348762b5708e2a207bfef48a4cbb36572e70e8c26626730fef64c2763caf600949b4bdd0169956fff6e2133ce1c62ed32a5360fd070e2c394373e55e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87d7046ed6a1128ee2c7a79457f46eaee58ef3a87bf855c3197ac3939fef5c7a5d3da996e1ff4698d30fdc6f86e03eba657d84598da3a66165b2cf423b6edea61615daed073b84eb43516818de0463a5414c22ff23443e9d545168bb193fb94807ea1392efdf1645957a0a7c31b7e91d89c80eee0db717f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3253b00dabcac002a980ebe1a4221964f2a7398569835e3847708c28d73c754272a9558dd67f1d6d61f18215e352dcb73b068cdad1b958f8f21cc36b7eca73473eda98cfe8d240f515b832281600f9c4461b0aecf8cec41e5988c8ae08a938a757f91e77a9c04e648b7c6310eeb46beb150bf544c18a83a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d939696cf6fd6e67bebc85575ba6a54759479b716c9f0b9fedb3d6f606faa79ee1cec2de9674d0bd1b619d8e91ebfd076b6e232d044bfb9aca9b71ec4f013f37f1461a02469384167d16048d24d154df27288fd545504adaa896cc2076dc631437359b83d5c096001bf02d88112ac4a0565ad43e5d51148;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f4663e9c166408d0dbed842de1a569c5d6ce20aa2959a4515b33e47dcaf34ff45ccc14bf0a588aa313c59d8a714e251f876b07df7c69353e2e2c806bdc76c9d3512ca034de62addb4402daf1fe55307e511c571af9b127a05f8c00100af34398a668322ec12d6ef222c25020c2287df148e9e8fe3a0b609;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3dbb692d96cbd1361a670db710c8b77df921a9db3fc425365a837d5da7d88564e8a1b030929f6b3be615e29e8f4899eefd471f85ea739cd5a7ba65e7c7a29cd7bf36f8b5ccf6f6847614332e0474e49a40b65de8da503d060b2ad571c1f24ac240f7c6a9fbb6624cbecc12c1e9c76544bff343de3d109fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183f9cefc4c492e301eb0d5f83029270c274ac5db237ca67e3be8f0597fca749cdbca81348409262713f0b9ce03a3731a1867089c2a2b82c5ef58c0befcb0c1327c8f088fb9ca92395794b5591c1e937ec2d3a10dfbb12567d4288b496bb9b10b4546227592e2b0469088d40b5abb7af535bffd4139f05644;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c6f78b7c5ed0302addc04afa77c726eade4284d2f5fe5140429fff72f8400b33a060b2c184044d072c32ca67e8f1d21a4602d9602d8bf127677e53ccc931462c3febc665997a0d64d56b420c4b7613916549be9b1e59671dad62ab5b70d5eee7e9016f7868ad7b8dd5c920b3324795ae4cdcfc9860b5a51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a95ea5c7ff91562b59d9ae31018df0b1772500abd2c87542de3928a2e005c691e63727c997634a5ad52e8eee0c34fd2a963cf77cb220dbf489d3fb228fc2c04122d466d5e949d8e1e64c0272f17ee0ef9371609d8969da91238f595c2b5730ce673c0b19b869f6e12b4e56728417443cad3f3073dcac887;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he958b6a8a8cf417b74f60997e74cbbedb076440df4fd8357e45180f435737cd1961974a7938d32d63f2c1b1aa48f709e996ff965274150a6072c2ab354a9180015476945edc1c454c5a88888c451ea1b183b1647ab6eb08c56a8322365db9082c88228729c1c8ff010137b25300e2a64edb5992c6ef4f86c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79b25a8e8541e62f91fc1753a5cb19b7676664ee7e1ac0d49ce360bf2b1526393ac2be834320ed6842b28b7b3de2c74a39565cfbab231e44af495018568a826dd67c0952b212b496917e152e749e34bc0826336ad130692989d781400ec2e3744e0125cd395b3ce881cfcb36fbc64c754259d680b218f781;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4993132466aa1bd4fe6ad0bfaa9254415e48ec611767a06df31aa278953ac982b56e8516b758a9de0a610ff6312f6dfdbed8bcaa9d3c9132b3ec0886168952dee472f3edf4e76f86d33287f50d051a51b4aa1df23fc655876a8cc5e96427c30c4da75a314eb2a27118e66ce07c73773b31b5d150b296d01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a066a1ab834bb4b9df54132e981ccdc1d9c87c92a01b09e00e498cde7e619b6f6d8ab825b0a9e01c50e1a06f8edf5bd5a780e7b58d6937cb416d518e47957a0346ba3b29322a77abc1aa582ac289951220a9ae3052bfd26c2f31826101c8f22c3fdafe0848e0bd9248662ee6e1c439bfe3046057b09764a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc71865c6c36545081ca246de9e6a876a410c0cb15f33fc897733266b65c5634c9cd2052a97a890e5960685cdca6ce35c875371eba0fdc2c804e04064760c3d26dfc3f14d98d212c9c84084561b4ec585c6e9b01b7b84bc4950f53172526f695fa7b24e0327ab8279bdbb1f8835fe736a8afeb78fd3076cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f27b3cd9dcfac17e545b566b54ddcf1f4a78276cf6dd1ebc0b0829632c0db6733688a1a1231a1ff1fcd2cb8ebdfaba31f7262e302173f3a39d6ea91d87af8669df87b5325bc58fe35c7789cbece11d9de456fdd261959226cef99de1f81f4b39f0637144838313ad48d8ae62ff219caeb2f898b79464543;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6c1ef0e1d4654fda987887455f639c1d1bcc9604abc40ed6c1e341aedeea396d8bb374787f3c6ab75de72d04b4d4e45b9d213a7602ffeae3de757f6f9dc5015a9bbeba16bfd317ac91dcab82ceb5206639763b73e079696f2a4fcf20b4531e25e55a8b6ba968d5e88c71f66812e197f6d27bad9dfb18e66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120bf30309c071cca3b0dbe642bc828b255bf9a4fe22945703f1b310ff84634ffa097bcfa3e533aa65f24ecead205278382b30f2f8da80ec0ee303910350f2434f664f3653f594ffd17c018d59d777c7024a30240136c93a9741535c6b4087bf9dcd2050d3028c5e720f3d37c5ce0153f7e5a1fe494c46a0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he932cfc8c7eff00bda9c8d0733dc9bc31cdb00614fa484442574e1d03053e05d0a839b1eab2a95ec3cfd96066b7b39629a8a92c88d68a48fcae9b343635f3560bf228f5edb9911cec33b5b7f8e17df52cf4638b580c357d85d03516eb36c918beb4febeaab3eb944a26dfc8f60ca84cb0330ecf5c53b1b49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b27f7044ae88cb51e520b0400bd814c4c24bdb76bd25136b0d5dcd79e4a5170918b635d47641073114ec08ae89481a2a16ea0cb88eb5bd27340de90d3131fb87c411c4562e68ee425a619e85a6b05b189a418bc283ffb83c45ada4c49be556332d94b48b644cb3595a4d1a8b12a889c64ee30744d571d3ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc4d65c0b6bf25289e0fa51dbe8327687ac57e35b7d0a81ac9f87f337a8707f2a3ef299ead8f36ce8ea5987e05b0a5d8ea6f7a5dbbf09fa3ec01fc4cdb2e3b05a7433b1fbbff6ef7a8f7447982a775bbd65acff22c67c230b48f1df321dede8f9908ca4446323fbecf97353113f76a95b8d2a21614abc11a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e114b48be230b8ce9e90f34628d27440b5ceca339c5a0e7d8ea5483f00ce9596da9ca287f73267fa53c626e40869b7de849944523eefc610f48ca97a26524b61fd52d6da89fcbb86f2cd9f00e3cbfe5bdecd75ee567a9628c565f14d0a36af06c99f2ae0f36dc0087d4ed36a2999013374ed3895f9c8d7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a308b517f9c3f5b9a2f43b20bedc8d41d519fbf0b31af26cf8b510d31567d52e0d518826ca59b06a45c40f5af36a6f58c00d6be0bc1917b34587afa4b8cd0c64f3335f4b7b75e0375cf7eea2f4b4c07580b3da8de63d2a3d8beb9f6df6c4036b0d188cbeb5865f7d494ae382a14c0378a14fe191ec5d725;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec2f5ffd374eb77e30a6fee45f8551ff63a0aec9d445c5abd75c396c25039795b237bd70f0ba594473073824ef33cded52ecd4708350e8a7243bfcb96ee1b2be300415fb3bbbef23deb74b71475cef3d73f34c20466cced48c0d955955b42e46b73282ee30d3b2a43505f09cb69b6fe5ba7d7774768d7d8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11707826cd633be6cca9e63573e97df39cddd22fa836ffb0e01f88f3c6624574618a772e0029bbc5ed240f7afa923208dcd040ffc82681e84b650d17d6b86ab995b01940b67565208a5ae7f81c2ee6e4d03478c9e94995b8ab0c2fb322bbb370b329d163e9abeeb8e14905dd40606dd090b0b4234020287da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6d5cf2351ae22c7c88d594356aa0d98af6a6a9af2f0ee996383cbd8e07358109192bdea06015ea0c02b8b8b658dcccd8841ac7e16b92c7b72207539bbe4c09770850366f5657dad335744b8d11911752300df458ea414dde0dcc71020f04908d0abe8dddb6f64a59ddef5b1234f078ea634b84a19605ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1537a3adb871cb7bb5f129cf77ac01d6f88cf52a9bf5ef942e1ce03b7da4fd4a23a67ff1c531be3e93d15c550c3b12bbc574f972f7a609e26bf4af6ce0e2ad389f7dd5c668b5e4ae59239f5288989b04c022a04ffac36c85f87ee20dc50436d2999fbeea9abdbee38c89a7574d9345f33f5e101ecc9b38490;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7849dad762d9b5f6804acb32ddcc70a9c01ac8ffaaa4f3a1676d24b2661d672036c39147547bfdcce5c001f0fe8e517083a71f947d1cc37b3be756c3ceab0dac3f775bbdd05b433409cf9d0063fe11ff874a66eebddeebf20cf0450ae33bd847c0fca825a0b20b0770252b075f721627bf9c0f33ad9442c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5ea94464cda0a0bbfa3b362a70c4ec3247b5581d76d348964f6e92a37c9515a4551d4958e093d63cfd8df37a962acf6e522a7d3f1d474d3e4fd9f6162cff125ff94af05095e006e0233954e1adad15f9c26b44850195a4ddde731d7cff64142a0115b10a4a9cfa0068e8a80d5453ab80fca074737494d05d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b908d5d3c05ea2ae9cf447fe5dfbd5529dde6fef716b8e11a5bc024c4d7cfb30b4b5aa4354a95fea328cdd0ef7139769ca252e8c243affc9bcb35df69c0388cda3376424620f6149ba5919f61826a14aff5ad4885264f1cb0af0a3b4ea8e63b0d383775350a0273315ba36f3f88a317eb9c66974732827b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1392ee332f9abcd0d8ac3318a95f0a5598b3df270e8b5abeb9b6ebec1fbe802e97d09502a1538b347cccc67b8e1c084d446d28bb9182d4a8847797be27b5e62931f1a596a0b53e13349a801ba56e6ece2ffa571d267856ba13ee197141e749cd6fe497209bd38176615bbc4d63a87fb060a765f15c13d24c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5a7229877a5c05313c53a34ba1a95a29fe914237f6d4c15a5318ffaa54901c7173216d2bab2958039d6f7630814c7f1335448849a5b41d5496aedc9f5c9e7fa64b1aa5a0f6e8a0542ec1269fa9b830496553f4d2cbc53afb3800c5c618b9061e18b9ad9e4b57d72e2a96def9f7dcaca5e3f54200457e697;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e88becebcaa00887f7b5802eda99c245f71021a5e09c50e3ba8c85cc27bb05b6836a10911dede91009803f9fdeef8314b68e5802b71d38b14aa85ab8e3feae875a176687419759dd0887223386928361e333b26b086acbfd805ad807115bf152a7035ac331f4e59ce2bed9a51311e09b1ea85514e116a1df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8966e049b8087d674d16bd7ad1d67149654063b294383081b5251c5e0e5fab90c146088b46a4d8653ffd730e653cc362dc4cdeebeea2f69220c72ede1acce34badd80e20814eee8001f3c3db16b74947e82b54fb45fc03a9d8b19f1990470f45d66fafbc05cf87dc77dd12072333dda0ee04c986d45e566;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfeb5affb4f07138c0c82765799ce9102c69bab99d1209efcee0c0f802e8509b03bbd5aee52b06fd6a78cf3b2dd8e2eaf112769a0974014abef51071f8e94e398fe67071758c11b35054f7cf3a11d9698af99fff80ba95e674f800a88b57a33c1383286e230ea39b6f0ee0052c0f80a23c380c52c53db5075;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52a31c9b293fdeee723661f0dfa5f40b26ff8e3135e2c8dbfdc65b48edd259c47fbff764da49a1988b73b9cdb5667e0ec57cc3cd2b1fd5c2e64c82bfaa4d831808a0de599947ea684eba66081fe66e8652dc57950e33856cdd667855c4b55a0f34bd927cafdefd3cc18ee9617a18bce91e4f3a9cf534803f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edd7b74bb67aff6664736b8b1aa48bb394ebbac7f3c8015c2a1208a39a11b8ac2319c0081e1c9cb35920c3b027905e6c1caf59eb8934ccf114a9420f1f70b4f8b2334b20103d4a636a94914cf8b25928c8531ba68cadf1cbcd7ffa05b69c6f5d6d1d25f053092cf676fc963e6a8c3a70a3a929e9c8c2a57c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bfd2dfa987d3e10a765a1636abd4f2cdc0cfe8c4db7cea24d03da5bf4d7a8a3181fb142591eb67e3f0d988d76f82a11240bfec05102c46851e4762a99410bc90ade2cf6529d456ab11e1b22b174ed71f4a833eb1b3170b4983331fe1614c8973126ae2be0198e973fb951d1bb070ee39ac11e53c04b1160;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f0c9f77483eb1ba072f03892808c63f6465eb9ea8bfe122b21fc93ede14bdda3a74434064134d732cdd010fe76289f6c767e39805ab9d99b1ba83cef04c093e64c007d9573aa6cfd19691e069dd12e614a05c89fdbc9ae595ac57ba28480bd8ce47c3b41b0c4b6e6098a249d100231841628cf0bee9490b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b3d56698663b4a71267f0d2c25c89484de5a76eeaaccb2fa82434230c947c56a1a31f55c8ede865379806331ed0b6d1c4c298601ee468dc43e9113271e20e3528321bca2527401f5bec7f3633905e36c7b67c342e20751daa3b8ae88185b510b46d585318c79c24830f5d8186f81caa1a2786a07072be1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b14ebebe6b71e68bd016809c8bb954825a1b98e42deeba70e9e72a6300c5db3e4f5db8963aaaa417af0b081f330ec22747914cfc8e6c5cdae5dce10ff2f2335e9c8c6c743f4b0744b670ab75622cb9a22e0c33a08428baa0fd6e76fb19dde13012fe133b7adae0c6e2c0d6e7f38f543bd5203eae145b4a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf5949511b13523eb55ee82d04bd26c7dfdcd9bf49eb2aca1109bb892da6bdf3d880fdf63cdde4eaf34d02c2078bc7699307ab85cca3a00fbd822752bcb81d9a730dbca5a8649cd0fef516b4918eb67a381b395a505e6eaee2375a6554e14eef1892790a286363122687bca33bcef14610d08bf720810ae1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he205322c26452f203f788403344f82d0c54fab9623cd1bd0ab5c6a98d2e37d1d1b386d4fa624c70b3980ccba6fa6bb2450e300e7fa1e107ac0c658bbb7c31c07f10bb54955e42741a691cc277de12283f55aada81b9b40efbb8b3f017847e160f14592f85265686d2bdcace138bc8834fca1474593179564;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd48417b7625794505b97172fac4b3ca53cf0199762a0ef291deda5d62fcd2f78d835602e87cf5cf1d37bed3585b78391c5bf1fbcf973a4aaf004bfb9b48c9c2322c25bf096741b477cebc09efa15faf3ff0cdd5456dbfd21d36ef8bf5ef1de01ca8e9be3fe681dd1e555473f9c4d65d0de55bde30db6449;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c163a34205cc84fbdceec34a2fc6f44ede3a57e862b3e38e43221c91c81a1479faa45ae52791d2809588a95b8d8d1a1b70771e24dad1fce25a0e91a1349070b50474c1d673dd1df24ebf91cab12cc1798900aeb1b78f2a5e2e0b6d4d2324d9e2c22cca8f71e9ac7234df4e94713603ac31dbf93d0c278ea4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b92a5c5d99b437d3c1ceed3d288e2e25b17abb2c81209b59d35ab108af6c86091cb753b0dfe3a4439ad6ce5ab135eac92535a6dfb38ff2b328bc1fd63e292403484f2e0a6638d32ff459ccf10b2424b15844d20162d61322989fa68ec5d6fb072923bbb887b3e292d628d6e6972a456b593ffae011973b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84fd88751db62602ea281dc6ad95ea6f5cc2b49ea666a6385feed1e4a6490b39631e336ec4cfb01b9171a7089e44144e2d6582a51b1f8b5156188e6d004a68df809020798c8ffa32575d187f0184f43253460a52ce9f369a2ba2337e498f9c0fe2907bb6479337b783340da6f6bf1bb5878ff6d02e454be5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42dd4eb66261a670c817bd2c2754d64d9be04a3703e8233bbbf85307c2597ecad347d6300b2a2b8c2755159b99bcc13bcb8def43ac462ebbeb3c25ef8a9a1bf4d81ce2aa591f65928877a6d68214c9de8663350ca186b52cca0cf7a020900263bc5430d3f5d6c920463f404ce3dc12204e012c1f2ce78c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h605558de67edbdd316baf71455730c6814b394b50cc3578ff79aade11258b7c6d3524e2fd85ea3b5a2520a4d94a8fc22cccf62c69a50c9a609ff4f568a71cbb12303216cfa450c6938353690c0b6876e1d6a39749f1bd9019dcbfb7d1e7f10357ca72a4ded4c4396033d9e6351f1415233ab05b1ea59bff1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1153c0345b19b21a43fae345a1e89407d99bb30dd9fef86302e619ac66805b413c4f137e7e63e04155ef69db6e56f58ac0c6bd62a4adfb08691415b19899907d934a7f04a6f93d40d6bb312b3d508ee2248105f5e64235eb33a2405dbfb800115066802f24bfed3e5ceb288aadf485dc84a0054c865e95cb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80af06e6f7765998d2e4e6126494997659171795b296b28925bda3dc203452beb4308cd97d0091e2074613b7a83c212b3430eca95e32b82ad7c6e7f5cc7499a578ecd706f347fe15c907edf3e892885ac6125b0d000f6eaee49b272c53c1251faf749d0cf33bdb29c1a07e5f06a2e70d042bf6cab44219d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7490ad8ac607657861eca7a2d127a31a85586aa5d97c4cbf50ce3a8ebbfa253c90e98a13efcfe6895045021d72adaeaaffc729a2290d8bb54ff9a3cfb85b67da8ae6dd5a0b4c773ce2927ac040edf922bc6d10a8e0ce7c425fb67dc94c7475ce5f02da6a58d8cadb19dc34963b27277523907578c79a9c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc830ada970b79d7d2aeab63a20d807b6351fc16f13b7e5b29cb85c324ce6608afc3be8bbd95c61f385182024b85bddf347c6c2930b7aae31391b408606d714157943f212c83da9dbfad73946b4397a58fecf1065be02a9ec1c89b8db93ae419b2abc1ccca8db198696f0d78698fec609cb4b4ecfd17eb102;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1358bb8075950cba12f1ed6bbf0a3940ac10cf725cac8579224a05f6ac31d09b8281b00ababbad98f61fbd86332cca27e3857e84198f4accb5cde58aedb57372e8ae0913f20bafc76a98f6650a3fe6c764658097baf5752ba9b6d26d179626d9817b48be11b0dc450d46e55eea0f085c8d09014f372b4e311;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47b3355eee94d449ae6184850b480c415ad529b57e9d7bc3bbc1c6bd30c00826269a5bdbaaa536f013cb9ba401fde331a02b6280063a8745a860a51c1ca2241144a894f94f068d1d4eaa8d7afe9d308cee8a26d4c3eb41e22026e55798ae26ef0928a8ab6ea92ad62b3b2b2638f5edbab25cf4a970bce6e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b723aa553f83669820ca17ef535a0878a810b12613f91d1e88092e63bbda6771458cf5100351f2fa00db22188e84786a97a9b95f334a8cee1836f73e742f30c99df871061b371b86949230ca4b6bf42815791b4b50ee221d20b1f4360cc1e23c83df00b70f5048942ec789008d5ce57537d7140f8232a9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a470275cd8567a4ecec4ee05673d3abec21bdfab1ae056c0ed18d9ac889c88f70e38b59c9f915a497a4bfcdbafae7cc3ae0bf9359208bc067919f0495ed5f33d999206f0317272a7131ba90385cd532aef07f40e68a49fe2d80b24d5ea2f73f20ac7dd67728111dc56676f8e607df23c4ff6110a10ce8722;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3a2898ff9e3f5caf67fe16d6060f23859c0146cb465b0641113b5db8437fb3a6b0f8456b50316a1c79fbd7ad1d372640e17995aa26cadccda55a83e5cd81f1bb9c947e837b7e25a300e4a893d50f3421a36efb834554f16b3e20317a0deadbf9a89c05aa4e9d795f937859029d4e4efddc4921d2490a8c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf69ad8822b0a117dd834c5351946a53b422c9ec964f95d2b015a101540af3b3d05df25e8bab2a3365571c8d39427203f74be2257d8ad5364c36855b71563f03bdc1e99f670ae1b85f672ecfe25b88396d7853a20a5b7475918f38f5cdff263709c4a788de68e6ba9fedb02b3ab1848a579fae9e86aae7120;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b7dcd19d38959ac34e852a1a20d63b2469ea7b6cd48ae795253de13c67f52c0d0469af8249b6e5bbd1dc2b10ff021e7cca76a95466970c11d505f505b0361a0bb9f6f45fcf26fa6398971ca3f98ef423cb729c615223f0024fd73266a5394dc4fd4dfecc15efe8e0fc2ecd420c05c6a0f5f9f6a3d5af7f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18502f73dd8b9c2192e182991d3f1b6fc1f40d1c43aae3b48bb60f32f557732ffb7887aec85a7a7ed925a376c98b15438f84a8bfbf32f2ed6e99a7826951a7bee7c9e9efc19ff1cd9148eaddcee268163a70b3345dc69d01a4c01d1ce3ce44672f87606d06bd6d598b3c8f3e53e9628e463415b7f15effa38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fcfd63329627dd5a1910158185a4dacabf8992c1e573c692a75a10b62c3a8c4d9561212efcea4475e9e92c34e6191e8a2fe1f663230ddfca08b7391007274b0e37b0a9cce1700f7642c671edce8ce6650f935e4b40acc81188f491835f94dd9d29e3cd6cb8934dc6bfc1cc9986ca6299b36387c5336f30fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21491af058521d0dfae9893182cffc489831ee05e0b6e99f1a642b6cf81a04da984ae0fa779fd6a70997e6f2439aafd67d115f56a3d5383566db222a37331666a4b3dabbcc708ab3583421c8089c041b395861f2d2b08c0a6aa1f38e9b17af2c748ae20951f67bcf5b15a0e192a2f46cf61778a8e5cb083c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68cba4cfb5727bddf87dbf01b54ff85d41d5af9cfd6e603260137b339c7f9bb23522f43eee5661859f39bfaeca0135e388c90b7fe44aef95fe096acabc9818a7cf3d56a1c53c67b1ff24e662a023f8af1f94fed03108bc98d1f393e71e0dfed8790c008b7a177add153898d46727c927a2a294ae0d16c567;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ce402f982a815b6c67c016be87ad498a31181a05dfd7eb384af22ae61294c9390110be43efa9a0af2c6e7590eee40a89315fdff75c868054920f4bd76c10758fd51592a34c18fa7827e9dcfdec7e65e565d0bb65a3feb5ffa5a26c2b2dc1f3aa22d80259f08f86afd263b71b6bf3f3540bb7e11bb56dfa5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1444a93f7ab1759c5b3ae3a0cc7339bc4f67c8d07fb94c363a438e79d9f830a4cffe0f076c30debb62fa1adf40feb80f06818facf205faad2b4f4496a7ac8079151ca8a0af3dcf9faef4050d5bf0732f2c6ca78b88cde04f820c0f1f5edba5dc88c3614f9b740cdf1957e1385e90bd5ae3f7f5f59313fe204;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1611fc44db85620455d37b68d053623d00bb14b4b3fa6cb437b796e6e938e2d5568287a5132821ce83b0203afdd218ff0d40515f8120ddcd7194efe35fc906ef5b5f819144bffe3a0790e624e20a615182e7d712b3e8ee73302b982b7f53a740712496256cd7838e64e1a0342672fa8bf838185648dba7702;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd49eaaaa6850fbbcd95b87ffa4fd55c6a367f7b117608ff27785da14d354fa9386b7ab4529eba525ae93d8634ca563d19b2d6919de442da8e905b48c05d2a1e470fed8249f174050701380641bd2ba72a41fdb4b2e5fda6e1bd230caf32fda188b384b16afc9ec36319e9522ab7237d8faf172dbcffdc6ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf604e5e0598e8af079426c58929c41fffd920b530296db7ae51de55542cb080e9e6eefa50c3057268a886f267b24e59ba700990128cc2f979c39f5ce67c3bd30e73ad2a356a28140f4457aeba2252f9fef7362bf87c20774a323bbf726cfb510aaf39af85d8cc915007313922409e3c356f17604c15e64b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf16429602e7ffc91e0b94637ffef025989bfd14fcc3622048d320e7a0a3bf1601885bfa373ea8dc9f868467a91e97b2c7ee82d87b3aee3b7d4a57cc8db204ec51f24c5dfaf408a92668ad98a72be4ba022d96ac7d97003bae990e0d59cc90f769ac5eb5e68f3c0d950f85bd891cfce2209b376f04582000;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132099633769abfb49cf2e8a8f831ce33989c3ec45243d90e9aa3af584341c7042f3b7ce092155c669de8102c137cf954c9f9030beb8d44964e0b7bd7ec072bf867cd9587b3eb72ed5a3e6dd455f0b0302d0f0229b3654e3eabcd2de0a50df6384d2b47f39928b494d76146d7110f1a14a7d9c37520b51653;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5117219b848f074decfefab3db56723d49168b4bf5e83322ec942d90317a3c659c413889f77ec475366a1a6c1c61394f71d34c2959d1bf3e1806437849e94b290ef09e14c7e8e3e04b9ba547bb5ae611888bc88692c8d9ca9ec17af243567be183eb36af51e06b1a84dc5ffd5870fdb2592fe56bc10ac0a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75e7727116f19ba1b5bd1ab6138bb534e31687e04f1c6516ca3c3f34ef12598a33218fa253e173cd8fdbe1d6cec57e9128e0e5dade5476e253780f3bd4b5fc753714c9981c8bf13e64bc47fa2f6aceef14503f99d1c8f24df479c5d9eeb4c78a300da81aadedbc23612820da8c53cb5718b418bbb1528bab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47360fa71c825ee2e3085fda92c458f3c56ca51e636abf778d4a4076a34e422655368f4521e4fa0e61d497de0c2e87bf34ac9200581363c3386db415ecf266cc7fec8b978e62bd2df76d0610f14d303de2cae3b21cfac9f6742428dd9221a3be168aa3d4ad97ae43399d4276a748d0688603b2a1e14570e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62cff5a15ca2d205a94973c45c0594cdde7fd209ed36d1f5d2cd4050858c2bef744a8a5159c69820be98ab11326946880bf4496fb19eafb53655c10d4c2e78976eace3328d085ab892bd92995e2ae3445dbb3c94964b4079d5fe3a6f772073f2eb8cb6880d93cf5490313ad27e41b20cd23eb9e3e7b7816b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a2fa3e6c7276522e3b7c184ea77b4b4ff703a6ca74070bf8c4b65703184ad23a57ee923787721f7b505dc5b449bbbfd465563a20326fa1259e5e38aac3edc103f46fd2eacd327d7ddc614aab317cae9d9f68c644b62380bf9e6ede1f49d165a3d784d7c0bbfad4eb4ec13bf84c30f4b831034cd8b267bc3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha675de3368d792330b3e09bc79fef385da7c95cee18b2bc3aad12e3250c289c4939e41c090fc56f513b2b0c5bd0422e7eb36066516a6348df484ad282c89c4a7f44c8df3c5dde887d69073506f25df70694f28e03ed2e6c672aca28120324e6cda9c8fcd85055c2551374e40398816abdf5cf745c97e9d23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12515f8a0cdc63071db0e2b55ea404645bdd1426c7f0bb6400851bf70f04ba3de02aa1559fdad03aabea94b605aee22d7d2405ac441e67c78c6e65479c9c0460a6d5db6d5d2a5dcc9334c26561ce70dcadf0689a2d0536478bd6e176a097f1fcb5646a0f9473b24215a6f0bdbdf0ccf4ebdceecec1701322f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h330eb9686fd8bff6a189ed4300693b53df05ecf8a215d765e7240b4d5dbf4163eaceebf02871c61f141ab8eefe652be96e918db627c2a35f6ac4cbf697bb36bbe5596a4e4cd1ef78354dc0c87b06e35eb46ba0164b7bf16375044357dd175e4125f80db87ff61167e7ea6fa6d67a8d5753a4bc22e7a05da9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b3c9e35c34b068c987d72ce984b1300432723877902a6d2370565a251f5bb89183fe475693e8ea5f08a02b38f7c41dfe557875d03633dde744b92bfedaf76d06964e6de7ff6d664cc27290b04cc941781422b9802aa89068f49a17bfd2fac68b2b85ce2a4a9ea4b65063100b4beb066c494bd2b46eee798;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1980c291f6ad6ecb274362a3a93eb88c596ebc62193c0aed6716d2b0a3c228ac61075e1853af3128b5abb6e7ae1b668829c09d880e97dad96b4d4da54c8e16aecbdfc9690d7ef983fe5e23552257027138e142de33a4cc389082b4db054c5af9b4e8c212861cfdf2140243377c9b90d15bf82985a597855;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e93bdf5adcafa5aa21d1e5dfe2b6562ee6d5a51d33f92a456d87f1badf814474a940f9d7cd39595e30589a6c013e4f2feb9295d487bedd6ebe62e0d5eeb38b4bc2296cd67145773990d16075f1d1557b16e715cc47cc245e6209a2a16c7a06270bef448f3f47da95fa6340291ea265aebbab75674e90ef36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4daefeec0564b809544aead4f9e215ec8a10e1c05c0d8e5c0caa13dcec38babb9d1847d682ef1535fd8a8ffd8f5f5d93140f6b60f827f301837203f2bd04c270d7839b0dc1b7f788449acce7a657d057e3527014913cf3f04ded6833ec9ebd6c1e230fc2a42006329a167aebb282d6a6ee6ea115e3d3eba0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2940d114f4eecbd9789a655279ad8b043181a9301b737c1676116c09eab6812346362076be869a1ecd34c593b3f0c368c67d8de91a21637a2daea890bdb8fe8915bd9538369eb4565cf48db4ef532e838e855701585afb9805e8a588b8c6dbe045c95dce2f8dbb27bacb60c8fd1448a595106147098a0f45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18424c9bccc582546faa06a28597173ba87f7284fcf4d37a4619807e13373204f92b0e85d5ccbb347784270e2d67768b74fbf37cfeacb7888ec50801b5362507133ba4b5ecc4e99c0e907b92968c2360613d23e94f12a4b4792f1bea2074cfc44b86ba608efd20f29a6e3561a3f796883fe973dd96e505517;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc0de7be96676d0f74b55c6654c8476e65221ac14ffc67fb567665aa7875e5a141e22329fff21c06a5353cf693aba7e7e216262893a62085cbdbc4b226d6c9ecaf0e78773281eaa085e7f5280cbc3dd8b2d23124c39ef6f68ae2fadc4a7bc77ddfea48d1bef099df7402e0cd06f84981bd6866e82fce52c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be80ee7b3005c9e5df11a63d4e9d9c3af925ac187c4b6d15e30819f21e28d2b1a698f2a9a47909e4bde5677d3e4149a1a37ec8fc35b5b9e351f3eefa88894c11c9fb0758e95824bcbb9e19641a40c430bf25bf0b71c64e8bf29bb67695910b3095f872bb02e419c7a84f8b2a51db6859b29a5aba94d79d18;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3e8816ffa37af5978f3a08483dc576647002af0516eef65559b7ba7f880be0964cda781eec995fac24182a227643c11536023c5fe72118dbd71d038a47b5e3f06aa787d802c5e462af8ac52d5fd7d006c1b54ade6299ec7c127460657b769e239fa75b8510409e103eb8ce15203479eefa0e21a267d3676;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107f00282d723f988eaca39262786ab529ba27e5e137c7a0d2e4dd103bb09ced4058a10d0f3a71493f7403570158059503ef67fdd4d8951b6c4c67a85eb802a6906033dabf1b63ee50126202d447dc20591d0ad893067dd2cc52ef1400eeb7cb473372d771f8192551644de12bfc98eb78cd9dfb9a5d47c22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b0ab1a2fd51715e7d1a470956295ac689fd3ed06afd6e18404eba1f922476546859b4383353206ed2f0904e1775162af3844424e41488373b801c2fdcc9bcde3e5a4522b5fa2b4c71ed1bc450e3177ebb32ca13776b12e894a8f0046b39abe8785f467450214d4c5f18855f837cca20ed5ea58e18e183db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc994e298f0c75c03d328590a242c5a7846c83bc0fb3bd1c4ea238a752c921bb19b0f4604b29e08161921f5af694474b8220449ea21f8fcf6fed4515b68906a71f19e74711b5c32a477a7fa74636f2ff00150b0de941f0fd37c3a062a442c44ca98f3c57903b9f3af9a672d93f6a3545bbfee28a72249ee5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64bf0e2d960b4b58d366ae1daab6544883fc22b8429886e28f72d092985fb5c77413a1bbdf38cfe2fbe07b34088c6cc9130be18c43cdc50e68eaa1a0783f59cbb15a1ce5a687504ce8e5239a8a90531e36899dad434a0de97178932637e7d53e86111ae452e33fc226fd5c338ef154e31ef76725ec2c795f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3874f59c006fbf2d2806a723a8f007b585db4f5def8da3be6bf6d3fa55bc9a96a3ebf4d1abf5ef143b2e02e17982b01a113ad42926642dc07ec255913aa5609be13daf4e65f2f5341b1efdfeefb9c724a11fba8ed815a3fa9e512b7e79b9d28bbae65e6922d98a71fc4bf937a4b4cc24602f2409c940f6b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b5da450d40e337a54462bb1444fd683e49515d30b2f13044e5c4063022a82679445a77cb7d249c880d2817c8a7cd333f374da3f058e2c5172a2ff9b975513b4c65e6a166e3c8617dfd13abb4072278ddbf9ce8e7bbf8b5199ddf21773521f4a8b43b809f97f4b959aec7b72bce9802b19d2beccef27e73c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81f135ef64e2cd6cd4c5f8e032c24e6103f1f913e3ab3267bacbd962304b8504962c9eb2ebb69ae71335fdaa36877d3cb81722cc5d3e2c527fdec97cfba61a9acac1fbd90377caa8804d283bfe534e87f97d9495d8b70d12f2d0d72b3a891329da7c4efdf5cd6bbf3890d3f37470c3b64ab04c19f34aebf6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40e04a903a5ec783834642453d55ffed376290c10be0910e603d886ddee025bc1caa7fc33adcd4d96f81ee8fffd42ce25a627292fbf157c23a43a6d618aefbdc47c429ac5bd1dbbf707e3b2775fd5d3131e6e6a47ba19c21191b50535958ef9220e74ebdc753a32362706e87066ab5bd1a992d4b7025227f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c3f78c9cf3ca6fb8ae7cc9741fa3859e14df59396d12c745e2ebf208b09732a4a02461854446c5fcf9473b4bd32b72e82eaaf462b1d37662828a4992cdd8ee82fbbde2a2e1a586064a482408ca76a9ad358a59b8413567d7a2a0a2eac187b147e3139f816e020e4dadadd706f2c7c0caed0ba718f91a4a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe7ac2d1c319ddb9a38ca8446f15a680b43fcf22a342fb4c7a7017bd585e944e32c60147d689892de3261b69b7108a2ab99dcf93a0e34f3842736fb2741ef37e161eb1ce2cd37ebb598aaf821ccdc4ab5249f017fa0c9246e5f50d4318e99a6b1de298b1a71d8c7fb4d9993f5ce9515b6c368da81fc8db58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a8d8a519a0d184e5ff22712ac7a306ad13be5bca7d580710c789b21a4d5741a8b90ecb97b6d2b77a4a146969b3c7e578e95365c0f93fd5a21eacb42a9983bbb015b89e15b6750b01b5ea060200a359453da16ad498eb31c836f93d03a47cf0a0c68aa7d753dee2534bdaa970a94ed04b1c16d0acf9a51c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1409f1baef8654b64f63ceb72d6666ac2b34d72fdd3f2240de310a4612fe796b1ae5b4c3d90df6d68c1c92e0304343201e5683eea6967a5a59e56b32a691a05fac5ca200d1489906f3768c2cde3eabba1ff535eb2bdbb1b950fe7e6d4444d1311190fa0216e4f538911fed7dc0c0a83c4bfb8f95ac7501d1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108c7492c7cd115bc2b4db8487e360e6ff8fc8a11f860a7457ca79529ce003209135075b418bb16c250fcd3f5286f058cb91770001be1a0b2c83965cf2fa02f1d2d2ff5548b01889c37f7054db5f6cbf4f58485c33ecd5cbd10937b4e5ae9b49d3eabae93e343d3579eb26380f2258b407b4c56fdea54d05b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he40c5abdfeaf205ed272ddba50917d83690f88fe049a5a6e447bab4e07363cd2bae4b4a209c9b3aa8e3ea6db86ba4e7002c27dabde0dba828c9fdf83b6e413b374fdf39371681c3262a34274f6bc99fc796bf36a4c9a083617cae40d3fce206b2bb492ea4e43d5a55747c95ffe5f5c771ac29dc2101e5f87;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3564e2d76f164ae4b36d5b6eed0f00c3630ed6f163eea88587b8b641b3aecab1b8c6a7b235d7bddf9a2e7e945f186d07ddb55c45a8c01f69549a9ab8207b4dfabfda7b1b4164873def79dace2893f8d8f391353c92aa4907c87283ca9b75637f8f2da3fe2dda6abc9be0c20bdb7e6a48367139eec03cdfbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae1fa9d95cddc16522a58c77d2f0ea1e671dc31fcb09b5c938a8478021b2251d2a3a6fee102ddc94c78cfdd004031de16b64992cfe8f0e89c8aaf9d42def1058d45524a0453136a27050f29ef1933ecd62532248c961e179de95f6742a48010d189a073a0af3fd7de02c41217ac9ea944e0a3b9384b086a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83610dd1d6b31c88bf78af9a75aafc8157d270e9eceea43a79cdf2187381f29db31718c0393387a327cf4ecaac2678bb57d5c45a870c93876375b64203d1791a3e366f7c3dfa670908f49be2767d8a8bd07b323d9d290752c0c2127b8545451d9c8f9b35b3f91e317190a30d6c4ce28fbf8180a4bdd9c2dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf8b1b5332c033c45472117b453e4a6b6b8af0cb75f13f5fa21f76c74fd0ea4eb2d32bf18b82674ed2e8eeef5ef1a8b67db267ad34376efa36c49c77f75b1240ce09f6ba56879ee610a8fb106cceea41fe8a8028180a1d72a1d294341563186330539d20a292e2c678f93ae51440fc3f428e1df0a82e0a26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ac25ea59f4f2079c492ddab224d216a74296139f58be314d02841676e2535bfe64dc265a943d5e5976c42dc03dc16c78a76cfc4f3bc2c90666cbac7f54bc08605edd2592636c5d6ad8773eac1777a46b709b4ef8af87a0cfd11dfab1ae2478954ec0a02e51d12492db114d1463b06999997eced9cb3d5a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5d7fdfc2ee29fb9567a7c4e0c6d89658bba654f24faa29ca0520c8050914621b7ee00865b4143b3487cb3d1b0388ceee43537b956a86558e82d70ea4698b71f3d4717f1e8fea8e77262491773a3570401813af9aa40c7264864a9aac3461a513b4013378446081291a10ae680ada5c6251e09d80234088d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h924e2a9a4f6953551617493f0b49b194b52261c5852bffa1981c97886eb1c6d55a1f85f632b81a10eb257c5cd0c8eae1f7cd77c1d909d75e8b4ef0cb1ebe471872c95c875b248fc8e65ee5e08cb958004c019c7f42b3bfe7814008868304bf482c6e9923902258ea682cd2f837dda7716982ef5df744a3b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edf45fc372cfd2a50c7d80fe644af19ae964b116b1695581694102f586ec37e61ec3f4c3ee8f532ce62a8b9c60b34aa5f9f162263081c3f587a4bd1526a73b5c54cb876b183b849fa5437727abc0306a31dee90f1eb1581d08426e2f07c6173a8431938597b31bcd16b24846ecc566adc4d9d16324f6f551;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8caf1883acbe96895de5b4a927c1fdb4f4cb8846379dfe54cd19c48b95665776518416e06971f570863441398f3a87bae773c046d8194a68293039e21baabacfe874997d3e6c535ea4979e23ae2d702963bf07ce41b8caff235093201c29b7b135a879aaf81257857b5ca5e71916e0bf52692c9421f3553c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf392bdca141915fc49c3b797eecf72f29b655d1ba3843ad415b578225d72cd30d4a9606a92a0e6f7fe8e8f4d046ef8b684c0a7c971084395934575ff133ba19fc846da431da4fa760565b835b60da31bb2a2081f504df86ca2a3bc8c7aa555a2a2c7be94d28c52a3e2c35945c219319029b84ca3904d0c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86ba3428ba70852fbc0059eb10b1a5a05158f568801a86d6e8609f086a4ca35cc99232a4942cbc93bda34a40a52e20ee92787b1bde253f16874951fb09ec789f37a4fcd2ccb5a72c0f92a0a133146ef9200aab2953c0485dd7cabb81eb4602c01f0ac4c15e8fcf1c3f396d4c71a02a7e4a5d14154445f351;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102446bc204be1db038cf470b89f1dc9f78705862841faa971556e0e79362b2739705cc9f5267c342e7f0a01ca1e8ff7f9ba75e238373a02cb692162180403dbb729b214c00d1cbde6519386a1502c7fac00a04990a06b67b3c154175d088fb4133f6ee430b006a77e62edfda2f23dd514fa79860444ed949;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2b1071d712bac406d74e32a4d8485d659e20a6123cc3011f96cbeaff7bd5f5996cddb1c3d4d69e0ae8df45833b78653b66a7bc4a32c3d6290cf283dfd775773a95eccbefe50f7c0106b4e643770c245454669e7ab5dcf4a99519d306d46a7f252e549bd7bb9fa2df3694fedde0224c1ba2e0a388cf6fb4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16339581a0f5986f31bc80d7028207416851fe455db2bca8ee17b7e30583175117320df9159dad7aa3937403a453a2fcc0e70198efa1485a8fd252ca8214d86a00756f8c1ce5d05eba24ef74a004ffb70b85bca5295d156d96abbc09cb4ab8b1425c68ed0dd8a19b6cf58fad8ca4c7c0b9aa6e70bc88bcd36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac052140cdf408d506747dbd7dea9afbb849cc56a4489e17f739f08830ae7c07f3352970faad450196a987feb7f1f8ee5229edcddd43d9067932737d450cf53770cb071945a3f9f93b7236844ac14648d2536adf61c2967fc7df135efe0fa32e178519f21867b33ad083ba8367fdc15b2138a458a150c968;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6ca4c2ec4adcbffddea1429600101b9d724ff708c0e558520d93eb9fdf1d4610aa654c1efb57775147e42dc4064f9d4fdd1bd5949791f46dcd688ffc99a6dbda420e2a990317138fb069fc0ec513f90e389a14d2e861e24142acf9091b5b4740e4b36addc7360ff50bbad544eb04adda81490da4afee4ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he28d82072c3b8b725a1196814c5b71c55e09ea71c1795ff5795aade40e851211e2b9d2e71b038020c2d3e509971867e2b322f68c3e859c8fc21b88eb91d189300ef887969c842f9f96aea74e8a4f800a89cc6b7e5fd64afa612b4b8cb47de0ec9851834a3b365188666cada658070d04b96b4c3fb246abbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6194806f712d38cd59f59dbf333015eced49a38bee039b7b61a51c7147ffda112e7e9ff2600c51e6f1c767c7f3fe892378473ad9649b7da658f1c67456dd4c53e69d54f66492b78768654672afdad3769e921e2d115e6e7b2d35d9e5015245e854d60df94b8e48a5817c59f608f2e4283177dbde4066f28;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1704ec386f12cc2c081c08fb92fa7ce54688d8786364a0e593e63ca3d6cdc76bdbab307c55e8afb29a5b0829c677676b7b730b7db3f7e6a9fa7469edd16a9717b19161b7cc40b3acc6b6da9caaf3983efdb0a83ea9ea77bc33a230109f0e3649184559cfdc2c28688bd44c6b90dc283a81f728122de733838;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d12fddf3c402c56e1581e3664bd68a411197b4c3e4e6c062821e0068ea4d53cf8fe985d74d1e572668b7d71eb3f7713aa1247de55c9a896060403b460db4c100d4f0a3b61fbcc827e5ebdf4b5d5329404fd12e3a8b059457ef2a1152b8fddcc4787e6eee22c5efd2ab9d775f03ec7993625d5e42ecb691a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f355673606c18e1d374b0c8e2857d657b015dfed74e52742c6b6129b49ecad7b1dc729660388b60f74979614410280229987a83490ef7b2869f241878f8053051c6de78cf401f3002b0026a060e07c1e69a6c225069baea73654f3fdd823b95341b32c75f14e5cf656832de154d90b1d202be0314054f9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ec7f89f844f0e8b725b5ffcd624691d8fbf402b6f87bd808b81069e4fbd45745530e511ae5ac88ece829e8de8c1479e3a485ede6feb6207b3476d35bd29d2f20f7b4968a20c29b0f23c1d7ed8b9a218ca9e04f3632f3594457213c68dbbddf32536dbd3221af1c6113962ec3134af8ddd4c71e7a291dcfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c82b7fbcb2380c7769296cfe09ab7f96cc0d51711417d712ef4637a223ede6a11db5ad85f4be7c9228fb4df133eb9365997cbe721c650e95ab27dcfaecb97ce06731989d0db72b39257e810bc3d52ce88585c07e02d2a997cae9e04f94e14dbf6a74ba74081ad97f34c480a3a25ba1e243e58c465297b75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b68d1cfa4a577dd0111465f0e2a05eda99ff5de4f3ef5e0fc7299131c0e5da553fa31780b1bad0a3708212b861e316412d1b38647b239fd379c667c79fd8f476dbdd4f2759a6ccc9a10c6da1e5dd591f473fae657178f07d266bbbf1046fbbff4ac448650d1b1bb8849f014df32bd54f2bce5b6252653e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12abe84a5e636e353c40437b8e9c8cb53b6fd267aa0304df98029ad938257ef80f592ea35edacb96b7db2d44bc3ba77bf178dbbdb50ef87379a154960a7649e5c3958fc88c18085a72f6454683a0b96b572c2d1270e889bc58d77952dd384db3762efd463099c9d91b5963969b7d026a89f4f289c15427bf2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2c63299c2e8f6b900938179baadb62008b34e01e8cdd7aa2e8bab7b0bc74865cab4d8b4e879d7bac12c275bcfc51a86060deff22322ba4000044eea19f64cc808ce0a3bd39e6597852ec90fe98ef44d5a5cb05b1a4e00a9ff8e292c00783243b4d8192b936c8ae492ec5850e455816a8b80a5999f8aadd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6634c3166be27f7afed8403b5f5c1597814a434da398bae0326b773dce300802ef1fae6a51f553f07a06c426b821c71514720cbb80db682b8f5f953d53675fbcaa0b269846065c8c366752254796bf5db019be94037107c281103e4407f06010a720ef0f065c23b8d1ccacfaa24b02751adf790a46f79db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35f4b6ba737f2cfe8f4362fd809e8672d4f46b49401a62e714ded9d069ebdd6a74f16a9f06be30f30de94efae93e475ef4b40cff3f4f7f58f9dadb719f4ae01642a204e1aea2b07b2df09e3db7a95e62f5d843871eb2a2dfc7b531fbaa121bc140bafa8bb5ab7aa11a623eebe6cbd5b713187c0934678d74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14bed0b85ac1d9a8e24e73fedad8783e9637025307ee189d9897da575f9e35a768bae41dfc002b172c7b6108f00e678ed7daadf4053da63408485c900ccfb6fa982e54f400084fa5cd584d455acba02d1efd3fdda397942f2f43af8b65c732a64889e3af27f10af7c2cace38e81da5fa9021107a8222067;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ace4efab42b949f4e24110e269bdd3acd60305277b725ca26cc9011ba6d94bf2fb840bff660d2de48aaeadcffc6db530a85e8f20681033ffd0d6ada44a8778332adee71ad3fa554729763bf3aa362e925d9f4276916bdc85bffcb6badbb4ba20bb3ad711c3c3340c93f93352c4cd6182e744c80db186eb2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1d7db8473dff4736e83f7f4738d6b49c11ec20d1c74e9b4a70a3dab9e85828b68c2fda4d26b614245f3c0d831f44a0bab679e2251a7519e98c54617ec2c8f24047a2fef6aa2f912ac39b64066f552c6b47d08c18bcc28e722ecb4b678d26871388096683e70cb52682c9cb0d4aad46f020e529092301971;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac813c4cfeb4038d5659198d8cc7340ae5ec0065bd608c83a009c328dbcd956f42fbcaed6c4b957a5e832c08e0cd9cb46c86a6a3b59b6519c4cab31de8463296f96820f7725687ccbe895ffab0fb81cd0db503294a0d8368698289d861c4d1744d91df350862fab0461d938520c134d4fa8be9a40ebb48f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e39fcb5be527c8400469d5708204ada19cafdd3f4582efeeb2ab2eb5e4c588fc840b5c06d409b52ca29b3449cf144dbae9657511c3760d8303761650d20e4c74a50e4fa20a8ed1823a34aaff7e5d622e3bc4574ca98a5ebd1b8cc3fbb04fa63d3ab846ef94e8611d4ecce48391c0a5ab721bab38db76bf32;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22b72e453225608e093ece6998f1015b1af7d47133ddcbc43fe091eac8ecd1f90251e1f5c5c0787e377d20c8b71b3f8b8f6da8cad34cb775a74ec0e09064b71b11f418b59e7496b46070ac57918cb547546f8de7bc2dc381156703c16de5dbd7c245d966922573a0ce15556b7939e39c994946a49f91efc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173416595aab5b5bafc56f1c003c2709605198e54d21b4d47b8123d69cbaa035e65ee7a9b753f184c409ef761fa96a786962de743601166a0f092c059e3afcbc0b711590fe5e1068968b4ef84e434e6479ba09034d45e84696301db0c314bc4708d3a8c137af443f22dbbc4d10d440242273a9e3a44b660a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10be15119e5a27b9b3b053fb9e5470fcb119354af665727bf427acbd9c34af818bfde5fbff00b3fb1934328bb078a7e0c82ea03568d10c1209687afdcf8ae706f2b953dfa31ee15ac8b2f508fd75209fe7e7dddb362aa1f46f3cf005fd22160c2aba42d8a68c6f2351fd7cd1eb73e933541a00034e6ef2a0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8045ff817f04296ad5b8f90086ac38c60bf95e64e08f8536e4495977b4610d97547fd9b26d8e0b14b32df6561b5effa3a6ac687e29f30d8c262dbfca735c249fdcb1fce139bb49a68265ad95428e56fb637967a63f18fb98917e9c38ef6ed6834363836634984c9efa205f2459dbe35958e10a098b6a765;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f40255127d18b8ed4230ce6c30d93c8347425e6427a0312f603b503e927f96ed39ee17d8101720c2a4706bbde64aca962f2cce0e7b1e523ad849eb13e748b6990d3cac715a95eabd9a8b47605a0454a67f7693960e7e57aa0916aa2b353dc6b38ee92aa5ee7ca711d5cb41b87e0abdf307ee64251dcbb066;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ea9dfe3bb9f805e89145361f3ca7d9208c906c906ff9c4518e4a9dac358120cd52cd3a63337667baba16c785926aa4e47fda83f15fdc3285c27a783a58e7108ff30936ac80e1f323c9b21fedcd7377c5fdc71c541891e20491209d000897282b2de92df425b12c726650ec75c7e24e212b66e0ec7e09c45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6f6e71376766d1f4087e7e4a091f6d078eafc345ad19cb825a70f3759620a965e636ab90a338f1581a994f27a8bd6a729e0d7d0c8190e06887e198259dcd9cbe8e30b18ac80f3d585f18fc8292e04188024a3e94e4ff565e99ba667709d0030e2cdb27d3adb73b9000e4c6510f63d660b6742c42be93e5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bf56d99200d8dcf8fbf7bc1c82e7082b5f816dba971af9dbf090aa3237a20c6b32e9564c06fc236466e7f816288b760dfbac85115de2acb8414d9b010e9d39707ad127e4661973f73b2e456f598cd1b63ae01c55d7167b24ad9c4823c5e3368df8713b00aade691bf1f27f459e45489a75aa927827eece9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1321691ccf751ac90abffcdf873eaab2b76d3f1d1e48f4b83145d6026793771828c5e0f300177f7b04fa83ef7f80cef0e1e75e8fb17b65c7d7eae755a1e254b61607deddd76ab4fc9c186756dba12a5b51090c947725c60e53725a1b1b2f5108cedeacaabfd0513e3a5d80c865b254622ad364b89b429f7f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10987408ccabeebbc3cd110aa63da277ecaab6da6b8ff4face62fa8059fec00a26986a06f831a11b6148d5a4222c3c278fd8723af8812bc6b49ef7f541ba7dfa1c140123082926ee9eb39c2d32fc1e228fd25cd9b8bf5e60c55d4dad73df4ffd19465640acb1d6ffc521139123fc747b61865af3cab04052c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144aa5a1c85df53e90f5c5c33878656794d8d2cc00bb80ef0f7ee476c71704022808074f69a327fe6241335db30c32d5659fd54264bbb65e4b8af6efbd541412cb5f81ccd4439fe5ac24b43b6455bc29080c4d2137b67d268228bfac0af17edbab44c58ccd720afa4897f9353babed19d180b0d18b6ecb0bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f20a040c4cd3ffd97c2c4eb797d9c475e2e70d33c03244519a795a1f1e6d4646420a94aa3430fcd18eeb8dc99f53b3c04ec80c209d6018e9f0d2e85e02f66996b154b5a5cb1b4d17d3046fa7c26d23cf4ad953b6428076319ebdb3d2d2c7b3353e09dbf0bb2c6d53096af185911dd8ce3d117ea1c27d3e55;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14c2f6e1e394b35cd4e18d1d44c37e6c1e6d56cf3092a924c6b48667d05973e2f4f7c8ecd2560caff8e7fb870287164d292bfbfd76f4cc1adc4bdd6f66b4383039eb60a2f1398d45ff3cd5179a0ebb24ea944b5fe79316e309194014eb26134df12fe38a1564601a7b8384c415144923d465788378a84cd1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129dacb9cdbce9f9e47d6d140ac76872ce58d3eb99e386d57aaadec79ac8231b915ce1eaa477fd4703574b39ef7faaeb7908c6722f3c58c110d9fdbc6315827909d4f2d266695b35130ce36c18e66960f1e601eea964e709323cb9ac19777e56fb5e5bfc49755cebbfd8450d1db5366903348800f21c12c96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f22a0537fbe83674faf36cc471d2a176a18d73adcf8a78626981cce152c6925b688f1ee5040f9e5c006548165139ecba47ca2a1610c424a41bb92c5535f7b7825eece811995f505fc38465d491a780401dbb9743cc552552f59b62f760b691ff10e51291b90a4318d0c68f0c3937c57dd0722e45879344d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4c8481b3fab53df71ce80b7df2a15c3d5fce2b30a9853b7b19e26c6ddd9f9fe7650c8ae1978355547d8f0fb99b1aa97ad80fbfe81fd77e82540c61472623877e1cb81e7f26dda4aa788e3b3a2ff1927e72f091c99adeb3f66691886ce8f911ed9b6713637e5afd10bb756cb1a2c4043fd830049cab376f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53057c86331851de7d1d89c49cccf9a57893d1b40c3348a7e897cc261c52e41e5d5c824ca77dcdd1a90f8d52a9c728fac41c67a04fed45acbfbe8af61b97c0ca8970081c8f398578c57c3e2d6d9621540f7ecfe5043cc393286de2777147785e3dc2a4966c6f813c097a420be2009795cb210f1cc5a50288;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4daec4a4a17c24261e5f52374042666ade2a6da8ca41470d1053fc56c2134c0aff262ab557af8d7e85427b150b27636bed446d266d7ff9b073f87015511b4597b5f2ca8311935dec44c509f1530f5de88d4116b1d9257f6e47b6e4e40666d5649033bab3729f6c2fd947651b2b3aa1f5a8ba60f78821d98c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168f7f960b7fdb56ed26a96b68af007aa45fc79117f0ca593010d40812cf8b2e2597dc48fe86d7ce563065318203943d32db96289c6de34425dd2acdb14ad11f7da0fc74322ae916405802086012f762aef9a2e23b1b53c4526f92b0c99b78eafbb8ed9c30043da2f4042834225bf8949aae3f756e242e160;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4065058a7a27edbcabe4ba1ff34fea3b412d323d8ddf1747be323d348e1c490ab99c269c3f05e12aae6b6e89ad3ccee9c01ed8eadaadd5cf6863ad20900599a1eccab1c2c8dce18a06c07558b0754cdaf1e388160d00bb2f5bcf34bcc2895e169f52cadd2b40614d277daffb969b811ae155d0767af17f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1acf7a8c4f5f8acf4d0e09290df4924acd39bdfb99ef06ff1ba0fab7a2fc8bc219617381e000206512b19a806ede7eebea440f74e35e9df42c0761bc46ae4f45b455cc558d033f2dba883148fe52f8f38cb14b36a9bac93ce9cd46b449e3fed4309dacacf05e621497642e402ca1f68370b3838c8864aa2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec11e40fd3a02c9cbc32059013bad532954dd7db92977263ac64ed75317e5e94d4a10f5687fdf0d442fd320bb3039ab3100fdea85915789413bbf8aff10edffa9db43f91dbfe5c2374b0e53cad9370943b28aee23f10a5ae990a36242fac8cfe617f2e43077226e59ad6ab8e0490532161d037481a2f9d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe5eacc5e4b7831b6239b9f5c8d674f90a4268b18d8108516e38d70d8dab6d7897d4a76a97f2e448bdb4df23e5509fcdf8808a7bd9c3b4f42e7b8ea68d9e70c27d26ced69ca393aa86e9640e02db36dd06d383fbf87c8d0d9a277a59e5fe6f72ccdadcafdc992162d7ef42a19cea7c5928db3a94da37b569;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b567b6c49d8f3f2b361820a91e680fb17dcf87a30e8fd8f07fb86ebbfb92ddc2324a580c4f1ba268e9a3da4d1c5ee62e1e80849a01b9190500783619fe65d29dbb7286744661b53dc64b629500598a37821b9ffdb3d6eeee838e6b508051c7dd4506fd29ad68d49036c1f623acad5e9f9edae0ac0cf5d40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7670476ecc68bdb8c3ceff653df323fbfc36a3d2c6840a267fbf112a64c0f5fe12843af8479175567f628fa511194c402bcee598479428a31cac401cecaf6090efcff086efc7e7a46cce98aad394eb674a7eabfd7f4ce9f06952b1bf323b9da10fc97ae3701754122486a24932e044be9f21352405d487be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f02680cfa9f1bf6e2f4b4ba48f79e3133356db9154c78bb1e7ef0ce5f0fc1c0ec7d2a6723ac1c13ae68373ef1886cf57f9a5ca8b04c7f3eab8ceee800614d656bb25cee1ca336d65457b4b00b3a6c1cf48edd86d96cd691276105c587fb263d9f0cb814fdfb03bceed3a36894a8de1fdae68bd8b2678ba9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59aba54a9e1e4efc73c763e3601458ca1046275f59f4ef81a4db423a67a4b5c9a397482a5dd82ffe4ea051be66ad9aced99bb6aeac4f22194aaac697d4671ffc0873a4447dfd58b7d77464c12d25c94c8abf871e9a1fb2032fcffcc81add8ba0b3b5537c6c369549629aaf553667d887b462e6e902d93dec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33585b84fc0726b748cb750cd506e7210925d4e2045f3c40a1f6c2e8d07d61dddb44e6f8022af3719063d1b0cb7921d756e3ab0852ff12fcfd8498bbfaead37047f1da69f2143156a3c95194088c80107ba3965ed0aa7203ac3406c792dfdf869504e382e77c70529e5801d831496bc043dcd4158523e8f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143922cbb0171fca53ccd7e10f5707393d8d2a1993b376e32936a825bc5bdc6735802c3bec8a274469be70df5cbe9a84b6b618dafd62b7f2dbf519992777771fa777b82aaeb3c6b6614e4a0596a77719519732e9abb5a78a2fe051d4e37080bdf19fca67566bd30c3105f36a586d7216db71c975e678b6e36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10893e0280b32443660f504e55b9b666c05760105f7b8179fc0a3a0ed794e455b8c8576c9904ca872b41fe4128f324e2b73c7684eab9e929ac97382e067e1e161c5a1820954c4f02ff94fb9b4f80f8e1972a2d902124a5bcc3d8cd1ce253e170c67e851c5f103a25e9d59ead7eef937a7279feb38b6665517;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58cccf1083d9869aec4f634702d5b0877ede3849bd0983c8c0a269e2e8e920745551b2c72b9f0e702072d3476c7fd9faedfe56bb2626fbcc9738bbab805f3f6a04abaabc2cb79c837cfacaa2fe3c770018ae1d0cc0cc724b811920bd5b2f07966b8fb8feea066a73e1700e68577123ff1acc62bb8b78e0e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf02c394c1089e909aa43a005d365bef405e388da7d5de782628312dd95fd57a91c850896015e27a7cea3078983da69cc533ac50accdfb8de5b68e9226183bf8cb12d30e7d0391fcecb070c9dfd9b775e43dd7dbbd7d730342ce207484a6654e1fc9426da4100a4ee57c8106d34649e650c6d583ee060aa1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9580e9ff089347fed1ed19aa694b3f0d0cf467b35beadbfe0ef51396814682a3ec5ea3dc82c76645b18bd24fbca2c331c4da459150f2b09acbb1af3bc0093fa8854abd1a8b0f1d72d1c598d0555967b1eb8c0b9ba86536512968763d9c06b7a2e1d8835cf2b3516a95738b66262e27f2757a35907e67b75e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e5c4dac96387cf994a3b4428715e74e099c1b1b0590ed6c7023c54e8aef65220b5bda77e30084016b5bf4b9868dc7be6cc83981c0ff1cf65628f45888e85e0850df0770d160e00018099c2a77939d83565172da7e7978814c1a4d090453977fc40a4d461dc3e2ef1079d0815f0555863665cbfec4ce730a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0480739c8e3cda87780c34894ce4b4b64fd5376c908c7b48971837d3a10de0712a8edf1b0f37e3019ecf8170dbda4aff600057001c227da3624b6e6a0f55b7d9543e83e835ac6221b82a68711b36027e6f117955588ef869a4eb590d62c9dee98203b20ff78f7deb3bfdcd18ffa30698d9d6d2fc6f925a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c3d6dd4c13fab756fd74fb5c7bb65691c41063a9b32430f2af5ca9c58acefa9f2191c5b735069d275537ac8814cd9ef2bf744c40b28e98e21a6b84032998671e1c7efa6365d9946341e470b9f5a8712b3814e6a4a33b323b70baf8b2cf205ff3a5e96c88cb82b3a1d2166e82cd88dc83dc63180f4a872d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4a8a1c64a5fc108de24a3fd27b20b80562105c6b0a1056695543810f71fd8be47d6a1d479f15842c456b926e9ceb58b8caa836c662726ef1e21a9075732a1db2b234a232e73abdecee69f2770ba033de241ca3044d618cb976b76bfbe3470b8d02ab48c619cc4855febff479127304d53617c6332c67acc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf84147fc9fc64f0acb7699241b146967ca9441d984bc767185e479ae3164ad7f7d41f5b23d01551ba947d575b9fdd272612c7210678cc23b41d1621331bf39355bf1cd2248d8544042a3851e16ad4aa7244a26b9c3f5f1e36657dd84de9bc28a31680c86a4ca28836bdf511f4f689e8bdcc6361672bb95a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45d1b6288cc5800f09c18220b67048759f89efbea6fad27ad0c1c58d4a594ab15d37672a8e0ee290c360bc91d15224e5392d1a60d30b073671df66ceea797efb60ac18f4120f40b41e85a952bd31491555269a91a51143a710ca1915682aaa561d796c022e3c2c08c24100269985f2f3d42eb62212a26691;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc95f55ff83d3e2954fdbef65e4c3b0ed62a4def8d33267caaca680ccfe99422568855e3f68e8ab38c24b94188d4d31a4fb732c49948dc4b6f2c5122a770e91adbfed95c572e86bc863a981aafe2b83b81bbe54adc7112d1ce402df4c0712053031057084963427dddfbb8ce530629adbacd6cfbc8ba7871;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ecc177dc02f27339f578bd67164ec3af79c4786fa9a3114289e9c1dba1904b27a6d9e8ad2d9af7b15b793f1eb597cdaffdfed98f24039adc788f16660dee4655fd653d66ac8471d19713800ce5c9a321910d810176bb06340aff0b92ab672ca74c8596f7b1fec54c5321e5ee75bbb9a223501cbbc278878;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h158f85576e41e5dcc958087380da7b2c2c977099a5be46221817555f3804be734c188d68259c835d175a4b10a8368baaf71365aed82c998cdb00d269805b2912e767219ee0e2591f0ce56efbe6224475b23003cb86fb9f4f37465127e5b8bdd8e7598674358e8bc8c4267953e4bf7b94a748bcef6aedeb247;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b8ceb60ce821872b84ae9f65e2e4a1a1d3acba744ecf677e071d975bca0bdd8a2517c3a9960df2f743b4b7ff4abe3dea9b8a4e59c8940b4a2c648f9a30ff68b3376b2b1b8b5d3d63761ef8c59d81fd846b092ff58a11f08a695e2c55bf737502e6dbd9b683686065f5e253a8f6717e9fda2c5c21c8af5dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e909e86454b64b4a9ef97181a7c14eb98e96195fbb5537cc5a239f77932a31e985293ac7e7d2f4a78889bb9122f2db9040dba61505c234375909850636c16a9ff3e6e0f48ce5b120b2552451c3c574637110c3f8ac22438f36f6ac640400136cc9745546e336db4a4197624e0781ff70a82f98c54378a63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a823998aa98ce118635a3565eb0c65562a08e1f17def7e9104bee9c4ef7748096a18f7d836d22dd720d0c81824b321a9f7a976425e4975718cc7428f496c15758d88637632fd963a4eff6730a76f7d64334b8f811f9bd5defb53d60307e9481c1fbc47f5d24f67dbf075645cac972cf72436d7014bae0ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2726db90dca81931645829b420f1c36a7edbca029ece7a85dc455003887d361f0ea01abdf02b8b3daca937b1591050367ab6b3541697641285c19d1aa854c3d37c7f3439ffa51f18eaa307445453da257bc8844f3c359d5b74ed2422665c3e4031f23a9017fcf8e6a5153acb3856129abdcc95201391a61;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25cb65b2f500c6a43712ff8a282abd61f025439f3cdc7a3907b93a8cdfd9bf72c5e6ded261e946ec887c9523cf6ce34392bcc1b55792190ed96d3201cf550fa91795fe5c733df9d1ae9d8b46dc7f82e90d4c133b6dd8db234918cedf5eca2ccd5bf9e336ac005a68eeefaa7b634e0762af5892cfbb9e6e3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb3e69348ba42bd9730932e0d247cadce5b5918dd85c421c70aca86adf8fcae344ff7eb60004ac23a224495bad82ef82e0ef416ab867d611e9e670ef69720fba461f87f1748003aa4b8d89d9997a9a6d34d7e627a421e29e42e7a60da9681d5a2da1c11116986f8cb99c146c4879c8f8386b799888b4a045;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5a6caa422a8dd421c0f894047395ab931f14575275fd1e312f263a317e4dbe0a2bfff012d716e5dc5714eeaf28a68fc7f81a9d0b2e91d14dce6a5e6f0b7c76ba1c2a422c86682cbb3fed633ac926a79a3cc46e6951b770d7b99618ee185392b54941cff20239d39acd4bc57265e6b9b82b902530dbdb76d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d626d8ef6947856de65340fbc7a34bfb725d1a9efbe52d10dda0e48af7dd54a1e7f538b1a17d4df07e21ae4bfb723b8a55062184a79f1315df0589120f8f066e73c6bc567eb61d5f53b3bd6b3bf51b11bf10cdd159fb6533c653795261b3726c05ad88f475745656ffca65d48297cd0316c15b0c5834303;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d13fcc116e57bb535f51c432179b01f6b23e531a77034d1d4fba9be2cfd29ae29558884dfdd49c7bd0598caf19a0df4e01b0f3b53da4d28ace527d4a8e051d493d96ac9e137df460d81fb620be4f89ea62d9f1f23efeaa438a2d407f03cebce868b2cfa67294b4731e309cc69f3c1d2ac3def448169bafb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69b62098f1c376121cbafb72e4494aa3a5dabdafaac742dd152b6155eafd457763698c7840146110d7593cf694a19c412ae9c0bf0f6a641953c06e1486366d3c943910513c4cbbe8c53cff7a3f8e9ea6ac461ef74f33902a35b776f76e90e3b4892249aba2217beac1389c537a77921a308c161a732f4f30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c69b6bf1f03ea887e90417f2f22b5e9b1f09442209fedb6bb35f7b64480534cff0bade0e8a8bdefbf0b77c6f31fe7bec0b1947e115e1936b6eb390786b722b6208c6ca66f609c48ce5237ad68e0ca3ef5bc8f60c56bd83fbca1e9be3d8f30b2f864dece14e6e460e6a1212cd2338034d55c3103a3dd867f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50596139b3016211cd2567a82efeb0c14b43392bf0717fdacdc0e3768910fa3387887e3fcf2ee88cbcbae902bcc4c0383d2df10a1b053e8c865017f035ca6f4f4077d2154f5a7ff5ce9ac1a26a5b367f3084294a81169ec2f3f06bc75c6add041dadbab67d617b20d8bfb19548e456825e4d5b41ae7dc2a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74251f2d6964d0765501ef09785413302248a30531c633278fa7abb7f1d5d012a445e838c7896bba86b81d958a06678580dcf2c266eb09ac364fb12c8795dea24240857bdfb759efb31711141eb3eceabb37854f2506ba3d967181d77cf5c1825a3e75869b731f8e0edf276cc41aa50ee61b12d1ecdc65d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd4fbd0552107074c6dbd4caf967064a641e06e0de931aedfebd313cccf594474c67bd2f17aecf0f1aa3d369ea13857e21431ad21b97bd4719372d612ed9576c4da348120f6922c76c336b42b59f2960281402b8d6ed2e462f6c3fadd57707c60d967dd399626fdbbc0cc51ee8810ba367defee618a5f276;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9219748a926070a995e077e6fba6e1c4c9107102b991f9529a5c4c52611c4b83180b336ff84a8d411f06e0d7cc1bc890cf8e5bb603ed02c7b85b866d301c53075ec9b2e47d784f8a3afc9ad017b4649142f29c21fffd5dfc046ed25a69bc29b7e8e1613f49f657659365cb5482799718bf7bac3d12abcc70;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25448bc692feff6972005ae176225cf2d2496a6aaa8cd938a5ecfdf31f9662c135f8df4cb02bca0d61251339099ee3fad8a3f9b2891acaf24a058afec0c0cf18dc9b88e20f4270539155e2b1e614df03a8def2bb14deb53777cb2f8c8115182085c53d7da063e1acda4b2ec2a446f49f7315e64cc6b00099;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ac441eb2c5dfabeb42d515e3e32c5d15061dbeaf7bf3921e7cb3955d2971219843abab6542604738ca64209b527c8e5e417e0dc699f70b33cb26aecc36a5ad79230602f2d3c8d2300c7be913ce6db63e6ee2a8d1f173466f68abd14443d83cbbdc6f2307c576450712dd213fc13225a017fabe7e629a223;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104f9527643c87631f1918883b4d7488144c1b5e70a14b337e83b58ed338e1ed054719ba7c6cf6d8ac49929ce15800c7249994fb834e308f67de4f93bf94408e0eb9975d8cef793ff3acab5bc215473f6743eb2331a9a2bca626ea452fd9e10371430b14187eeabe62b102edce28649f73fecebd3a0be1554;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed5de265fa4c301ce1608c8aa770822b8bc0c6b549ac0113eb78fb65585368173516c02549c36d067388f8b25c5f3e06885ab9e7af162c23f1245f1dc6a8d080d071a90676f50e1831f165448bcf732fcad82690ee345fc43ae7ac46ccf2b095f67a33f2e63403ca945605b38a7ddf80142e3c1497ea51a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15866df06a745ff0985961fec338fb6f994fd13ef7dae0de51a4264dbac7a955d720568dec4b02ab6fed70e357a82a9c36e40234be9f3c2e638d24930f94ba87c03a9626cc208002f3381cd38c1d4b40e41d2f0b535bb8aff73807cbaeb4bdc5790cf53c74e4a76b6ea1fe4d8e734f83df744de4b9e510124;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bebf040ad4cda7f71e6fcc4df1884068e4a42abda365f58d0aded4e0c5f542ba0466673a2e23708a15a4098a3045fde70f2f0a54841a87e4e305f588f27f4e6d93b9a93ebfdae620bede43647885106f3d8d41cdc5146ccb6b2940f23ad76b06c1219fbf9ea855221b66d8201ddd1b99663afcd24495efb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e64978a588b95b5bbeb08c0dabba7e09bb7b604c26c037c76fc3f0e1f15ac234aff5ba5d7472eb21467e262d2601d3aa40212c85c85b605cc731fcbdf408b88871e55d535310ba2dd6eb264d151a709161b8fbffffddabec3823902b4f64cde84f3791e45a6176061038b25db99b24c6f54704ebd758429;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1832e7e0064342017647ec8c599bd256f713265a2b2aa4554933cd5b039f72f0545631be2a823daa795ff699bf8dc89e1cf4e1f4f7a0d5a56fbe4525df18619c7d06b65d6eb347293200035a189a2b4d4e150f51ff9eb73f3257da7dab8aa174d823ef9eb6aaeb4be30f36da365a68aba5501054ab1bcee3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a025740948f92627e193e65b385ca04d105b196603974c5084fd1fcb25c9837ff0565eb01385295b74cb48a2e83cb441c4151efb89d3e085ae66a9a36b8ad6618d968bb09c863a86b1151f61a635ddcf4530368a2171c3b5070f6b4d6241fc0cad5058a2158bf6efaf0c221d0f05d8e8e540cf4138505aea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad2245507bd519c95a4f5c1117549b996908db3dda2cd71b53ea954e9b8b847442276e0ff0c07dbe1eb4b610a8156669e4313a6602332cb58c833cb57eedd7641e710fcd22239a4862d503218fde6dfeba5a615771c2cc651bb563f0713794429ee227e11d1f7def3c3dcd6cb9d14f30da3a5866a1b68703;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37ddc75bb74d41ed79fa1f3704b271b5f1dc197f4fbf87dac1485c08865326d3361c3fc963284d9aa8c995f72d3730d2f7e9ef9b94a2a06cae3cf526f1705fa4d36bbbe90f1d413a130780b0b0731c2ee0d8406cbdaca7f16ec35b136c8c00086e26aa1e4424b4db05cb97e9d7938c0f1bf1789a051bf2f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efdaaf1333faeca1089210bab4e73f5859af5a4fb39079d9d3667c3aa6af42c9d160091af8dd41865b512d93cb884f1c819b222e5f9c83f1beb2f1b54449a5719e5eec5fc2b39135c82d05307c44036a2cb28166707b3e08d2450444ed42ab4cb1cf60906bd363fa683cc07ba741c8938aeea5b087f49e0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c7f20def1397a8c90769842ff9c8401c3b27d267c4a1a0e135c97306af81060dc5a68a685a1c4e81411ad12397af76c08701d209da62504db41c7470835539c582cf527438eaf40f9be90bd4b04ae380121fef726743a0fc266aaaee6db46011de1769ad06a16d0ceeb5544b959597cc2fb9c1a164bcdfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46be162174867144190f125bb3c7200447ccb2154ce8905bb4fc1e8bb80756ccec3e13db7a365693ae902fe35c9bb1dfebf6d3ea54f26e7d474574c0c5637823b300dc2d63f7f73332b6568ef6a966518e72fcbca7496249a56c2362a2db10161d62d0a9ef5ed6af29bd7123c98c3d1a7876aeb1a8ed8646;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3b668f0e7051f98e2da5fea0d4e96b8683f29c0056eb420d7104c9422102426a16ead05d5a4a7c06ad86add26db5f23bf3266d82778721dddf9f44776c17ae9ad078fda4bea0f4465c99879d9de75909ec92f87daaf771b24657af9e53d80937a8981c5cfd9c65def679e672296b278f7e2e25feb14ad10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89a85c497ca599e95363a6d108be5e73d9c8fcc9ee42b2ff144672db4b5f9c6a1b62ae389e6faf667fd39b1e85a6bc85a5df67e6895e440314cfe8d12e886d110249cb2c30f3e491d8c8b2d543d474ba05e1f52806683adb5dc9b9c4e9e3edd9bab74cdc7c996408edd38e810ce3f8a6173fd9983fe7c087;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1936c55be7b290e01c649af9df18d9b82d18b33207a86ef568ae526f699460b049023f0ede06bccf2a52fce754649cc96db47b83223c21a258c7b25d4887d13ba149f35bcc7379da90698c95d1c1c0258f96791356fdd1b566d39153277e5254b145b453a1ddf6897658272285d3cafe5ac4e230cfe0fbb83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3e71b7a06c2d326512aeb8c177d902c43ea744b5391fa21c878909b92687dc3af03eac3cb0a26147a1a9948361c985ac79616ee5868c38c8fe27e0d6780214bd4a291a1e9a76e43a4bf29ac296091076e65e4020a63fcc3fdf9aae58a2322bfcc69f23eeb11f3ce322ac4175ace42b51f9f1564f0322af4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h322d8551891b037eadfa1c9ebf1bb8469bef898e6774e86691c609f948ecee1ee349fb740149689813461219a0c36460d4d8b8c47777a53e37dfb82cbcc5ed7369567095f8920938801a7b67d82a77d15b4cd7f9c03eb855f5adc8a0feb046050c48881473b675eaa0135bc485c8cb2357ecaa9f9ac6c49f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193a00f464a54fec4e73f8119d9366e84ce0e5cc6d4155fdccd029076ab2b03ec0779a5bd2860d05fa3f0c310fe33907e8281246b6ad303d57e83d64f051deb6fe94f58f2ddc52eb74645f04b5fecdce0f41eff91985a0ece09ea79f760da3f1237e9dd87620256694a5531527d0601eb44e92913e273d7f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6250ad88680999c1dda40825be65bb1f1a9fc1746c4051b7cb02121c8b8fe585d6ad7f0f69ee7efa2db072ad6f58d2820dfe0bf282c3bde33f426743eab7a8b44b94adfa47241dee77b976d91a1b2f853a5fbc2a95fbdd30dd06093377bdf352a351b325848bcb111575b958ebf0ffe337854a66fd3e0c7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ef905001a3b9efd24fdcea3a0a6eaca9e93389b90ad691a095fc35baffccda01da3e1f8cc93d07c495c0a11369bc71c1494a5436279f9cac00994c80a6aeea30c59db493b61755ee209d619e2b26aae616af29d8893bcfc014df4d98e70b1d387a1609df4007f3eafe8d73c60f1ccb05d19f73203ea2c11;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f352f8b743b757887c7d4647e0be9a8ab1a24092be85fa51a01e76d3e56ea3b9615d9b3a3a1d7fa7088fd5c9f32b5a45b5790b0d24f89d6ac85e61691a9a1f3e36402facf6b8de823135a37a3c568d2a853bd0db77a128f65875be50a8b8c54e432d32fe2b0752cb39cbe87a12a20827efb4fc5431e855db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8cde0ae3d28b0d8bf668ccffb1ea2350bd93c656dbe42e2ff863cb07a99c4e87f0bc3109adf901497234d0a3e959eafdb88e6ba013892426b741766d6177865fef17622f3383067ef435a27720668f05e10ea3ddb6eaf2fe226e00b5573179ff4556100db38ea26341fd421d7a4ec1eba7434fd9039fc7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ebf8a997440adf104ce33c25130c9a959138af6d598977ec80119c7df0d756f23a2a50c2df7c85b89c9873e476cc44fb5113b3f044a53f09d74f2a4c6d5519ff00b277000dd54578776806b917a50d67f5a45b8ff7a9ca24fc7a32e0fa17d70745b33729a994472b51a5dc8505d72b00049269b77f27da3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a5774f67b9e9cd3a6d97c4537602094a090313aece6385d57cda9326feef6bc874a7ddb74a9e705d1f6c3e754a6ae507de1c7e550ce60ac833f9f6c0331697f6b4a9d61e3ad6c88a510c961b4f0190df99b54b73afa7250db0bee0ca408354bc54d30c601f318fca5396e692338470491a8492a97cbf652;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37be097ed5af0ce2244d679220e771d8ee827a767609f4494329922d5b3912d2b93b8d0eaad561a762e9a907000071711b94356ef87bef1907ee0d83130e2e1aa8a5871b5daa949a73447a01d970e8f5107566a1501509f96da974adbbf84693e618cb7e55c2546bc3f4107cb2982e5c4e1f9a4c6d5b0f02;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1855966baaed6d2805c2b6cdfba0f4ba2e804d9e317c459f83cb6846a22c53eec53670255c9dc50901e1888b9ac8be43679dee473b6357585fb215df57a1a5ecfa2975138ca873a523f69ea1a5f3d1e954a4da9907ff0b2c9f158d9f44cf03d64ec6d72dfc0c6aa31a89525e308965b5593816804b40ecc2c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c128642319e42b367162c3777288cb513640668a9590c7b9f3e1179c38b69b379e7ed3bf0110583cd1d231dfa2c744dd49595c8b1b6dbd2593d38827f6b5ff21339a042f6b71203718e49ea0b01e54f1e0c83b64c58a1165d7b1df7837f1a65afe8c3c2381ce1cead8c34807d4d423ab7038dc7f0b4a368b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe3cd3257f9fae9face5aa74caf9beb5b6bbff52e89d27611666dcba4439f9c6c7d98ef3fff62d95d473205bfbaea9898a4bcc729c1e5db07340c7ac886bc88dabc25d22387bd3b37fe10b2b2e1d39c94ba2aedbd689471225afd30c34aa7e27afefb52b54b90d336b4a34de6bcd752e4fdffa48c2b8810d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h308b7b70ac45dcf4a4aadf38b5a53636487b972306fe19da0faa0dfb6502a74ae1c628ed42e614632175430d95564f4f521820e280719fbc69adc2b6fc053bea8cd38e322b55fb9e0f8f2721389b76be2cc90f5405eb1895c9409d118e40281f45159016693cec9d06f68dcc63e6ca56045a7ff516d8c889;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e31cacc3b2e5c757eee018f1b8e14cf09739f1939dc4155da5a6aa2ebda74d3dfd33eb49721230cc7e5902d6edf762ae903a9c2a6026da4231581dfb3c3b6ca1f749b52b4bb2660b5085361ef9a8988424d197613649c52874f5a90993a97ee1272256033a6ea112b26a31ae0292f2d6fdc74a657fbcd086;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ac9f8ef26b5bbf72a06b730eddc165f828080a210b15f501477dafd896ae0641a1dc7daefede78157866a459a4d84463a42e5b4a6fb08b4a8088006f7b4d17c371fb45737b4941a4762e09f4031682271fec5c91fa12ddd83a98b2f57eac4c0b3cf93e9651ce361461369546efd13d9b0cde03e8b395329;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h177964d926de4785630d2a69e8af43a28ffed44de01fb2632ebf464bd64000e66a1e2403d8d17942e924d501dbcd1bc241386d3909376627e08b5b3efc0ebf3cb375a86bdb5d25420c56d0b248c2d81e83c66526b0e8805e0eec58ff38661394550f40f3f256aab84d306a513c41d4e70262414e3b80b3c9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116d3313683e656b83c30381cec19e2b3819e653013eeaa66f41ab0562213d52eca34a69cf0e38d17a466698efb958b3dc4d4b2dd1da5267f3665aef2f0098857aa300caef92ede35bcefbda41b308924994c67c1ab8b2ed33bc0a153b8a5c829c04eba6f35639869cb734a936451da995b4cff76475989c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19610ee6361272c4d89c7569cc748fae87821574e14306ae75fe50dfa26f69ef3f15d6245aaa1509b4e96e1da07a5f21a5bf66ac85efe6bd87ddd4cb887c42edbbec987621dbf93c2738ea4cd5b786468109eac2ad4eb07bdc70f4685d21a0460e56a4187e4d697f361e91b26a619481c2a8d2553b8c63a5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacea2bc6b70e45f5e09445cd6580110b81a9258dc71ae208ad86315aa567512f74422ebed0e4110dcd2ab2fa4fb22c6f853048d9182e4d266cadb70207f839581f744de3db0d58c2b16d35069901f4a0c52f16e6cbff0096408c83c9fcb50a49c965f6157f524f431a899aacc93069ab2503d91b62dcc2dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44df774b3cba61da20504d22c89e4a62df7f323c48b40e2ab4654340c31eed4975e72b021dcdb98403a5578fc158e0e2616c2638197088f6829f317ac6538fa3132ccf5f1cb30b5ffc65fa5da57b6deb502a225bc00f0fa0b277daf4d0cf7a2ece49dc8098ba2445b1d771e88dd77a28d22d6921aceb2a42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138cb7c231f9197668854a89013096e2e6bdf63fcfdd9a1b71fef427b3cce27e4399530bed18c674ec2e37dbeb2fee0890c4b7a745a6a8b33e3e7d3b726644037a85bed269cfaf9529fbf1a9f2dceb28294b2a46fccd957279e60beaf154a1c7df4d10d987742d9daf1080ca4f5cba95cc9ab11ff580154ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18307e1326feae93eb96c5804cfb89e915dcb80d9a78c4d4263257464cd575c9be1b99371754075dfa8f167e3837c22e69eeda076331f73480bccddb829ddef5132a68752483e014c7372733db4f2eda07b9f188d92da084bfcfdc08885289d97fc1e211a90ed40dd2b5d507d0698a9ca96227205b2896398;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h847a21ca619c2dc3ad44879bd993986365eb1179555733f818609f4b992b96eb3b68efae64284bb1934b87d38ae5840f776076254917ff1da845cdee61d22175899b01d63cf87bfa12fec970f91ce67f3644e42184a1c8f3fb12cb5df6e1cd7dce30dc241de39274f80f455f2ad1e4b72ed502944a31f03e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafb47cd6c8945325f3cba1c87d27b83c2e7725fedf1e425ff78a06d8b01721c6e861e21cbd820691fa0e7cf6c6af8d273fef586fb774f9d79700037b2bdc4c5983cdf85d6b61b203dfc4982076f6e02da213317f2a51db05ae6b223b7f0c0f30169d6e95d2c879a52640a49f1b00cc2411c03704e4ec53ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc493ae00870822929b411f9d15ef8447b40b6db09e7fce96da422401bdb5c570ad1d69357e16ddf8608129fa5bf9787392c5f63b5d6dba0514b3f321dea0c72f70b00817b709393d4ead0ca24ab59b94d8bac7271369ce9f0283ae777ae4ca368ccbe48b5974a29b0de54e89bfad0b1e39f38a9e91f0618;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hced224f6ec6c3a7c55b7b46e03b5e17a155886346abba3c2242e9c50f2ec7dd8f5e0d611e78c4fe16ad03a0d5e468b46788630e594f4a2a41f93fcc39971065f82a85216e8022d271da78a34630760acaa7d838deef83e39be685c34f7888cbd942038f6c21abada0cf76506ee3696948e644e1157b52795;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9a47ebc6c1618a7f30eec6108ff4290158d881b82381583ee42c657d971bed8a3a91fcaf80a3c2f5f4bef601f4756049883b16658e842db8360576fd993273438039d1b767dc7ca9f2e63e76c1c4bd5eb952719db540b0a98b0f752d8997a277ce890d373799b229d570b8d6a4f3c2d00ae72f0b2f701a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d38a024481321ee23f970a7f5a48057926c3a95ef56dc0f4824d496ad4306d15688dce573e84cbc54384dc11831358202ecd3831645c127578ff18b274e549e815ca978926c2871d3c064764924e5112d3e68329fff267164d99801af4a1c94ce035e3c5305e3986de132daff437ba8b10ae7530a1d5bbc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h55b30c960b1a887d7e5a12845d96f10b95edf48104fe7fc21ef18d81dae53c87b1a992f3c03e1472575388f0a79b83eb687d8a888bda0ea37e164a26cda03064683862bcccf079c5fff4cf2165808ee17195954f87c2a00d31fe2278c6a6e428eac72f68540fd695514f09d6d253980e2c28a3134af262d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a309f909a29e981154920cb9f3e04b11254e3d47799aed0b99e327c9a9a1d86c45937085414c5e59ac77e0f01b837f2c8b8cd8e06d443e1102fe2a0e2d52fbb52d653333421a48bbd7424f0bc3d980560c8d104dc849eda39abee019a0976ea3f8a612d01b2442d155fb08155cd6988b6418711e556793;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1661a5644621e6a686b46a8e6683a2920034a3377e37de708bd5ff2a6e53c5f41688eeaf092045b4bef954fa1a1503198083950e78458c3eb31d6e6c252d3a74f11840485e0910708e9acfed997552d7eb324bee05ca111064cd5c741cb5d0222bb0bca248e0acbe1573563a00afabb683ad4111742b976ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3145969d1f55231d693aa0a1c6f8b1c4bdedeb5a5ccb879b38a82ec8b6a7f989b591b95352c824e5ed639fe1079a37e24eaf696f9b7cbc1cebd41eb33c68fd1d385a1603adf72fde78462dd31e0413d2f8882f9caed461b8b1da5d936bd8067f0b7585001bcefbf75af794c16e1be0a88ede071352989de4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1443fd3b2bf8c56449b0c193f755768141eb49145f2c60c1c45ffd4546ef8b29d96a36b4981d305718e1b8cb4b7456d15ec60110f3f73c5440bfed54533a29d5970148d9a865035320e52e9042c15309439089c7a808d53f316cdc7ebbf525fcaaaa08f1c4614cfcb20f0c5af1478a6f9efebb508e02052f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3f3ac1fc1c3492074c5e92cef442de866497da73e73fcb1a119340333cdc8311101a4e392685859b687c795513d3b58ecda596740e8cdc220831e7d68da5008fa6aa2dc2c6bba65f69be7962b1c210f5bbd5972ddebecbf67feaa4664708a3e52655ef463506294cdf54e44a9ef7a41d229a9ef3ffb8581;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7d13d48ea10159dee91c9039b7774ff8d1e7ebd8b88100884a77ab2c50a40fdc737d2a597860249512c2d19f769baca973b62890e41a7bb1be9ddfee1eb91e84d6e32c107bd60a8a8d56cbb3c848eda7b6719bc7d02cd66ab02d3ee449506c71d67437d0f46b970ee4db516c1965cbafcf0f02c31eee856;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6cbcc012909b5ab4ff29caeb2163ba6eeeb2b0850a2dde2b80dfd23b9c2ba4bc304d66521132148304894dc23abf907a2ef4f22def2939b4a353b9fa670a23a7670ddabcdeba25e01518d54b8c65fc4037c0ad60dce65125c9447af44925fc8fb30f98b5c4988acf637c67853401ad268e5756c0f4556c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5496d7bda2f270dba7c498eac4b6c0167f4f8f8c46ea20d712e079c41dd0d051f8c7526ff7587cc4aee08050eaa46a4487c1f7bb6742b65895340284da2f8bb4d74064e6e4f952f36fe55eabbd2afb1d753dd59214185b7b7f1069f9a5a72db277897bb6fa1a2bd399f48b783b876ec4437d1e697e7c81a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h479d74554682a1373fa463112fd7ad5c8b3b3632bca9fd2a192088f992153fb562b0035451f46ae0a820aa03a1dd7e0cbdf3b7ede1e05946f0440f41bdfaac391e16c131cd02371d634c474c318e6065aeb2232fc26e8b72c1173c0120d9e547d68d440bfc8e85c1f05930d5e81a8092df5c3d863307afcc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168dc88e03a3c680187f6df0b18457845bdd9cfdcd7d57d5c0ce261d5a3c64f318ec2941d4f6d8fc40fcc27f44bf289e5303faab4d6093d49782f23d7779c8d4a9598ceadfd39a4ea189090202ec313fc85a596a385b840426fc029f9d468cf80ac9ae2a8a2afc7d2711c20be5e7dd16eb271b24c90fd2e45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18584c3f5612cb372331469b2a0fb71925b078998d5bcb6565a8fac8e3405196c530d90226f54f65c4e714366418b69c6b0dbf02bec17a60ef02241817a04b7b1bc28aeea9f95c2705e55fbebf55abf6399c7ec2bd5b37fe00d8d25a8b2e8e44fbe7ed5d29cfcd790ac4e8613138e0bcba652d54d0816d6bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4aa31255716842287de6df0d670f3fa567491f3964ee4c1ea3c7409748701c694e560f1de7010734282f3c578bb3313ff1e28a23e00f8d08c8c023aa1f1b684143da3f082867cffdae80d0f9ae5dec9775ce94ae0693bd4fb7b10dab535432bdf221185692ac01dfcdf6d4905c5ac30cd5ea67868190423;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186408181769796489476785f7ff8ca5d1c7ea690d5f8f33804199f22508595df023bbfbb60fa5e372f4c002902ef897e2430481daf6e0df0cc0630e33c1dc685b4e2c8de55816a0a28ef7206ca189905015dcd1f699f29afaa0a656b3b05bca536812dda4f445d11d69c787cb932848db297db8ba99291c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198ba868714cd5e06c27166b3fac98deae8f3546a273d20474739a0494bad9c1caeb75a3ffee0a34b09c183de0cdda41f987815920b4228a806c7e9c7a6d11e8ee0e6ae6b7485e4cc46a1006a6ec2ffd473c71d81206aca66756f1120f94aa4191e3e44c513952babe2ece911970ccb38588c0ce8305d7bad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3edc4978d1b64eab0db7f51be40f77bc724332c9ac587773df4d45a091481549ab43798b512d845a2c717e277e6267e9edce3bdc0de07f4cb84250e3d77d2445090ff2f631f3ae7f4f75a4c560b3458cec4344fa1c3d8dfc7365e3eb2c6206115b6dba8e1bbc9026a3237aacab42ecb9aa1224526a481686;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f8d688598dd3c71a7a2c0472ee9e9dfe9d950541813666278cad489de0c200c93df0412fbc4ab598b71f560af8c39f11769ca8bdc73a1064ce65d4bd96dca9ddba0864617661278ecaf30493cd7414ad1e6178c44991248e2b49342e301faf908a6761a50c2eec6eb6e36cce2c470d785198e8f5a65b5d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161503931a173a7ea5c8b7004bfea3e0ab7b1f3b75643b2008e5be7a6002ccf8bc973c55376d55f355694680a03d82181040f2326d71d2b8f5cc0e894412aa4070840e9af0ac45d257d05e82b91f22171e8aaef3541bf384d2b805e29d9c6217d1bf91812ada9e8ec89b59b9ab1a97a737533896fe82c084f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b54426534bc33e9cd6ad3d26ddb781effaff80e5abc145b57c6a812b3586b77def08244686f32615e4ec7f5482f6d3aa836bef70266bac884118b640a8cd46fb31f9b0fe207ccbc56faa9442691950ee699de05133e42a35a6a089aa8ef9cc66ae0d11145342acbce54cc7db9a643df3c26fb2f33a48b06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h589193d64c1d46bf9c4f19d207a0f6f4b982c440ed9993acda91accb328a10b2773494155d31875420b59fe5873bd582ac82fb23d792e42c08856488e2ca84544fd80169147b24891061e8a42932cab7b89824b6ebaad88373f22cc53ee40c96f92d0e9703408795b58adeea9768e753328a50f4b637ab73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9096ab599537dee2984a605af6cc4ca2f11bb376d8c0a5b647c75abeb7d555956ef3f27a0c7d647ced2dd1e0bcc1f53af8df80d0d154b48cb4b486e1fec14c12b9bcb37a81c8e90b3ff1784f02f31bc0acf5b58e83d45b2c6884fe97c700cd6d208fc3ed51fbd01c0e54faf29306dadd96a5d630961b1067;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176c229c72294882bcc8251d82e6595cb16ee6800b1c7813972d72041e5e47f7befb6dbf06da75ebd98399dfb96a60b20807fb092df9f1984bffa1e26b4245f5d6d37ac0b10d8702e87b9047e6f3ab2bf23bc95cc4f4285b82548fd9fd9bb9052f24e8395baeea86ee85c0f3d0964950d0af8bc1d04827a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heceaad9be6b3f5b91cf93ae4a2690027cfd5a381ff62e4e6cb81f218bdcbb395c059dc8cd54e3c1249c4b897409331b3789c12616945b4cd9561a07207c07b517a3fc9a5991fc07b9f9139b99c4c2536d2c5cf23b1ec4a4267157c38f4872df494f52ca95eddc37a17d9067cfcbc4b4e7b65c9631e196b18;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac336022a45c9120143dcd57dcd5d6f9a7a47d07d031728061c962dc253ec8a1fd296a12e7d06980a3c2eb56d66b7ac94ec687e9dc0be04665f50a592050927592945687e99d1b95fadbace757c2fe9c35723cbb2c365c5d0d63ab46c54c78870db2a30eb2b8b8038f2149d5470ff50a1fb2a7d041c43465;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb081624c3c37980e5248ccf9a767c4b54d39e3749794b2dc957a960b09e482543ec2b42ed0b7ed90e88baddc36fe822f5a3d5929c5131507980e5b8ecf949afb8ab941029b4709b4c838eff74c02da0d5fd71dac90ded2ce5becc6aa18ffc5da78be0b358f333823a58c6a70610ddea17a0d6ccf4087e7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15be6f6446719258b6fa477d71cf3a6fcd7ddc58c5018d25a6dee35c6cff1a9d48d6a8dc6077e2f78113ce1d51b4432148aad7582690fcea02989bf9caf0632562dc3051ad9748665fceea20efb13a113423fc4de70be0a4b06e87e767de78aa59c2de19864794e98348095a070aaaed080576c6d7fb16d69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e8dc1bd4725ebb3f92185c6164b905f337d8e35c890d2c2d47d6375e5b17d0ea820592e2d45646f4edea2481818a3a43ca6d4fb4cf83bf49b2fb0dc902f53f3eab95ae2c59b9f0129e7941b40e94680b98cea5dd3851e1e123e173b92dbbcffe3cb0326c363462b467e3c1e61f75c74ecc07c99ee9899f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e20dcd3842dd4ea823a5de5172ad4bff6fe90422c3cb792716de6c4f3d4b9fda64a681ba39a603e9e60aa5e938b6bcb3abb299fd6c402c8d8839455a38c0bfa883baec61c1358dc0abc98a5b97b054a4eb8ef1f2f88b0d77a5aaec0f04ed374125577730837e1ea18f1c73524e217bc3b7afbcbcba0a160;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132597b2588582f3764d5c44372218874829e5c22bac877f403e3b7183dd1b8f6ee91271a507eb9b46412cea3e7e5d6218713c7b1e0f956ebdd58b2fe6f470e590bf1ad73ff439a9787a477ab7bfa5527f226d44ea668bbcc8dee71a7d333a8e7fca841bed850127b0bab439fb29e6b4b1bb8c158b304577a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1002f5cf34e9158347e221b20f292072fa05ae7793ec896d3e8b98dda4c513b522302054fbd5672fe61ab71e32863bfc280b6404a33c83b9e8c080756fe57926ce2ecddd941554b9dce70108aaafa85c8f6a825897c741d278a9b22a9e19911428c07d9bcace40bed1e28762d66ce264cde1538b77b5936fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b73816b73ecf92f7e13fe61f47b9886309728379c11cd9d03525c27cbe1d8cfa079ea0059812d15f91152b9fdfd95bd6846d24b9c8fd056a2d30f8668e2a2e7857a3e9144440d617af954278baf90b2e7e5989019a16ba3264c2716250bef3faf16117b126e61493f10f0dd2cfd785d7e27f1c7d97d642c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1925b5f1905e8a46efd430a09ee85cc23d9232c92801bbc0f50157816dc7f0e3b5e4f848641e943645a1526bef809d0c8884d04ba53008c205ca2c624868e30032b9a3437c12d97eb8351b24ba83b3e0455c035832063c8037d66ea5a4e77212d638a7c84cc53f5cd058ae175d20930746e6d72e5a77e96ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb19ba3368e6926da0c34b4b7e50311bef71caaf8f150ca7b505f07c926b8dd84a274f36cacd5fa64d3b0887559ca413fd0b44ac0a1b57ae3f5baa34787253346e93c7d8146b4ac386ebe92db7e4b00f0c76d9e5d7da76834847d9cc7fdd86737d0a03295597bbecafbf0b9bc86924c56ad433ae318891c0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f6364aa98c8472e6d2611b3dee352a247cc670b5e2be9e9ddae366036e03d889ac096daa11fe35122f0984420c91b802d7a3c1bcfa94d81a448be846851ac9cd7f5375c2d169c83e5b53930399343884bddfddaa258f035c67b430700bdc9b29ca1a7330827afdd01022e0606616607fbc0bfc5e03b3721;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1811dec6d59af249a5ca699ab1155b376dd5eebc2bd9f5d35a1d4c1e2fcb8f7f76a27ea5634bb37d327de559659f868eace12430c74e3d753ff75c5c3dbfa7d851b53fa4b7733332255cf7f37a7ee520e5dc7514ea5ea2680732fafe049a32d7d50785aaa468c17db067f7bc764ab27a7adc289a4f37646a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c497ff217e05c9c1e3b0523cb05641149ca1ffbd9c1e27962889f0864ada680c956313ffeaa7428ceb2b4284c21b1819a848ea46f5ab2a47828b24679577980307efbccbaf693570b1c64b7284ca4e9ca2455efbbe7bff69eddc64997ce84a7944ea5193bc15d76f2f4c37f941ee59cede53f1557af2e1a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79d89f0658e388dcc4aef1acfdd7f0db24b722c940bc5e8f8421516d4897aabac3736dd006aa7594948327a10bcf9e012ab1bf8f5b7755cda1a2c6536282db86217ea1bc07ad4acb7262e0c7920a4024e0c59a45a94ae1b1a7a22eaac3a77e14768617d09858f4fb4901555093f8225ecb63eb2138c843b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c5ccd3e367029973792cedc6b5839988761f8d4c4df6c4b304873fdec69687f9680cf3a320d85e60fd89dca6c343bfb138571599be2e8870c171adcf38fe38a58ae44c5802e8001c9eba26d171a35c36c6c16191150ad034284e5424038c0c4d4a8b2f32a1ed465e12152f5732bf809293e9dc5603779ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c65d1d3dd41822e06f4655e67de95044d399463e5a49585cef9d87c45f7f8f4ff12aae674b09c8f19fc13689fb2b00ad95e3a2a7acdaad71e12f5a24187eaad2bdb3e9025343f9286e26377eac64ccb49593117c94262b1d6045392a81052bfadc829401bd2b6040f04c2457a21f0634d80fe66d8c5ff783;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165a97cf7236b79e7375f6a14b1c0a7f9cabc0b3892345c5b0e5761a7dd1f67b352f0ed3ee3c45db4c1e3f972e4b61cf2f00d13580d02d367591134f55434cf948015245fc841fa177dcb2ca0710fc2299af7155fdaf90f834f3cb6cb7233703c23f4ced80394a975266dd4e37110913b79f7d3056adb0961;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e2b53083bd5ae017384c3c3cc3d646f73ace862bfe93b0323bec49795076aa19e62244be3d406e07458731f0bb126dcf2bfb7b6d954dd80b231ef672647cf6bdce078f9ab054fca1f920f09d5dfdcd8614686aef2225fada4a11e47cfdca9a5be279bf645b8871481564970a3b3968f01d961acc20c17e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdb787eb9a47ebe0a022fd00ee0041a8e50339bab752b0a1c2fd6a399c0245bdaf4a5dc33f921b36bdb746fbec41525035bea4d3256585ccbd4842b09e4ca46a70abd35fd56578e0eccef0fa93e88fcb8ce905c91521cd7fe9cd3a7bc8d537e4cdff5a4889b3ea30340600202a77af3afc73bc95e96622a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d20f1340387f7f35b48a33497c0d9eff01f3a30ec68a44b2fb3f2c6322eb0310c3b71239862d07dbdcbc8f7ba1a01cf8c510dd57142beb8cad74179640a19e0b80e39b3f380904bd0be9625deac6b8d5b7786e2b1ce3f7124b5e07156767f5e8a5993f2830b95f06524cbe5624571b0d48beb5336819864;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1275d8e5e02b68e7a1a669f65b7fc07627acaad07e97006491b37bd36d4addaff3dfd796b4417db96ea13f4e0ea7c1764238c63f276def7b6a70fad302e3e19ccb29d5813c5a3e091851dad109313bbeee34fcb2ce5acf8ed72c65cfacd5cc1500da744b17835b2b1da44f7d608e407c525389ae786e77f1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f73d6c2b15bdb8219bd1634ea7e2397b765aca212faa1d96ac4f79e3099fe4a711581755603e2e1623ac71a3021e354e9e95565e0f8aac1bf2ed5b3aebf7bfab9881cbe1bd6e79f8cce21aab6949f526b27cae493dbceae1dd3ff6d5d7508aee131533f8ae2155aa786ca130840543fe31b43c95f16293a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12dfdc785f60c648c6b2cc9bcdbd6c554eb1bb9a1a6df70a19c72403fc0405ad1ba633f2379a33bcf12210ffc821899dde096eab0d01641812cfd282175899264e057b9c6b305ef7c15ea10dadcace30b6f077d4230936f5e1f4f4d1aaa951c90a9a941f68b2b4ba25d26b0499ebee4918bf0ca9de5bc5ddb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140b8361124fb53276302df298163b2b28bf60b9be899502810fd93d97a4ccdf34f626a2317f2ef8bc3273bf6ab939828ead9942281f36ffc5a65b45d1ea55f780bcc6c540cdfe3f5ec16ecd8fa95b9f37db9a88297b7b9fee8051e71745d60bc182f385c326441a40142252ba19902ecd0636289b6b9e6db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee5ba58ce39b2c3b2f6e2af0fe492c21f4c8cedef487e3ead16a087b60ce99904c12fe1601ddd7c2948ecc1675a173f7992afb7772bcef24675e22cebd2babe924ad42201aca838dceb02fefe1a67eeca301f185646d5f53ca78d821d9e91e971caff509a88a039906ce0af7b882d313e30cee06e1463824;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad363f76e5df1c64a16e54e3668d2bb7b4cee0ea9b866aa5b1a217821c582c42d6ecfee14c40bfba7d5df3a08f5e3903ed34007200b4358b6ce96a230a2c0ea76a82a682a5a30d69b6df41af8f35b235bbc112751393248760d47376cb09fc97eaa087d999ed54ab73758a8178f87a7056463404fc0b1c7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a28633dc5b90f15bc770baf25146bfa2f495f8f9562fe0de2475b594b3544b0103d4c4dc529cc03e4cf7081ee68ae9420dc5b0bb302705ca7b85a96e36138d6c8ce7ae0e7179a6cf3b653ccea50aaaa7fd43a7c286ddc56d2d527a5b0be6480a2e895dafae2cc0f0e925c8b3d6cb0d72595f875b1cccc550;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h791b4fc84571f00f57b1307e3feef922448f4dfd83302f7544c2d894086fd1d51124d3380d065262fe680e893d596ff2130c63ac80de8003398f01184bb3a792e8bba975f91b33c815b191cf4395ab71381aa7a3ce0ddcc0c6eb4a16372b80628a3a615926a8f444755842d944fda1b566ade94840cfcc5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffcd31484a352c03a7a48e9675933a34c3d0d20336089c5b9f2f0a8e88d466f22ca09bda63cd7cc8d14e1725a71328cf39969650fa1bd58007f32f21ee7d9bcb98a021af8d12e8bf7b9f6ce13a0ed67418b5c3b5b20b7c8d942c4ecc68425d089407619f08c5dc726305021d5e4c1ff791f419595e839366;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128d0069e9ebc54cf37bdd0638f3e4fe36f5556d2970536a55720424ad59fc02da5eda1c3ea7592bbef7cc45046caaae93f61ac6e48f3469375244aa4541852727b28640706773f23c9b1da2260726e2f620f135918fc94370362306253ff5b047e24426091ee835ab41d16fdb963db7cd831316e10ed0453;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf56ed622a2d547faffc2b4cd93abb349255b2ac39b4f9b665c0a0f0786979abbeb5320f2b99cb5e847179aed650466387eb04d0c4b3c750511990f05c2fdcea042e06254db9cc9975cc55b536161f4b0257fc3a724ac49eb4cbea025a96ac3fd433a2b43c32d2e6a844003ffb28af7d23858d881cdf6b796;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdccfe2c4fb0db58b638d816e944f04913c3541a560e81d30d6f32fa1dcd4d5ba2940bff394c7a8975db47e9331559cfd2f4786d50707e9a77f025345a445ca67503dc017dfabbb3f34f250fde3e44bc50c48e16c401b50633ce60c206821d255d33fb29e7a5c5a56b254fb85a9d200444b101c3420ce716;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h969ba62ede1d10c2a28e717659cc7cf0900df64ad7d9d182005793ef0e7986e15a2a59e32f45cfdcb999680e8aad8a03e8ef8a415cb2ad2a4ef5836afc4e5a3c9d52a38c33d9cb2c2175a3ac70a2b38b2403609cbce2bba294f2655663ff0d7780609fa18a6a4015194651fb3dca709ae900ef418652240;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51eef8a0c83ea1f9095c73064b5d279b805f3945734fc0ec68a76377e7408db3a01ef600eeab640337c67aa132d4c53f726a255424e6f7787deaaa75ab37872a62cbed87509ed046acad1dc6340b806b64fbcbebff8e0709af4daeb4bea3469ad331338044e425d030de0654d151fcf3369c085435e2749e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9044a8f11edb7efcd0b1e9902d4f92b258fad34b4acfd4e422afe314df80bb374513ec4808dfba3e4134a4a6057559b8733f990606e4ca5bc01842c9780258d64f7261cd73d7f54851b6cbb6de1c81eef1dee3a0e8cd5f979957c434950af68323cc86ac4a5b0c452a1264cf31d62518bffb648d62edc50e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7092ea70d8bb102005fbc39df1a32f30fb4ee220336e1fefb591532fa6351901047f1dc2845d071af6aceada4d62b61b9113630719668087f968a286d8b44776ce7c9ed227e21ce5a5b499214500df8d8193af09f5b4be7cb39a26c5d9dac5826ad3f2007ecdc1b423831cd65e75d9b3275d2ea9cb7ddd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de17df187000f6f09e8a5dce106238b3b7b63ebc45e70f1d7fe955b5aad6e036364181c6b211be87c2f2efefca7c9d884abde224b4d471b2154da5ee89b5029b17f7984095d7d260cc3d5eb61b3f207308f077e32df50690a55fa48dc5afb386ec0c0caf9e0abffe5b1cfa32f7e20c27d23c110ac7f6a64d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cdbd4e0871fecf214e143296c030a5429cf295ea8800f45368c9b938a07b040361b21f27b6f7ca31726d1469542878ff9bc23bec28e99bab617d32c3d3b694801c07155cf00eefe627d049c7ddc5bac4192e4838716cc94627b6289a4dd746f8d346eb502ae48e47db641c4526515cbef30c1a26f933cc7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfeafb90e81e4a4c026e251b803c94cc0156354aeba78e344124a6c1594da0908946a2ed872e7b6d3ab37ea91d3a5ec61d6bedda923365f6c0696c608da7a3cd9e6f1a5f46603a698fdb1d05680e4d7e7d234408383a93239ab4b5e311f5584352f2a60a78f1284a18d0e0dfe19aa28b5e0077171f88207d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40574b562fc25a4fbc1a3d678482c441c6a804f287e07a2b110f0f5cd4df9708f6518a4bf6ac0f9788540f4c73463114c4b423123596fe32f8dccbae10c8ff34b53ecae7f12b8f71a4f69825fb6dcb5b995d341f84493c58d80a28a0b4b008df68f23d2938c86d421a71e7d973a627ce72de4342ce72b19e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b072ff2c7c0b948a603b085a46f92c1d620876df63de3d4a72cff810c2f902cd4be7505c8d2ed16fbc3d4b9300e189634c21c0e6813b1c01280490141735694b403de9d694d3a9fdd4c22625778f4ab6cf6174f0047c16ebcbbb060787a5b703dcd920523aff842b37d074ff852d647355072174a2819cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6e4e1c290fa6229d12ebf5da33a564fcea46f9aa355c0775e00e3ccc7ee8f4f7a165b06e54e83ab090ff4e39580418d6e9f587d7dbab23aeab049699ab826e8fc1a85faa9e1d36cc9511ec83c80d4acfa9ae919cceb2a2cd6ce2e3dc19120843ac1ad9863cbb31faf0edbd2f4ce1bec69c46ba146d3560e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b67564edb7203e4e65266a80b6f71b7f0a13cd8fe2360ac00a5df9c0cd63e73052c2156cededf907642b1b96d14f9151ff12ab185eb945bd4e51aeb203f14d5a9ce0c1f6043905b2caf6e25fe16bd294211a9bc7e2cd8f21d078d79356cb7f6a8022658a51275bd706e1462db94bb533a58b2788a8807c97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3723b281887675b32b6f8074a32a2cfe51a18012ce9a0cddd5335c183f606973577d76bda98a022aa553fd182ffb04273cf7873276cc8383fea88e36f0c0425a641a3df0d6b7e00925c3169aa70a20eec7aca496aaa8bfab788ea7f385cf0681f260baf5d3e63f0258f0aac651f105929fc84b076cfb5ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd09e8ad38f61c850373550b484ae6080aa6cd60c90ebca8cf3957829439664b3ec33c569c6618b8e68ff50d34d6f6216a3885ce8abd68b5f805fa9b738952f4ff41b5f0eacaf231bc892f9a56ffad26cfad7986794fc6bbeba27d5db2c75ca776a00d81a953051c04f166fda6380ac6a8528db76e03ae85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e9b880a8181d4788e3c3e7d2a32a201a54cf7826db65e0632d0b8a5c5f360e7e683ff39f54321fdf1562a608fb6c3d64534d751bd277a0039223b0f0f4c8499474261d1f240abd50fadb1b82f2d8360f6b017bdb235deccd9be84b812029e34d6491dd929192914382eeedafa49013f6fa1547a9e007484;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfff51a40ae6ccbce690d21a7ef816a4609ad0685cdad32b4f1bc778899c510face3873b6b838472cd7fa85ebd18b01d4c2210860fc0e075bc4e3e6205c17ead4a153f178989ea8aea87bad2a95d76f787cc6f7772e4876fefedff001f0c9cb2490cc9126a318bbe37b3af9b929dba3dd1f13008e10dd1a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95929e4a63717d5309db5485b21e960a38a8d88142e1d587111a9b90c597ee73e7e96951d5d8809de463d8b2e9aad9729fcf8756b8940153112332534c4613fa578deb72e43b1715c11f0422054ed8d0f28561e6023f70e5ff9deee63aa8ee55655977bd2764c1a2fe5c850961c6ca16e896d259157cda9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd14cb898e901aeef5245126bc70335769b1b28c043d88d45cebf3f8afdf4153bf16761312d91e1a1de2e5a0764e2b041c49f7185cf5a0a1497e5f155b862886ac513a254c8034e354a7a34b25f912388c75aa01064592d1be5f61668905872e944d247434f120335f3ba8afc19dda0e40afaad6d2514029a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2eb1089e1bf57306ef4614d66a0423b9536b37fa740337c58245460eed369dc0159f2d5b4f5bceaab03107b46e62a015ad56967f4e6cca99f4834e85fd46f956998fe32ac52e8436447fd0834138ff97bd00a012f650c5fff2cfe228fabc370f96669413c042521129c5f78ee271d0f8df87f2825ce16c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18bcd136b8d44697193c7e05bd916e04368ec10d51a91d951648cf90406a73c6f40575c22a66ed5f173e731ed5336a58da7940cb4325e49c2683c8f9b1208fbe40384acf921dead6a0a419b4d98cfb82d4ecb8ef936f10482c5c49913df6a86b268c49fd2d7dd42cb6d9d8e8fc2d57e5bb33477a9badcf103;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f1d2a15f99340d118933750540d531c95bf842d02d4e320dcf095d5230f7c1ff0bf30ab81f3696967689e09bbc92277e3dad3bf487755d1a570eeafc42b08fbb150316cea9055828d2f3eb4385a4da4f712e4f0011b14d7ca0144748b8148bcaff856b72542b3a4919c74b274540bace74280aa928a13f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1a264b6dfa9b29e7d24fc632a351f1c5a8ebf976872ab05ac52c13aa9865ea404722c90a9a5c7831e46b668ef996fd6f04950275b0b1ff2f4b9026cb2775f067b1a75251ef2f49c8c792808e230fc0e984bcce5b1d6ae8f43bf50b3e3d7c2e338bcd4065f983479ec5f22e6ebe2ec941c9b331d1f93afe1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf15b64b96b38686bfb754a5b77a790d8e526095b6c105ce1616dc0563ef26cd4abd29c0d67d7c4ab717d460d2daff05c28c72c609345e3c97ceea7ebcd68196b7c59a950b7bca00c4504417195d92fab94a3c533823c52ded492fa809ad6f418ffa9112f168e40a1f2357f32dbc52cc86092784a44099fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37889cb8b705913c53c8960f6938b6fc0ade36f099082bcc6bc4d7d23165be09c99f9136ec9813fc785f5262b12ebcdeb720f63b949a875b52d839b904bf7bfeca7d78ee0e2a2c8c97c2c6ef087cf865b48abd144b22090b62754e7d1d97325c9a8342af952c94b811edbf5381d2525b117fa1ad3dd754d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78c5165e2c1430f9768defb887e5151773355457e85b6ded8cb86fff617c5fd91ac22d952331ff03bd56b6737a498b5d2ed99aa65b13329a1577883456c2f091c7e864d757c843897c4b5c5ccd4edef86470463b9849884c5e258baa584c7cd0cb188c19102134b0465d2c1242eb163919ffacaf92276b00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b22e009ce99fd40f240868b7bcf2cbd6abfae8a67bbbc76c97c16f58d81c96f6fffb1a8b9af3afe7d9859b9101ca0767dc0536376303bf8c894f3b9b92a5e748b565a5804e81996fbaf096fb87e678355141ce008f12e741ed6fb6df9f10d5872d0a9ce0ec9aff90bdb69e132969c29a17a346d4fcc09f3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131dbab8e42d84cb645ffc52fb78774a7bc634c6e3c9c800b5d9320ad59d928c8c6d57c5aa6fcaf45f5a5db85761db363385cb2eac2b9c64b4c7a1841d65ffba5cd3f3672e914b2a32e3bbb23279a2d1446d35c9702d04972a75ecd5f85f5679773b96801c56ea5ea9db4163585cb645e3f4702736a703344;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1966c26eda761a2e52bb259ea66092bf377926961187984e7261350beee50c33d6d7a1c943307eedc23d3c020cf8f283694498dc54c6033c7098885f00ed13abff317c37711573d29a02ca183389b80084cc01e19e5da449c8609035ab2d205f132feebc0fe6f16ba4d77f6ad85cd4cccbd03f479e7fd489;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h326cd5b0ae601eb98111f61a83c4163967a1f535e3d6fe5c67f7a7193f52212688b15a0f643941aba11692a93bfad45868f26cb147388944c3de525cd6012c887e4e710f2db9dee6b2456b63011a643b8366e9526d2093fa247931fa327bb7d137284ab580b45e194dc5938ccf03b537253e69fbe785b055;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1023e68e1db4b1a273121fc3deaacff385a1c16c93b58367cff69ffd518c55f082bbcf16f2a0062d407e526a2f0abaca58d6917b7281c3204f5f5a461fb2226e99d6da3e602d9146687bd2119a0e0206d06baaa584a4f10cfb60f362c62ead55d7e761f5f95d9f881625210d79805955f464fd3f8a185904f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19951c90284d09b1d26bf0eb5f820f4db7fb39bf6466a3d77fd1d5a89daae1d475d9b338f647ba719fd6386279a33fb1219a1f733adb1ccd17650fe47681a5cc8bc359d09edb02f9bd8e2e4e411b4cdced0b5c7bc74dbe1bda8fd442e8a74b281bdc34dea1b6da3841243ad77952ed61cc5f52f1c89beaf24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfbe5c4ce911f735fc490cb071e3d0f624d97d2bc84489fffa04ecc020e5188ae75abcf75b633e718449f343f9021d02b10a05361eb26f074d72d47ed8e7d4b36bc907ab42c28aff2c88a6351a0972d3182908c214f8869cc9dc51abeae6f68ac5f885677091620b8d5fc5f45eaabefdff0563f65ea2ac63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1021f48d84ed2f7b9842f85a5ac31d3fb17c1baba530a767a58772bda62dfa258c3db6fc6209a7b778037abbe88346560d8b415102c578fb1cb19102e26b6e9ec854aed77d6098b154d9a9ef8d3affbe4893322779a76a83e1f9a227ed55d4f2c53c5e54008db904a75c2a81c500035b71288fd7cb3a1bdd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6bc1b5c8b4a48c86d3dde56af4a1f91c3d120f800040081455035cc009fdb6edd7a638bea2eede0d762d636d5cc0954fc369c20a6783d1f2d1724b8fa23210a285edd6cd09d921d216a6208d3a46ac0feff4799305c46cbbfd756258039d8fd96733be256a20c78eaec4e84a22c17c91dda1f797ff032df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87395513199c16c94989c74cfffb9b805848d52955c6aa12048c911de7beef5f597a91aa4d30cbb49e285e9a5a34fea19b2b2894884cad684af2b9249436fe8cc89b773caea46c24106e4878f837d510957ebfa8fb0d7c4501c1806242eafbce815dc4ca66e6f559c85eba959617e6a89088f61c8c097631;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d5550a2a344399c902ce99cb563b672e12af0bb7807fa400fad3f9a7a88dba0fb3a4a0ad808b1b22421e7485552f3b773a55abc689c324360959e66a81e4f539d8c190ccadc295b51ca77ee70f42458f81cb4d249423f6a8dea5b80aba80a27287368f0e71a5a1cb922e3a0535ebfaa22a068b162558446;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13287c9f03fbc81821efd9e98206914e0ae4dcea7b226c5eb26d59d53cdc3a75e4eeb83ae0b136268ee827bfa5c79d9eaa80eb1896cbaadd44c01a9c062507fa7f2e5fbdbf22cd59eaa0da713f02acf777d94bd5fe2719b4ab7cf482a8e350d9e88ce3124eff4fdce794fbee280b40371c43c8efbc7e32dcc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ba6d8c3d521ead9b65fb01d35fdeebfba99cf73700f8660c4ae70b9089006f7fedfb2596ddd602c5b517e33ad37a351243b9a6dd5352f17c2aa2fb52b86b82dc28406f92d6abb3fa43cc93cef7af5499856100e399cd90dc430b2f323579157a618b3275b86eec23c5705d3ab4e23dfb676c8e686989c2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1b3007efe24e30620530344920a6eb55d3612c37bfc5b6a3916d4ce73fdf45a3fcbfd4b8f966aa0c40df779585dddfe9c54506b2e9620bcff5ecb414ca7afbcd34e4f2c905caf565a04e4116a343ff8bd3dcf93222a78721c8308f1dd1457b43fe270370507b50a91789299ee0e5517fe1e4db224b85fc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4df46914b05e3b455fdd75aac988a4112b2b4405ec9ba33ae19f922b616275553875af0f6aef48df2762d61fc34a19e0308b5e18d63a83a9a31d1bc824bdc24799c077973960b0309c52eb3e125bfdf1ba0314726a51573dd8e1e8a662d4b47261bbee63d83552767e5af381bcb3b6d119af493540db9a82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198ad61a9f4cb5d200d1e3292bc8345bbd237608f95298acfc6b9c99120bb407e9882416b61b46b9d1efb831e601d6c02db79c41ce674ad27fbd634782dc004709e66fe6df0b2b7bd2428ae251a8f661299ed352c9854f77e2f40d10999333a349756e04db9b4591038ac86e3fe29cf02733834b89d49edfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15190fa1c840e5ca0ef3b39780654b516a48055969c61ca20d90268eee270617eea985e6289ad8915b856794e83e8f82e42ddee32e24728a4e5e09f1d3884197f723d2c52e7dea1413a8df7757808ec4c81b5be0e4e4fbc99dd9b85f8ba1fb718fe8d66a1baf80efb9e30f57cd6468b9be953bc50cc7fcf41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc6bcc8a83d8bcbd2af7491458d7386783f4eaaa9165b5c3dd2a4bcaeacffe53aa05284d5e03b9b656eb1938ea1dcd0eec450c87980f66f7732f495dde865654002cf3ff25f93e6aedaed32f682632ffc341fb4f38c56d7fbba7d6eb938755e6a842c684199c705254da24cd45fbbd7ea6c4f6711a165f98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1370bb11975aa92c716e2d45dc1892b01ea01f97aac539cba89aac3a9e8d0e93a93efde11e6908ad90d6d9b0a97415d03958246b3a756391fbad147770dc38542de7a2674d0973d4972927ecf44edb3c847968f4e16f271abe00f3d3a120a14b5864db40c6b3025cde84ce948658ada44294afdda476a7fbe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b89ac89c2acd5a8f18502baf9f9263d694e9ff057b76a2d959847b7decf537ac0da3e6d42e0668a14974facce2642bea68bba3f0127d272b8f6638d73f9d49f4ad10ef3bd56f08c2e1618bee95e00f7559f9462809c6b9da8405e2d9476af9b07f5d94aaa2c57be53773ee5e091bb93f49e444803430879;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c602ab8e82f0e9e785a7ebbc7429aa10a72e8b96454f4826cfc3a940c80c3db9b935dadeaafca88c169b212f66ffbc8c8bf668983e1676dc606f4634086b0af30f8d8cb3bd4798577159079d7ae2f0f7ec49eea6feb19f6001cfd930ff77d9f966d1bfd627059384bcb97fe972f7e58d90bc82e7df4bd59;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185790a0a4fc9d0e535d114f73d6db83ab984cb2377f8eaf8d1278f4b85f9d79f6f516b99ea03e0ade2ee031fd93eb855c35b8d4192fac73950aa28e5c7f326aa4f895a035c11d07720c1b52862a0b16df849a28e12fac41a1bb76d7b37c66af2b6edaad29e9bfd6e0041cd03ce74a9bfbc5f16ebe2fb89c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129aa0c49b1cf046b826d64be87d96d2fa7a49ebafea14d2ac091bb80a12e6884ea5596353beb475255e75d3378939ebb876e767e0c304f3c4929935c336c739205de2db2de02b25c5a3cc579739ed1db7ba8920a9b7b066f8aa2cbf1d561b0a176fd1692c2ab2e91a4bcfa7bd8381e6a2dbc66f34af1a1c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a523aa8c035101149a20ffd59e21f31299a41c7afa43d858b1d3a542b182862253a8bd83e688996835560a0f0aa5c7a2e8a6de3441f5be4d0b4290ea33afd4c92c760008e8ee6fbc75abfd894fc1935f913f648e861e273814a8acd595b37966709875b284b5f01babab4b80d5d42bbd41ebde899e05e6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c366e99ca108e5388c06e5d1abf2c0936f9d79550356fbd89cd1df1b4b88911888dead690b576b79a1acdec70b07143a6ae487583d9a5dcef12abfd378637eb46afe20cce42b4e959e0f50dd07bdd5b9ef8fc8a52bde0d3480ab047cdbada83f8d890aa5a65e7f0fadc546d32c42c7b31110d4713bde334;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88d180c6c5f2710ff929e7db205cb789cf08473b29aab5fd23df4150d54783368a134ddc207427b9c306e8d1d81c79f3debd80e32431cc189b0cec396c14e8990c34ab6836115484b450af612477d0dd1e67e2adb92099acf305cbb7bcbb0516c6c9eb3cbd1f08ef1d14b3fa83b7a0b0ea504e92f3b24c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150171413370ecf3def218798fed19087912f2e230abfba5a02d526520675c26e63293399c5128d5c62a6a05a97d816b401d08eac7bb3d94586527e32d9cfd96cda1edbe7e0aace7bc466d64749a718a0d3811f732a4e9554b1224c8f0a36a67954ed1a83b3a496490c38ef2bfd6d80851e98b38041f73aa7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b54a757f00a3209185fa70af5f25db573297a9f56155cbedb7e9301ea247fa4392058720ea62daf368631a3a1ed8c9efcc67709beb650c481d4fd9e1aea4f1dfd7f9c071b9bdd6fd62bd271ad4f749e218bad865e6cf0de8bf6e139210953b2d64585fc0d9ca7b2744d18330b78529d6569a476abcc4350;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b7c97cca6debe26906b51d033553343b544a5a34d45193b0a89c8414755006c288960818a8e73732a04aa9d3caf637a284f23e2daafcd1454c5c363eb5c5ff4d9b158d4ba24556a17633ae5ec2819e3994f6a98a0bca80c3ea4e70cc56c32d0b076abd59a44a418fb34d9dac9f113a75b4da5de99874351;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd2333730eb62f6848c1046e36a3fe58f7b0a2dc8655a3d4da2e56785132869e0d61e90c30b150b0b717d816360eda7bb885e62f90db17af6bfbd7ba8bb8e9d0999d44ff7f688dabced8a96882ce19912fe4ce8ce4e500b0968544824242906aa9515d1cead663135df20b73e138cc9f485e073ac5ea97fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h913951c973ff16c202eea0301e66d582d0f6c2ebc80988e37c35bc844982d8734deb6fbc992cd37ab7615fb98fda3d63f15f9bc6ef33c93bc15b7516ce8164f109e7a4368843949c951f89213f309b824ceb89a5d3a7ed41f288d85312b96525d9379913b52ca5940cb9af7160e81efe055e5a8ef40c8893;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7efc6a9f45fefa44dce8360de66ec0d85a2e9933d9ed708ad2058da05959cca305e9278c981e3cfee21b422ff568f20fa68cfd1c4858cbb019fcbf1352812bb86be5f0bbc553c008e66bbab8c8b6eaf3b2bdc31806a3f0dc96a48e85a1cba1a8d2b5bc7e4a7f9441a24ea5a75c12797539baf18af66d5b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192e66eea8234b8c72970e35b1875b1d2e5d5e1e7c022939f1551a097b8231d866c48c6d18b93b3d7aae8863258d458a2783f72d55a636ba972f0b8da6761057fdc483a93e3aee0dfb12cdd48c255c1ee2c44f933f8107d3fe3db3ddd5af648401c18cfb6b7d57fc6590b664741d6c6309e6f475053900231;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25d7bd6f825163baaaf5c70d5204e55c8775a3728df7ffe2a3852f4bb9cf3cbfd2ad13b65b3d21c9aac62570a9ffa41f0694ad89f6a619b227c683b38f8f694f574ce8e1f26fbff083adeecd13bb9514bce6f03c21c8ce480750be99d8d4929e757d4b8a22606f33e9e1c4e8e8bc1afccec7d00a59a2db4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf70f5b480d53ad5338dcd773a32a5d92bcb153655bf8292225ad37beff14e0d30f68c211a46dc2ff811b3c0225782d5466724841bbd0e88695224f89af64d619348db64edac0dac032f743ca1993c9a3924593360d66acb36ca219f04971b1d683fffd66e6a321fa397aeb32eeb1d6f35f4208d339ef238;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66823a06166e9d720e01a2c69d1f07e5e7c8e34e558431eff15def1144fc72febbefb27549b75063815179011111063dd3f1cada072759590d3757981da2995b24189339728c1353056456078ff83f98c37872dd2836d4d57126d5dc7b37d9731d78e3af10ea65d9ca9a906e360eab8edbab12d77064ee8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f853c98dcdf975ebc5c0f84d68ea231ae214a8841ee23f970173a253b35e5a4c075e75881a6fdc2f130b1eb0ec0adb223fcba81d29a282857be529e6872d68beb2d86b35b820c9deaf0667c73455793ad4c3c441bddd477beeda57250796031877cd32112b1c772a58334ac1d992ce1d3b934aae7fcd037;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7637ce690b939064295d90fc6f8bd2799175a07eaa872499c45a653cea1d1b46893e7d378a1e9d0576d812c3f491a2922fd0a62d96284c26ef3535612aea34df8d2940be99c29be096ff661c5ef73c7ea4dea73de5394d8847fcfce57247aac4fb0bf62b60f8933fddb0e05f6d99aa793b3699943c2bb843;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26aa873f0b4c584048cf1b26dd68037d7850711e116727f8c7515e170fb6e5d752bc7993c1c88693b395dc41f13ae0ca623fd13128faf5df74d94adbdf0be188ccf4d2433a2733fc988e72f7e5524564fec366ec4d1903d2f56c2a86e9666fb41ca590975f8b620b6b6bc7d65349419eb0d88464e595af42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d08f981b421741df09b534160a457d6e70b3d666d26e8d3595177cb0199ac25eae0c62a67005287b6da11e9f958ecd8e8da887ec4fbb84b58eb0bf90dc23f9d6258e550d2cc5d38713bc22308c1ec177151b051d74630a06d31e690d423ccec2f7ce8e47635c9085fc23d4e4a6683c5154503ad5c662bc5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee13e7fc87811e1f2835a447170ad7cceeb8facfcb4adcf05fdae12d7a3a84225942661593c0b7eebc13b5b79bb05147098a7b3e39a00415870ebf26963d8aaa0ca00f238ccb06c07203ce832ee63d39b447a8aaa345e2a1710f916e38fa0be8437ac297825fad1cd928627afdb48ede240e4883c1388b05;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heecadd6d66c3a1dbc2ce027bb434f63beadd037ee0cd823cb77c390062a0806a7ecc70baeee6cda82b8b2db664dec5a8dcd484073d4f0a241063e8c0d65ab369bf641894c3379fed222d372b64b3d2588f4fe82b2466c8b932b085a2895625372d0dc8af8391f028e321b5d534896882af8a3a3fe8633633;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9938617eab20f09748a63e82b9cbac0f4e10df3feb7e364489398f52c981b8c770ba5e5eb6b213492b533522c7457bea282a01d6350e1ec7ac451592938ae9f0c349562dadf56f73697be4dcc2fc4f6477b36c6b643edd78d0726979f86ebf80b1c6d73da9a9405ffae815297cdfc9363d773066fef30b8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7d6f30703d4430d8c3e7fcb0b9411f0acaaebddd095bb347e531b90830570db98d2d3c5e50bac0f7a87ecd6ac5c4e66520c6268e546bb2cb562e9fcaeac68e20348dcaaee36af4d43965182d336e508cb8fbb0ccee111f8ff9f02e288cf521456b0345f6604b5105f06eb59661f7794b72ca99bfb738c13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h495fd7a16c45a1aae1254ad4028d883742fda3c89c9970d658df83941cb9997a3771a4df79f8f0530e0d5dc30afa4c783394320b72498a7c5698de943964af452f10d5761d24bf03a199de1d2e8feab5e6501bf5318d00a6b4baca0ee8437109469116315e425b47efc17e291b388501a9253e20b24a4261;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc194125f1d5a582fae91249a71cb1e4a51d35f3cd79b837cea2d8fe64be2642566df6885c5b8be4f2a2f738c3fd79ce9f8de1d05c248cc12a1486545be1978dc7170becafbccb6e9a59e93a181f0f943c53bbea275dc0901b81d587c94c0168fd5556ad3584b983f00900db9492283d58ec899a0ca6d989f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1865be9bc082a9ac2bf59e07c796ae3e3f30065bd51bdc118c30af2cd777940b92940b9b0a0a6be019ff36ce8e8dc6cf18101ed510dbc28d14c245a1f9eeeecea7a0e29d40f0ae6c417e8073200a3d4c08134f83c30e75d7e413421dbe0234d210e16399c86ac0ad8dc1ef174df77abd662278d77a5636a42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13dda8e05ede7426a6d4380b4334e4cc52193dae92b7fe44653316970b7e58ea58edabecae8f3dcc5af762ddfd6d39490361991a7308e12927c6af6d7a90240ab50fbcf7d734f12633c5b944faecc5cc1090008551146b1b5cfa192a49d30d40e75b62097e5a8b9345db1afe726487f5e0816367656d26c23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99ac1e3d250df839b2dafe7e4b4f7a69c17a1c81112b8ffc1c260120ce9c558dae8300ed13bcd719fd470fafe186dac5a6fa675e1f0434bf5b76096b73d0939684770b1fa3f5c591b7b83291c83367f75734870510ac0427c8d4540fd5e1f4e998d7490b2a2a72b7a7ffc707e15c3989fd81f4219d7fae8a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58ffbd2ddebeb5cd60160f65190d5a4bb89299f7939f0776d1cfb5896c6465f900219dfcc11e11010722dcd295a53e896ec5776701e02187733f5183316eb75c1ab02e86dd8ef8194c960f9c71eea2c608553fcfe3817ead0146092dd3067284a6e01742aa8083ce88d39ea7b5d006c0b544c2da57f7ff6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf42e0221b15ccc69d89c3c30efabda00d2bc114fc4aa3d190213b4a2c20a721d51c7ad43c4179b4a43d20718bc0faf3808ee98b004bbba3506ddf2bafc50cb461d71aeeeb4fbd181385e907d59568a7ee80154486407b091fab76f93b635f67e7ac7e61ece381c2b3a1a9eea306a1e09c4961c97ea75a222;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17900ae63b91a8d363b317401c4d16e10d9ce60e190d4ce602867225c95845f19feb4695f584fbac4be27cbc1e5d8369716af455be8e4c44a451952f456734dcdec12a437d3c251a45124e2d976cf490d427d12425bcef0abeb32e10c5b88e116429ecb423356749e919b450db3b4a52266a667d868544072;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e680306c2f5eb7f950420783c0e3892895895059b24fb9ba4a7618fd50cf104ba38491ab57011ef701179af5b96f3fefc969cf21fb39d1918edd134aeaa1660c29a37c3dd925e0a80e80da10a1ce9cbf2b2182a39ab6b0ad6634aadd5351f81ac2a48be44d335203489a39e3a98a2a4701c15b5e77c4a7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5afe729ffd319dd5200b1589f9f09cbdf5dbdb5403aa19ee072c46c930637bb95ef8e191b0f9b005cad0a28f24a41f0e4e6482576d6d95ee8f99f0b7a642d3b64703232212d50aeaf518517469cb1fb1ebb6ca87640cf22c0d1e0bf671fb2c1caee04e6e2a53de59c170b1f4380cd4889f9f271328073e22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3c4faf898e71dcfd687a66a2897e71a8f0f3550e1972bd87fb71127d5f7a7c94aed90e22eeb2623293d6a0591961289ea70748387b3d2481d92802bc88e58879ee8e6db6210960b64f81460287e862b1df46871ac655db0c9c4a2aac9726b74b20c6380bfdb1e591a07c76d8e7c6fc25b3a95cff6f3c86e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3bd52407fd4de06ebff68477de500e7770af84f0194f1add7be933788102a74c00026450b98b368ce3cb9b4fed5afa86015008ed98b31955e557ee0850ffdb5b3ac1727d822e937ef59b3e5733d4209fa73bfa1bf42b1ef30a3bfef5aed15056523cee6f6314e4e259281ca3382365e813d752ace4abb35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e36088afd1306819e1bbc1105884ebb45154433b789f4bc9daea7292fe07a331218fc2833e4d66f46fee6c510fe5079171f7c16b4f7bdc919a2a71f74a9fbd0eb77a92fd5bf46160d6cc7758bd78e991bdedf0edef010785d108abb1f29cabdec2f10b77607e580bfae218131582313a28f7874194b5a5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6aaa4f45ef8c9e4619d3093444bcc7e99fa5220670995cd60d5a780927d05839523f73175783624f6ce948864605f6a5b40dd66bafc2e4215aa21ee782e3225fbee5e262199f99050dd17c035ed6c0f923aa3271af53e49facc7d8076203a688347362588e3e8f269d540497e0048c1db0400b0f975e2d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2d69f3f0754c647fb44c6609b05c1cae6e9f614cfecc8a1644f190c4fcd997bd8a7a3ebebb12a6620d11a8a896d5029d9bebe2c4d110f8bca46a84283cf34c6244c1b741cb64e06eb7efe0a1ac411d5ea283fa30544f64e4abec7abb6fea3145b1fb7c534ca42e2af06987b55161eac28ad36c18f8c63fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1039cfc4030fe535d4dfdc65935280a41ee2bff197189ece8556a0c15d9360e138a28a43f11fe9bcd925b4158f01e87898e6c710f1700449dae02950084a8fb98a87cfe86c7b49a047e2382b321f726ffd5e734cfdb891379af43feb4d5c2241fbf0640b45cc4556e149d83c96769506e3c46c3d95e1c0145;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1275da125a22653a6dc6ca1aaa44f343496d202693b076bb83aa98fc106c788dd64dc1e1dc25998d17517c1cfb6ef8038fabfcd35ec6259d44ea2806ada159c893304f344ae6fe2548ac298d7e362634783fb2bae519afb5a39a78dd9abac820d9554b9033d7a828a894a82cb42ae67af5391dad4d6bdd152;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a7f907df59157b229cb48383cc9eb65de2b0a874c3edd16b253485159874e803e5b722c56f6eac3e5b02e9705d7035fd2563bfee8e3c73a670a997ebc49910eadf5edcf1b6732452edab5c7ead32841a3ae22985478f67c6e1ecbf1c520936efecf5f50e6fc4108101255a2560e034d1c2705a99dc40272;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31374ca7fb38d56dcf83ab56d9ec9de8ca70376967df8acf6b0e63739a7499ac21d6f98112266ad8c4158d95a6f63a0e104fc8b8e2fda91bc218d41d23951c8c6d2248e100d654d7000d533239d2dd161f15a9b596a08976927dcc76f3449cd331abfbe036c095cf0d09e0bad0d678d3ea831da75316a48f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2b6ae7a41ef4cd18377305539df71b95450a91e23da4e1452d93145aaa2075e46e222f713af2ae89a99e995063bbe30d464948e7b18e4d573bdda4b2b87aae14f94a737703d7753a7c0094da53ab40689f5d4b2a54343f1736e32ad768a417660fc9e526876aa385175d79f7dfd871b396f2adc46285973;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bfff06e20753c1ac802a40af129caf2c36c6a0179ea31a457a713fcc57a3a125cc67d356c17e201c42075258226e23cc3a7f9df729e1538a4d2d58f52f705cdd20df97700883f100cd3a9a1c825ad2f631bcbc5a22f619b14f6e6d9c87aea4c21e15431eaa087864ad489a1201926bdb5d5cd6c9c7a4ff2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1407bff78a2e15e464a02cbd762f7636be83cda9be7983cc415858e6a9036ae8c4ccadd2ddbdba965c9cbe2a864c85e9be23b0285d182095302357de8ca435fad2ddb7ee43296bf56eaf97fcbcb5bdcdcff3a01aaf5c1d00caef5026d6ae7e8b333b4ee1731818321d53f117eb8831f224f61b98b1a3bb509;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18631dbd35b8c79163f2ca3a6234264db012cf30eca4896e62394e74b0cf4d989cf0e8ece91069d2743f57719e2ae2d2a5308d55b719d38226eed5d30b4bcc2e41f2cf0275f7b4191b5b1b390ba4ddbec883daf9de5cb5da033e71ac37abf9c0bc08fda2d5b1c1ce3337a42c795a7e160ad42d6b3d2a94424;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d44dd7dbdbf10372188ba372b7a974d4becd6e6415b041cb2127583f799cd32137e249875b8bb42572fd3ac6709cad055371ed8cd21559ae052d4db752f8174e1c9c530554680b1d3e9c8d5c362aa3104b2621e925f6ba921b3e88f899c8c6c5ba0d431ee005cff19f6553267c7228c72495447a9e342507;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191ba78e05c6b8fba43105a3da9404d837962657a2a884b9071add8890e862879b5c5aea5b0e64179851b8fb61a4abe6c15d7f23f4f254614dc59dd815d4521934e8a83b1c0fe273b9a8eedca69fe00da839806710e6d5a8780c55663fdf74634d960c3277c350da8b6f73313326c73bb922e5b93d1b81d95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d600a01e34be5daa5de345b041949057d2b728e2e1ca8c1581f4ed76c39a9fd6504119acfab7665cf3da7bd4cf5aa5530baf8dea0be8f2f83e1820e97b2ce02e1642d379b193009b4a3417605ba1360266c440372ba7f3ed7812c8e41e58a7e34b881fc765a945bce64ac738bdf988cdac3fb2ca7c7947b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc43e97d009b7207cdcdcac9fbe6aa95bc277f4267b898b1c1101c960a595d7f4a3a0c6e883b8e449b0d04b0a43e2be716512181fbbd8e8ecd0aea3c748b70ac123a2611139e384b446223bf627572933019f289aa9359ae8bba355f2d7a4b63ad94646c9b81a5e6e06a94b76ee4dca368b4c9e46da7814ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h689e0e44e2c71a7404e9e3df9ca6273eb9edff316a41873cd05c509f6d21cb8acb2926309f2ec1556cbe2869c6e06e7fc580be18d0ce3f4f56e9cd00ca0074ca5e230b780001e6734c70b194cdec4960de228a6e23059864ac909589f4c556df964bcfa5b28e0845b2514d56f201ca663b5da91aa42cca27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53bd3a8b8564fe9d9604e0e8fb7e90e670e754cad215e5499400b2f9bb28145431bb103bf023fbd6dd35f8f2d61462d25fa1a7d29ccc9294fcc4d03f29f7f1611d069106308829bf65821513ebf7ec70952367afe33706a6fc4daae20340f06908e35cf8cc26c312ca553f68aac1b45262f41d24accb7ef1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h817722b375d840ef8324445b8d5597b6e84993b6815d867e40cb3d7978775e42a83a3947277ff60ae082f6258ab30ea5179776aca8706fef7e5e3b17b80cb844058a25e68e94c4589907b1c4084369f2cb023c0ba93aea3fe3023c947a1f455b1db2787a9d2dfd2c8b86e9b35737619ba8e754c80d349148;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2bca042390eec195b6a47a21fe3aa6a32f1181ea3c8976f434bc9f77add1c66437c899a2b0488cb7620046d7d617c5874a30f55c4f62d415e3c02592e54fc1b0a6e8fdd4ece29d43720ee5265ab9e8c83f07eaba7982b751c99906863e1d551692d6856817f0a34631600b380ff07109a3b2424c0765b52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8c942571fd05eecb4873271a37162970eab46c64df331d1796b5c7edf8f3b66ee6a18a9dacf233d00adf14e1a41366a4ed8bc03a531cb1036d3ed69a9c0ede3b9dae136ce96517888ceb54c3695e5406426ff5118602f032e5f5441761bab718c52fabd38f1e80a323040349539c9ca9f6df584cdc9475e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1462bf0b655e1ea503dd0636f4cbab62aabc3e45e02ebdd8d2aeb558b8e4b14feb5dd5cfabb81adc6e5bb81376cac1b562ed65eb010c9d504bf41037fb254be09229a75f0b6988fade54e458e5f3e43910f6074ac65088c82e7786f0e8c7687b99caecd44f22441bf86c97ce660157a7f049738abf0a0d92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb7db0b2ec9090e0d2eca2705db3dae61e906d6230fbd46e75c5b6d6c06c00a965a92fd7af2cfa908e807bfcdad5ccc40f75785db7c353822973662d7490fd647a078f5f33f089137dc5b708e307312dfcda2fececd42fd4a27587ac174d204d8c852a1544fb9ed0fc0cd8b1e4332e986ca79dd5349720a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c531d82bf37832b21f0f672172f8128698733e62e823ae32b3a3222819587412ef23a67111d24d67d01832efa2353f8a20c9acd993465b0007de695aee5f60b8f039e8fcda3536d19eb8e41630aae43af412a2c70e7186daa124892ccc6ef769c14745d3e5bf6ae5850dcc91c0955133e8bc46a5cc250d89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9ada7ec1c2c1bc3d0436969a2e97b9ef95f2c9fd6350d9dd8416b249d540be464957956f81558b9e751604556a4eef99447eb9837e610688984b9dde0a3ca84084035398b5061231110e7c219b5fe68f956bf9401b598277d88c7b38ce6f5f881280fd16c6d3c75a7ed5750e4cfa08a0df118d70258f70b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57e23f544f2e5c8c6eb262915545f2443f9dda1a9ce24b88efe7c1de5a26a3c0f8aad75d5a8cfea059211a0fc79c3112614604bd4b4ce9aa8c0632f5b5ef4bfdb5a0be8495641530fe9e695ff8847082b364cee880ade9be7b21612a8ed9cb90faecf62120d17269ec6d28e88c46a1db0c46688734c17434;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b682012c3f13040cf9c4a34ba74c9137ec61da6630de9f4ff7ad4cb41ce4a33ee3cfb39dce3591621cccfd78e3a29a529d10d0fa321226a1f99885d8344b56c9a4898e9362c2ebfb8f734f843625d68d955642cac8a8740f2785d37edeadb32908bea3bc9eb69cebd31f1df603502cae0a1a2bb96d0d4d51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ec1b1816d5d21ff5118d5148859267c04bd04ab4ab1cd4b7be21f452bdf0eb61cd1dee7a2e3e50fb423e808091fece7dd530150c089889cddd7c04182b0ef72ce4c7f633d4fa1a4571fbe9f9a36d1f8b7dc82ce6a34d3cedde354272f5f7140cb4295e82c7dfe50fa033b0e99d97d34fbdbbf4b3c032d0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc3af9eda08ef15185f19d14f932996ee3ede222ef582f63af1de6b62f5fb66c7e328e8ee1695fe462d7adce648a459fcb452da4a5cac30f7d8e678255a74550b4827fb40d37ae7959a3789376ee478a684e8bb4078c189e2b344d802393348a4bb8bbfebb17bf036ee5f8c03b91a048520b91abc2906b81;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae52d2c3f29255be61f396f6320d224dfca5aafe5883ee64da840dd2aff864dbb32a5c29c542e85b7e790ac42b8ecddd4e94ecd61f4e50b1a11b73c17293a51a41bb78596cafba3698158d9e395d2105e658a22830b7284f3578f13b2a7fce63fbbce616e4e6be96128ede42f64dfaf3ece4060f70d990ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fa9a50dd9666f554ad7a854f4a16a563a6be76f39aa28e8e91f76b12f22ac384127d8ecfa4eff0d14f3868dbecb59f07bae3634e9f2895ead48aeef262484b070d90d7c23ff43a9c2e3bc83fe5266a4b1af6c7e7a3d92e7a822ae648463c30023ddb7d841ee9cf6ee77bd8751daa3a4b11f2a9ce3fa13e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1713196b7fdecc37604c065ceb07d374e9974368c5702fea23c8c640936261ef2f7df5ecb655dbb4a534e046132e3905ce53be279ad446c0cb355141d1d567e9db39ff0513defe072d37d9efd4cee221b690098dcc37bcbdd9610af44622111db9e358bed8cdb38dee45ab6e5979f648cbd8b7b8069351ad3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1504a40eda83b28ef2e13d0c1589bd2348f889588fcf55211399021036dd64ca5a34a1f6f6de6ec3f99877bec1ccec040e005bab159864be147118f2124753c55fbb20119995b39422c09093efa66ed6d0eabefc85dda1b803a8be3c7ef06ec8810b1cccc3256815225d1adf9e1f7671b921be68a7dd786;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d6e1a76b18f1f9aa4573f4613f584f135683375696e15edb7f77fe6a5017d4079d7ca0a8c3a20749ab153176d3d9077900218dd47e132fa5c192706d4bd2c000c443443bc89ed8d5f8269b876960a0cc33bdacb9bf090ae70c435a7e5691b7e9b0eedbf93fd50f4cb1f0ddd611affdc21d59bf26c8b55d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd15aaffaf7bcc587250383161a434f1f6cd0d65b89e0393e06a6886abfe4c199f3f6e0a6fee6fa078b7e00a58b99c72ec7b71050665aaf1bdc303fced6303dee42a2b8707f0dd6f154548c15c607e20e988ad07d401b02f04846a5f7cb52cb2dd17cd3a123f512c1d6ce4d02698bf395fc2169e9f9247016;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3da57a4d9b7a30bb1e287d4c4adfb696a4aff62b18234d8874f298c2eb7e45696e90d714da677e72271566a75351346de6dcbf13cd746079bf0e46e43e753a1b17b601128fbcee5b472ebd98b3dc3a5fb96de2ba0f0bd32ead4a74817709866dd0264a53434251623d25442d9ce96c6bf5c04561bed49bd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151f288d47f983dbba9299ee192b5ab6a0ac309ffb88896a81e9fa402a261bef9b8b96ee3b936fe449878d10dc1a0f925da92e635d04b8eb906b1b58a353b76e93d0efeda07bda53e14b4646ae4d88f6cbf8dca589ef2f33525d22679712b098c13e1f72f43644418a4c3dd8058e3df1ce25a16938bc22512;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e679dd2bafcb530d75180b889d7c44afc28532a5836b796ca660298dfc58147e15673ec76aa7f5a1ec8462bd8cbd216e76299d1044b1d41393772368163c497d637309be9cb69ab5317128bd4b56d76a909ea9b467a67004f70cd46a39b5e4b599d0b39288793891d1f42ab1617201dd700cd6c912745c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180d532c5e190a0fcebfc7c9d1e0b3e9930796df39864ae51390c437a861018b65ff24b4c61d22be3fe0464e101d2407d219a904b63b87bd3a267488a3e8550000460afa9080d179d1c55ceff0a34bbabf745d061cd8c9bd95a2306e0e23944d5134db47d0dbd4b6050fed0c388932854188e59011a07df11;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2de7965383b8e4670c9f8ff183b1ac6670d9206f40cb94b205cac3cedff32f7d35c52debe1ffda851b6f74dd0427e4ebc00916d36f7d30bf1724fc3298453c5b901495292535174544e6dd07fd77717cf8b1221366fd996aa5fcf1aa3ce09e5793db6045866aab4dd1985fa6c2d30cbf96b390caed66694c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d9d2d7ae1f3f1cf91029334f18a7332a4828af7e6e437b795996fac05725371ec89d0cc49ac0c28423e9d79cf01bc23ba0c2809532913f4432b6206883ff9ad4992a573e11f4244a91ff3494d6c810b3c7e64caa34cc5ed632311ac661d1196d95d63d94a2e9e0ccf2006df60fa0b9feabcffa57b96ac49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12df3b9fea3221243890c973617e8650f61662c43ebcec8bd4f22f0a9d0e5a90703a8a28fd43f20fad4a5325697ba25f8e3e8b4d071804b9fa33a6f5b216389f02ea3f145d6770ddc596bdb151242c9473e6a693262028b1efbc1fcd529f66db5b7abee95945a0d6046d5e4bd47d461c0b0eb8f45f2f3d47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1061861f1444a5fcdb3fb3fb6a467592bf1d4b544fba4a55b893946c1e4397e54c7662ea56189425fffdc2348f36e60cbcf0a88cc5f41ab59eee2615eefef0d114888469681cab18f72d996992c18e779129510ea9be0501e3154e45c09721ca2a9d7984cacb4dc45732c239c85f94f48969a6dbdde45ac88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d3e5922a824d7694cdb3bb22f5e555ae2cf3a984ce4b41449fedc8aea650a2107b3da66227b9485183ac0e86677e137ee81e231dd72f6d48b97a3c9aa9c4309973cd681f01c000f94240cdd15675341b911d93e299578911d8c5a2d3e58ee0ab7e897b18ee7cbbd10e10a3f3f9d30539680dae52f478762;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e570b962d0394ff6f05a680aae9b58c77c7e5f9d855def74ad8a6186203e2f84807920b137225ca1eb18b4135a56c3377aee7a01f9f0a205b2bcc6733d7d9be5d72c0b5be74a2b545a3f804164724207ab406c89728dac7aa157feee0f1ff295767cfd9a806f718ea65e9d1213443c5434875dc2c02eb16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f8b113ddddbc75b7b668c8a6f260fc65019e4878a8a1a3bb805cfc87b63ef9c7242cbb05fb7d22278621bc0be6aaa180cec7d1e4d88550714ad6005571bf4d28c9b94314945079166486c39d1bcef2bb392619378887e6ef9d2c786d7f7f4c6178fc3968d26e5e3a29b8bbd9ab9a18a1098b2e3d11d9a46;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h261fcc13c8fda69391dd88f685498170800040bae0c1dc06090dbee6db0fa7e7a1b4ad6baca71c829ce666e6febb44c3367aa634cfbcd0946dbbd07fa8d579a87c0819f451e205c4c655adc420b53da7d8b74a74967d682f6d52e2f6b4e8e9dc55e8ff80d24934cac2642f0631d04e9b74a4d41a8293dbc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f37d5f92bb10503c7e896a77d5350103c8697823b67c016650650a0b99417339959c0c8a49c1ce4c1643811f5990c5bc89f8906664fa9f0dce805cf3396fa476bd065d6ff648861276ad973b60b0afed7f43651569a8fbbefc96255dd9ffd4409db1f42bb3c566a1b5d04d5e0f1cce5b58da0e0180185b30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab25fc50b653d275ebf2fa882d265c3281da874ea6df5ce6318cbd15df3e8fbea7131cd4011468c69389e6b025d2ccf60dcfcc0784637a2241ea2fb7c52ed7ff1ddbd55a2dfce8ad4c2939aab06c2612c775b2897ad0106745b6170be48f3fa0a90b1eb983266276bf046ee848b88681eb3b249e55ed6e71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d274a00e18b5cbcc96e0ba9205d3a04098e964836dbff417a1d461c8aa3a620ac4f7daa384b41ecb879015f2a428d99fd9cae5213dabcdba8b362aceae5a33fcf78d63c697738f6cc863fada83ddcba7b6125cc9f3c4f1531dc98643887f99d99fd43846ac7ab9aaf142904ef9c84750c7cb2e3192d831b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3cb6484f6c3bed72a2af9049f3d58c5524c52f976b62ab152d1f9351522db5d229cf646ddb713c004a3e923a1f2b7b42422fe82f3eb996d25d3bd29a55411fdf32b2c5776420ec039ca2023a18f06f969c113df6396d9cd33d62a6c6416ce7b7d82e3f29624bfb627c99a107d7894b4e91449cc69b74ed64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12baf8e64ead6aaf725cf8319da0a5c3ef7b5590c68eec7580262a9d0f7652194c84f5956bff03dbf32241e9ce5107990f09e7027d33c3307966e2cd4e2f3d5c876c32100d9e2e68522e594b23f585f4aa1823177070d2c4ae33be1775b2336f784689e5d4ad1b975855c2316e72895cd0179fd00547ca115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1958a9740b5d8e6e16461186f6f172eee6807ee70195821b55b97dc5c031dc41170327465cb49fa6e3532de189165fff27ea4759213ec44f03ed72bd8d3dd8d6839e740239d401fe4b5e95ef191eef601e7b80ebb883cb0df4cc62998abc0e98ffbea385a32ad0fa8ececccdc91bb4f0156eb8f5d07fef248;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf299d227f6904067ff648d750002023d8879c29d1c842e95a58df7acd830b7525ab7d973c057b22b52eab9f263f8a222bfd9cd95e9dc7300e4d388ce69bec37d69ce1b67d325d2d3bf998b8cbfe5f9f1d1e086aa16c57a4eb37a82f78d99aca162c2cc4e1b61368aff1d5d9789cab5493243a8b07babb291;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bee8d611c65e8f4bc6f653e2df250615b4d9851dd07261109550d3f360fd47e2a86d7c383e4dbf4e71087cbdb93e6f2f8dd41a9094376e6e14b77834a9549e8fb16502b57dfc4e2a8e3562558e5cc3169d0c0548445aca4ffb83de382d74ecfec1d23a7db041dc8df04f930a97411072abc022ce94870cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3081f846a3f17634073582ef74f356e7336d0df63f855cef15e88db55763278df28deba2e6fdc97210528448131b1742253453607b832531f301dfcfb835e94d92ed376944410dd18bd5205f05aea7fff2a96681c9006ae8dd51b041d39b51454e67712d20afc318d261de9cefc98d89d148471a61641b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e39543693e0a4a64b8e6aebf67bca94940fe82e2d4ea8eeaa1a2180ce70f67b0599e0e5b0766b1e3306f78fb8c992530f06b76fae2a4c9f1276bb7eae4df49304169af2c1f9e798113f362c597f811b938d43b9871c191516406423f8ab87324bde9b4e14c991c723071c117c16ed05bab641d99baa60e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16233e25bb4a4b885b204df8fca8639223008f7786d9234b01607070d09ac6d8fca47a4c686b0452728eea593b69d01f81430b7bf652eb2abf3dcd8035fb815881a9c038a15e9d1605631c300c0b4c56a66c4d0620f7554f25b7108ee271ea8c61114d9094d4df641cf963e8510c23d44e61365bc4348c2f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3304bbfac4f1c3d77ce0603a486c823f39f600346cf86206b568d1f450961ebe0b4b8d499a5a4ec40da887ac7194e80deff886f0c97ac1635d1f431e5ab30d82dab9e6a1deae298bfa03dea98901e17ba7a345b2a8dca46c38d4ddb973d129bde304ff2496fbfbee962410865a898c42b1824ef2432a0e56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc33f4e90625b72484aa11451298b9cdc0b3f89cda560baa489a52bef0dc915d9ec86608da9f5f1bde3d467ba416f9f09097acf925affa2e427f6be15d64a9a51135cbbc0eccff94d529f34b0b66f1c0ea7e06cade8c57fc78977793e23d2332a0f95492f9312d7fe403ebf988e46adfb3a6026f3cc774ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182a87035a30dbfd3ae6b0326d7dc8ef453eda8fbb434444ea98f8f8ee4efb1d2c3a0ceb95bce9b8d5a149e2a875cf9d81dea52ee90a150e116f7ea34ce0b815eb525eabab927487ebeea3c19a1cc75536d54e790e213c1bd15a8b996a3fc8919334f31d2ab2cca86ce7ba163862100a2b02e243b80f2acb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e07a4b5db324f780ad82ace1a67b6bd6424fd58ac0258541233155efd797065f084a80d2c8a793d35612d25c0f5dd4bc4bd8ca5b2c7520867d659cd1c166ccd53d7d6ea6072a7ba038fb2cdd189de2d1b6eb642c7e99d68138a011c12304de40e94836cf2c45ab3618f341254a655f8081a616509aab124;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb5302070e70ec4f2ef06bf973647a4520255b2350edfb401d62067531aba27bf8747a7a1daddb791ceed94efcefcc5ea8efb33745b71f18ee5115d035c253c62c773112f7b00b95d44cb72e90bada1cbcf77d87a275a2ba90b68e092cf9ab1f7121f9030a7dee64138cff1bc62d4b81007c1b1537d56fc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fff16914392ecd8fc6c42715f76df2cb342374d4f7ff8f779c01f4e62ce0cbb5ecc15824e97ad09a21c834e29376eff43a36fe34f1109454dbf9ae41642a26759e9755a8e7b2caa9523b9229970e4b0ac063efb77dfe3d6f7f68849a8c077545673bb2ef24b3f5a76cec661fa0192f701a9de694e4a78e37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haeb14972a35691341c363701b9a2f636db10059a9cf35edbb18c189870fbd8db96aac66348b0a56dd0efa9e6fff34a9ec058066bdcbed6f4415f9d123258d8a1e4249fdae4746460dbfbfea30817ad6ffb21be38918f2a63917cf5ef5403146df73a8f47f3b63d415959e44ace49969d9e8155b082a41957;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca6aebf0240ec1bd36c0c9e013cd51a4e0ab6d3d1e82fe07998efdaabbad97e9caf33db54e05303f3f50337f16540d7a2f3cf371edcde2d839727918ac6887ad86d233883c0a223af00fbd5f363214dfe09c1dc8ac0c2c638066eee940f99daae6cda5ed2efbb8e70f1f80792877dbf6f65f66626b62a3f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h315742685438722258145e3c66bab466c4ecc0936c9ea252c1852b02570fbbbfd596fdea9a85731de589c720ed5d5191026e0d4de7ec7851fa67cc1dabbd84106eff1fd754b6d9b08e58900717841d86a61be5341d46a40ed1309be9c5970039602126c204315629c77c8212965e670442447c074fbba1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f51e79fda65d4e7b49ef218decfa4d594f15c7990d75e6806a88c11c75b2ed79e1ae7197cc095faa7c3d3403ef28e4a7815630a541cacb33971be8002b3df8e01cf320d4a71c0fbdcc7e2c46482728f5b1728db67eebfa2a4eadbcf57b1aa1afc659c9608e7a7ebec609f0d4d4ea5cbc59bbafbef738e21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h946689fac0b1ccb7aa4ab0c68ce08f9c598f2fd590be767388fa0287bf78e87b6a1e383462665453269101bb42ef58a1e3fbeebd133937c595d282ee3c7da349e2bb653aa143c99251ac8dc915943fd5eb43954a639f90d6d613ef256fe0a00dc244a975c410750f3b3736fb3bfdea3f6845c20447273589;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h784da28c15ddebbb419c06a5f9b2d42389d56f86f722c2b92975580264a666cf5e17b63e92a4759d87847d6624a761686caf060555718fdb2cd9206685b919eac3aa3b2581e4d8974237db5bbc42089211d9ecdb54f9f6e6e4c50aa7691c7019e19b98418c11b6932da0d8812dcde15bb5fca99f5e2fee1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he12e50deb37634e2be45b6679d3b60883781a0930cc7f6ce310c49c4a43f2d7677aaf50135dc7e5ae76ca932810a706f483e05ab008c0a5669b722b991d46d2183a3da82edef1c9dbf2a64b1498d790fefa171cf9e75974d5682f5ee9d3df10ec8efe41bb002e4d23546c4749ebd8688d198c66aa43c9a1e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78cab946b8a999d62e60224f653b766ad01f4f606cf78c095f5d6eefec011985943cb5c6f3ea1f9351f7f9e487a7a0329e4083ff939a8660eead55a9240334f17c8966b2a446779e6dfbcc8f9a66f385f20e5c47572e76be3db21da6c1bc0960d6d7edfd870d8c85a34cc210db26e6c9a1f5b9e61c2c964e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3a7f116ee65e9f51cca777e4180ec2a91bbb896256ddb65b1145285d859e099cf2dfb0eb683250a89a3b570cbc8de3b2f4dfb81a3c72085002aa9b67589a676ced1763256e64fc84ef6bb0085e9d697d726513b119531ac4c355f6bc81d606b00de067da046bcb84e8bf483e65aefd6a8fed921228c25e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140fb9699e548886a3db946fe3da46cca38dcc5aba2af7a0ce59cfccdd1a894bfe2fcf3366851fcfe05e5f124785628e725133e986a42a55f4abc36ba4c11b788da7a596b562231726846d18718533c5e4269da130b2ae97943b5149ca95c3d69bd69add9f8a93edc61847ac9c6ac4ff6b942bc9a14992dfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b614cb19201618e134e5398e375ab09d0333dd1e8bd7de7f72f742fa328018211e7b5d37d055155e576dba32f540f2c08c65ae3cf8aee2389e6f853bd501b6cd38d5f28e57a1d84ca3bd3f7f2f090422560671950a549a0cf9d3884c34c3e6e3695e247cfbec4321c7dc5939b51c3fdc336610f68725230;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c58e60a49b8eccd20d524733917c756f32ca6b19954102c0368497c4a7dc4c100e478c5091e3c7f321e02603c58451f1543bbd9fec9955c8e5c2eaf5f1f59e4d4d0b97c69815292a6c1dd04118bddb3d6972993e543df844a2ceca6493e87fdd66926b618338f5563bbe5862406885c384704fdd96a9054c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1521073c654b990ef75bf041245514083d3b84203a1545f940cea005dcd6a6acd479547dc1bb3a77ec7e75ef3aad5f51f60b9212a2da742bed7f55b03e4da0465e58aaf84c8dcea44780be0565688566143dec39138d65ed99a48cab58edc73adc954a049c47b929f85a41b9618d7ddf6a718056e6c5efb21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139e265e79b6298f24c0aa16bbff316deabb1b966b55c9e66f2a07d6d74bb15a38ec34ab85f23fe16a8b49d55d15042588122ee1254d3766fc2c105beb3c8dfc1b5fb6a61129f7e099a4e00cedfc8466888424fa0d5a627d6843b013465a211f3db8c7d80cc7ab5ffa986ec53dc5a17d154b944359d0f7c84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a13810cbeb9c4b92303240db6d7a55b188e7715a3a70026bd50946433aebdfe809605334f1c521fbb077f933ccd0f5e16d018f11b06bdb7b755963fa80ee99d41102f85a6a5adcea980e4337a6ac32952c3de740568359c06d572f13d274f38d91860ae1c363c6e321103ff582e0f15e1e976c3d7adb13d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e6b279107adecb57eb2ada0b2f258eea29d5e73437e54cae6543d155c442db7d0bce9660deb4f10da0c9bb2cfc390778ed752acd8a78e86dc14302a81dda1a45889eabc7e347d4e956beb9a161dcedd0f0b80afb9c25083e044f2146c867ddebca141e803d573586d65c5da403e1877afd14c0d07769fb3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b0b2793ff32f5255e1acd619366293443d6a845746506d5fde4eb2bdb34bc9fc1862f38718c76eae72382d074515935403383713c5c64ccb59cb5d1a26ba47f50fc7b4d24f310364a56903c2c114a45fab8cc63745f534715ae72080baf2d6deaa4c8419cb7686c2cfa44f82b9e2cb79565d072d8a1b98f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea7ff9d429bfcb8645b606722af0d1a49457a30fcabe4444f488abf43a2696c17253d3818d6ee89452ef7380672d64b0f47f917e97feaa5571f537e6ecaf33497055d646f7a21c030378d29efd13bec0b27c93ab1a2ad94f5b30f1a4db7b4e122884f0a16c313f4d64f588fbc4bd5fe6616399fc3ab475fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18048ccbd795bae41494993d53c582f0e4575f6d3f9c511188ee9e752ab0b65d78d63bc6c6c319ac36f20cf8c79ae821a1ed8808e9232f517caf6189754db956f124961be2d5cd8da9afb93546a20498fe2003594d92bc716c6d08e437d509d2ccf2f929357a64125d5617d5f50a1794b9ab7f964f717067f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172139d064517e1dba9370fb0eff6c7cc42a04658c1f3b374c84ebdc9faaa58c7387697da5774b26d51a2e5e2cdd1afbe53881e861a8d4e207ca1db49b526ef94e9543fbaf24dc2bebfeed4f4ffcb3849b38cab5dd71feb5a742a2b19c57f42dba66f90d5cb69cca024f664c07987cc24b8050fe8bbbcc28;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4eaa7a3c2b5ca460be85b4ba5306212a38d5f1b4c324bb6104e49b19add41ad4c9501fe360270b8bbd0e145e297a57edd55b50f4ccf4b284042e29edcd089e493db50459850be5b4c305defbf9585abb96bbf96a4ec2641ce5cb800fe0ff7153c8f4d2d3d6a71ddbba17eae1cccf21b1649fcf8700416ce4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd689f7ab63a7894f929d1749104db0d4094ddfcf2007a160f7949962e224eced3589a83271b2668aad52d7be2283a4f39428746655255075eade33eb24c49372f611ffe79cb0e47845b108174af8f628b48a762668000ac31f138228fac740a006a37f9435ec024a678a0990d9fbeedbf2df68675528ed7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189bd859dc4fc241485d19f7fb2943ddf0ecb8e197b71e6a4989f013ac95289494ee70f7c6dee76a0eff03c6e5c70bb60d8717e28ec74d849c927c330f498ef7441ffc8162ebda4a27a7f674c402703be729e0c72df0c3a4cc54bc6cad2f1cf68fdb4833fa9ea8b6e83ffa8dd2eeed4eefc94aa7825f875bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d10f7ccc86ebc7e892dcdce6b8927adbb944eb2ef9df3b13f83ac83169931f7df067ca66d38f713723163ea6c0a5477a43f13c3e844e3bad434ce8160c92860e2b659fea9721783f21579236ff86952c72d780ad831b996adaa3e58cda9a653b4be27c1504812a791822d0a57667591147f9173f5f4ccc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc3deea48c13a2c08e5b38bd6b4c07be7a0d7fb4dd3526667b405b253bd27794f270180c2caf3ce64eab8d2ad01ac88745d3a7999af54c179cce05c67d99960597ceeef8d9ec7fecfea107c9014e7fedd3240f6c26763cde06f2b4ce72790a48cbb8c3020ccccaa2e9db0cda9cce3c70cd27018c55932029;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b6f644ef98333beb36d44b3626633c5eca50141236f6a8cfab1e4bf237e47b028c3fb4bde70b9badee7f4c0522bd9d52404c1e687a7f408924d07a18bd2fa85340e8613dec9cbee6fb3f297849b802faa6b4070333de36488229013c370035f6368b0849ce9ba7066b675fd2a955dd6cb8d7b3b91728a94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35ab25b22fad3c6636994c4b05f9da90e0206ebb95eb7f9bca4c34b55436ff2fc7944c54a554bbcf3937d4aaaa04500f72c436a6ee2399ff1f46c61ce680f5b061d44464ce70f30b2929a9232201f9aa1437ef7f26d951684b74b0e2ad6ad68b7d7ffdfef948ffab1b7766a9a608710e4f8ef8ffc93b4a8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c37766378e5a7e274798089f76c26fb9381a7ce780d847e79fd272806ac1f832f0c5bbeafbe2776dd39f873acba56c7eada077a2057a90c7bc8f6df8635bb20a610d65a2b2775e4fca664d1eab5cf0dfb7b99c884b12e402d1ddaa2ff68ff4cef7059e6229e3b7216f9dee9f93a1664416f4c82909dec656;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b9df28fd338620976c4dac83a766d1377247bcbbc1e806ace5f08a999056d3011c2fd023e1aa33ef47a6713b37c22987ff420d495c270fc4dffac24e36048e5633c367638a1109fa45c33fc61f22db7bfe92c978e2373ac138344aad841891fb09bdf18e7c2334aafe012f3b2b5f30a0d4ea6672341fb03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a45cb1c5087cc711a4442ed2fc7bd8799e1b6392af47bcda1ca06731ff6087810862c368304c2768ecd6089230357920c78aa598ed28db484ba0fafb3f2be0e7c87dac14a0deafd91546bc9b75fe110d761dcbfd8d5410376c814b0ef1d7af2fc1f9b2e363f5348cccff0f5bd072ebe39e7727b7b7eb0f45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f806ad5b65ad91d5b834852d6835401e9f27a12f41d2f39f75169e4d35959b49c6a84bd7c216d03f2f6f76ed24a0e08294dd59132b0607bc557dd0b41ea61319956f01972c75f99b48d826144d5be4340fe54d2e89cb4a94569ac9b0f0bbbf6b0df7d2904fda53b698115504db1826fa9e849cc81c752037;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h373ad527fcfd41d75d5c11a78f48aa756a395bb78c03e154cf33c5846c9ebdefe4d7c511f795049980aae1f21f7b8aa909544acd9ffb6fad8cba4ce20347744d9259be01a36645721383e3046ceecae2f41e3f5ef45a5132f73e3e42180195c35a526ca7166236fb780c9dda0ab5f66d79d17459c01e9a4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee0e156214510b45f883e51f5f9d656b83e920aa2fdfe8c0db741d0b8567ecf42879b3f00e1630d12b3755b3de1388711af67901942212be6f2fd39dfb10b15885ceabba721786d1e08d64b1c07a2c981cafb9dd4b4cd936288ba860ed1b9db2624f7866f5131e0ae56cb58e7ed934ec50f52e0753d48bfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebbb427dceb44db042119abca222852309ac918a314209e0903d468f20e372ffe538871cead9d5dd6490cdd4f82ba0de0224359e70dc75c795692c2a0751ac45ccd520e6d4d0250788606080a0bde7217941d83e02f4e6575b42e4c5cfd6035a7a131d28e1b8e2c66c16ad786dc6973220523f0e2228ddd1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f5cd69e68961c1b890229f0be7d8db93d81a9b34ebe580221fe89dbb09a5741956e970770c35c5abf38df44efd9aa9c157bc50ebd0107ec4dc7e241738965c5ae3caca706f71a53a0ce80985331383db6120375fedb4c530853d32d285e42b91973809224303f847f9357d696a9af01e14822fb45c263b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15352bf2eb63670d987a4a645c5d237c7b7d0a32960f0d6cf0e2e5c1d1b26abdda018b9e6f4a666db56e0b17354b7db06f89418fe4013be3aa0c1b9f769e30de10d997b97d86ca48e79ff087b20fc0d3789f3ec0ffaa9047f1336fa1e4a81b76f981911ef52ebdd28525d77c792899a6ae7c5cb9b7388a02;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf3df8f3e85ef3d47cf38434c21fb6ffc91dafa738ba02f3bf8d7c9a72d98dae4e4d75496c0243760dc3d38579601719054e565511d7026abed38b7c94e45057a23b8451c018abd9b80d9e79d06ac8bd0a5c6dc7477670f5867267c0371f9d389238d6ce4baf9ea7f14a707bcdc595ca3cfdbaecb946c33c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12994dd3f3ff328d3b49b9e3354dc813e1657ae6425f6d7291a1430ce91939b3d7e7e05ba4569cb55debb4a09c0649998472396b40567e29484586ed60a5ea48abf07003b3e56c6ae81d38e14acb0a9d7863ec2d58e9914f2609568179851bfc29129ece988e841e8a7798e2479895e14ee80e10b0ac76665;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c73ec3bede2a9ee1d84cac8f5a37f4bce8f0025c273f4bdca7dbc84c3b9790478b04168da4be7e8e4725b1703aa5f7a4dd1ad14fca3f27f0c0259f42c67de99afaffbfc88c5dc8008bb5d29290258c0d8a094464fe03e82dde13e3f368535bf1cd657233a44f3e98ae5ef27155ab6def6cdbfadfde516ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea9178df829d10214a913cccc4e334808301580ad0895fe7f0db95424338fae297db8b5b09e857114801235c002030f753f9e09313633f4d455ecc62cbcbca759544f117b6c96d635580183e6f15658c62e68c0340bc9bb38bd5e30b11f2776e5f1c1ff89fefab048e45e3e351a6c7e70f60ab3ea99c4fee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103bfd9e2763b23bb581830c7efab06a03b9de479e2644bed5ce4a08cb0b4e01c539fbc85be6579583015bb1c2b60fc8c8529564ac1a2eacf66f45c0c0188d0014f9847606ccc349d726886dcdd3e4e3492b35aada3e8c99dd3ad66bd2475dcb83990ead0ae4e3ed1b58bec1710c11ea67c607205636907a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heae64f1610c1a13f24f8e72f6e6e3530e0f03677389141c01589bf3eaca91ec30d4a7e71f1c6c34804f6ba7e0d005131ca484be0c1e1a9b8f00479bcf0e02083945fa4f2375ae012eb12db1b0956e943ec22ec0cf2ed322c88afb2927a7862fbaef2e7fc0ea01d1c22124ab3665d12a02d62df951e5a58d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86954ebd7f2559cc51655e130c8a2551d642d949d2b7163f0dfdc79fdf8308f4c26e01aec411b681600cffcdeb16515984efb73238e6feacf29f12a4eb9b9825b8910a5f195655f8017bbd5270d375601863c06ef5e42eb34412575af0999a9fe811b1245e2bf564824b9ba2ae2fbdb04574b3299ff7d407;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee3522d2bc1aaeb14e2238c839d843710a93df3515e675b9f29e2b7c806cd0a1a7c75ba4f3dd02a0cd12fa296bb6b49e9c942c0d3731ebacc974da888c90388ed20cbaefa52753baeea7e754e7a47bf15cb5d0852b497d603e179b302f4f7781fe6be18304cc0ba792b1b6e08caf5bed6c29f39d6b7b17a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c68a99a27711687e976d5afe19290d3e7e075ef5c0942abfd0fc63aaa7eddac24d0a54ba4b649d4b0385e7bca8880aa43007cc2eb356694b4c99466e41445328c0b610068ee68dbfa8b171fdc1235b0e252fa1ed6e5edd96e546748349ea00f726165c3522a68d396f4088ba4417f08421756099c9e42a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19579590d6747684faff343caa639a739b4765fbe8333a87573c2841c62127f23b3917649a75ed009289d3d8f514bbb2c044ae222989700135027115529c70c47d5140fbdcf2602bc56d581e17b39bae6e702d7a95a53b85914f7da649eaed47341c3f2b43a77e4617c42cea59349cfecca16f3adf43b8cc5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc3e8996818cb5bbf633fd21f0878c339b8a272c126581459d79cb471b11668c9d0983e131c0c6076891707685254e0fca287760494665a0beedc2c5930d66e2e43b2448566dc0dd1e29e6bcfdd7e4edc0357fb486d70a5f418cc05b8c9078358e2a061c4d1bfccc57256fd998337b127408bcf3e9c2885c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101497ad62ace0f712086daf42f446a755aaca33a08f6fe828c3db4f9c8e517f6ff72689e35455c026a638c0221b57f9ae5ab92da80c1e46b25ead6d94cee2649bba2cd71846369137f61d1dea81c0f7cae688ec872fa444c4311e2a552b4a5315bf53a6c103ef03d03946c382052b92632e97c788a60e807;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b9babaf141c01ff396da43eb2687076841ec196935edf0d5b4ab0228a05701205b68979c5fb8c80786c7a5e0c1c3903bee8e519cfd3883a12b5b0904e48ab76611a42e3857914eeb1a3c7396aa59c4f98e14d6f77116dbb68f199e4889ad27b69e95da90d3e85be1471af63e0c115ed651d9b0e11ea5002;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h331ebce23bda5ab4d20b34357ab9acad6c0b13cb2c1581e42f050dbc651526c37eeb99105e21a3103198fd06afb0017613205219829873846df7e9f438a079313d95cf0f7af80a9e8ffeebbf7340ce8ec1f6e5ef93ce17c55d1d51d2ca6f4203e03b87c520275cf082ae0d126baa40ff296996153bea96da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170a4964e3c0d684db997d3c5c58230556c1c4859c7b9222f1c98942d93f3dd10bfe22434da6ce4cdad691732cebad696ee39ef58109e8d929524178875eae5aa62baeb2e96cc95545ebd823dafa141973833c946331b86259e1968faacc019093379a5105e24787965e9fbbc2ad52bb0f821b007a52548dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7fa99573cbfe841e8b00d988c4190372d58d28014d2675bbcea63b79047cf90166def759c470748c38ffbde24f8eb50fd4cf4b6873d64242542e33b9b7262d5e30f12927536e5fdbf4549f922c4dc2142096de8c6d98483d6ef6c5c01447fe34dbc18a5aa4d0241ff208b2b9288f23f8bd0b4c5229fd5a4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b45cc24bd05e77764439133b4e4637c8c8b131fef58cfd7d44f33ec34eee1332de50308b33a9ea9708ba019cbf16e54e7037dc8175e39b4328261c0b6735c4aacfa368cef0a4b5594703bd8ab3976f2d4d716bbdb3b35b94749300b99ee1420a7c3c479fc44fff6cc59f13c48214d9dbc6b840a01928af0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc628f8b2a84c89b2f2e9d9e20382f5df4ba4d337c3adf24157c7d98a4cb545a2928ecfdc23f885d171277a0ba8ad7389c9551e09912cb5b91371844f608b20ceb886bb4a9f437fda3250ec944f579661cef7bd33f725713fac3c5f068e7b46191ff9fb69f9af807f9090805f36104fb0b49c330faaef189;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had476e31eb462fca2fd74f2663e89e1c6207d705bb7b5d7e37f4f0aa43c74d5bfb5b928edc4d6b69ed0d9bc42fec6c73dd64b4ecb462946c37ffd694b9401e519e13c45f0c295358c708b8a5a484c3dc2a0e8d9024a3c4413871d6045dab0a5114b8510b2a076cd7fe9f483ca70c2597e8f1890ca0d9615b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3af0be06c09a039c23053e839fbf2ea66df73ee58962643eb055f3a9e04259c4b6d9e12029ec83cc14af580dde5834dfb25c703078158dbd90a68c9763597bf1e5ca22a70e34634d5b696ce543305a7625ddbf87ec2cf8a930ff2d397b6abbade6f9b507c6c55700d1a3eb6716699aa5cdb9b4d15b682a23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h463bbd8132d24e803b4f6ddd7833e0840bde5e56104275d86e06e2bc03876d7c2e16233d3a4b2f44a1106076ef0ebf36114781fe2dfbd127a558254fa8082d4a82bc74808da445c694a1801ef4b723bcdd49871404c44b340a2e78f20bbc0f9ca65190be3baf7521086499fd920f0c2e204a51f72e932e4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161ff5c34fa03388eeba06b2040b187bfdf59dd6ea5efef82250b98382890fa3b71860f90d27d10cce3349cc995ad8e0ef39f6bb94669d3d8cbafd131dca37a4aa21538b385528502b166708cadd301833205d06d50209cd0fe0651a7f6205bb9e0872ffce08add63df0fc13e7427e70a3711aa7ae99809c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h852c41f98352d852402ce3ed2b5331b2aa1ae7c224bfa268c3e2a0f8328308d7582e3ba51ddad476795f8f28273aa18665586496bca717189b13a527c9254fb5bda3b1c777927ca462658bb53168e2d2acaa2a935cf5012924c624126638223c9535dee59f8d96fdae986c4e0cb1c7ff60591ec1301657eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65ad7612b952fa364d3f928874f9d7da4910dcacdda72e1081e39276c29d064dacc5bb13fdf13cbf36320416223ff35e20c7867372fc95c6e2096c8f5425e3b4b8741db5ae097194d880664e76814b10dcb4c20bc541e4502bc171d71ec693d0ffcf3af0f3b14a13de48eff836297a9c94750085ab595171;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d2f845255cb623332a28c2b932cd80b14d00003ddb2c0089d7f4abc35036ee22bfbb98ac916156e1e78c84091d4c5c0ea5fabaaf6cb699e4879687f6dbafc37c13fc0fa43c99aef5be3c1f1400c99169a94fb8bdf5050d4b25d66b44f076aa471a75921e026d3a0048591f4f74732fb20d71c9405ccdf4a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d5287ebaecaed4a513dbaed04bec15cae395435a1ff02d021c5d8ff0dd8bbad3a0c43e82bcae763338d47b2fe71f3e6ceac00fcf23f426043ad8ebdc7cc9822bdb5b5931314744bb0dec6b90664c1c96c71d71891a6ef63403eb9f786d5e94a5269701903bf10a80d8849e259d7977e0b3dc5ffdc7410be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he887b2ad879dcbef45004e676369b1afc7562c4c6606bf366a8e2190eba6be0f38c8632aac773ec285199cbb06dca522a1c5ccd2b69ab3227164dcddadc7ba10514d4b482518fd0c79a43885c22ba52161cd7834f87bc87d6c75ef157b21f2139a69d058bd86596e1a15335de733a022013222ba526d7d22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ba13a7912047e49a9ab42b78b2aa89f5f9b7fc2b6ff1251181ca6f26802a6a26eab79aebc828f131762101e3c109098e29a29581101e564f1000278edfc9c45b640b12b54493a53ac644a403cc004d887035e517eb4fa654c021d20b3bc14dadc378dd471275be9ed77712577aeb9444439450a1a2cfa92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57326037ad1d5c825cfb4c2e675bf3d524928196f7d296ad491a47775ed84fcc1c138a61c4bdf1a2d4c4ab69f2d43a85f924a19e67b2df8b38983cb156df2dd4b58ac1f609e11364493832a7b44dcc7501b2988857264410e4d9c9b41c8a91bac3408c0fab423166730425fcd73fdc7c50ba409b56b0a3b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1021e4f63a3bea66177ae84ae36a18834654a937e23164b40260ba8da0c593f7c25e158fbf5229428324f4590bbd297519c05d3433db9127c40b77549d985be47f95c8dae1e9f4de35ca59960297a3a89723737fe08e23a77ca34083712083a9dc44a46709100c6db722f86a8a799202ad9b21dc6a04afd37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dc1fe1dcddfa5204ea18160be45fb2a6f314eda9919073c6a8e7feefa75679dae146399ec286cfc68b921f1f20c1b386c8332a2f00690ba86da534f9f3ba4326cca3368cf4ee2ad15ea3eb71bda54ce6bc9388ea0dd3760b666b203ad826a44188a3d0435732573da8f2f592c376ed5abab078a5e39ca99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da131afc6d93d55356c1e2f2b97fc59b0c67d73a0c1645fdc24334ed96f114927eb32708f93e750bb7d4a65e502ffb962d8edda61713ee778b1f2591b7d0a542e8af56b2347db791d1f85d6c4c6308a06a94b02086dc8c8208c49a006be10d8f955fce9ae277c8c8c5c5f4c7c3e22a734dc20b82e4435e00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6456e5d781eb176b30db1c33bfbc87ccc1292ff93f6c68e35c3b236e1f3e4aa9745bf785363f72d7a7ad21011688f50f69b945ab873afbcf45fa207f62e8667ce88fb4a9b5b77f50c14bf168392d76d3ec96443e7e2fc0a0a4fe4b5ddb2b3548df457d3b077b79e1c340dc1b948b1dacb35f1a167e44b33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c116b366dbe11c006e696e1478caa3108f27f20da8acc2244887f5a72e0e70793a2207a3bff4ef609acd93ccff2d03f6d03f6502e4b6f2a73a9b805cb0077f22aa4af2de63a5385b2181cc57f5c5da511e6185e68cc65c8814cf8a7ad4fdce26447baa7e4ffc664fb5c604aef215fb681329fe189475ba41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c64e347e77b3246c10b3d6d9299a0086689a4ba6d13e2a7c1dbb28557889eaa455df98d72fd299ab67de1eda7a55b737602461add92b4e8690a4a28bd948e4ff1ee83dd7d9657d02fe7d6685ab3d658a4d70cddc12f98b8d8d28be95d92d45cb9af7502b2f4b43694423e361b195ec19c746ff58fb3a225;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bba6579c7d8406ae9897120c42456963cb6b6c0408326a4e6b28edf5e6a1e6cb26bc8c67d979d751136e7f4ed92ce243b8e6abad69daa9c1a823f928490e858429b8a50c98de9a25d497d2e9b3dc92df5b8ad3f9da6fdd8bf9e45a7702033c69afcd0072449aee9b316fa2f8071ab566292e11737723810b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e748a621a9bf529059b952eed121e567cb34357490df471243b857051198727788dab5a41adeae35fa866b0e7dc72b0860f4153f073ed991e4dcdbc40d966d462152ec0596d3c0fd1a6cbcdbcd99a32cf15cb5fd5db36e1742f32742387e000cba17a0025af7aa86a4352e36abd1f2c81c5a2453c738c60e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef4a73e7eb99b2a66b1ac35ecc3bd02b8b0999c44ce0209782aa4a842feea47dfeed8ab2a6ab9ea885fb3557641438fd302cf4ac31afa5326f84a0c0eb5b46c1e582c64f76319ec4c7c3b40b48a9ef6ad41ab1ec959cb1d6a0af6d67e87517055607816ab2d40672c93af142c8e2b4fb55a49ce6cb5450c1;
        #1
        $finish();
    end
endmodule
