module testbench();
    reg [18:0] src0;
    reg [18:0] src1;
    reg [18:0] src2;
    reg [18:0] src3;
    reg [18:0] src4;
    reg [18:0] src5;
    reg [18:0] src6;
    reg [18:0] src7;
    reg [18:0] src8;
    reg [18:0] src9;
    reg [18:0] src10;
    reg [18:0] src11;
    reg [18:0] src12;
    reg [18:0] src13;
    reg [18:0] src14;
    reg [18:0] src15;
    reg [18:0] src16;
    reg [18:0] src17;
    reg [18:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1752ea2b38d70005e80fcf363f2b0e0046796aaa51e1c9d73177f272f979d7a8b0a227f766025ac05aca44a8c56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fb57f3337c773b3f325872fdd63d38430a82ae2cdc0b18d2e552fdcdd0228d0af22d413b95c440221dd88cca0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170b1c7351e60e44b0277e4b1393388994fcf375fd704ccba62d37a37d69f6a31a02306c89f6389ba5c8a27c2af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d06e21a9563d33ecf60e25c6570cd548af6dea79847f1d4059ac3b7cb6c3cc994fc79abbf61d398f1c2e2c6d83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1115e2499391ca91bded29d7ab76011079dd81ffbb6cbbc93624a1c29fa2003dca8fb668fa80183733969f858ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167fbbedfa6a0edd3d21e0ee3441f57841949e7e9f27cbaed5bb383074ec28d71a769509c6c2f32c2623ea7c4e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11395b763606a5df0914c526437048741301758432e65b74c95626b8bd2eadf03a2cb94d4db0297ba5fba411fd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197252042ce80a3c4f0c0850d0b45969aba73454b5ffa42617fa02621867e2f28e6f7429876a40c2c90db004184;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb3dbc56505de478506cfc34b398ad470143385f102f5f7c5e752bdec0f6afbcfaba7111bcab04b2dad983f822;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26f6e7eff450b51e763290f71c0a51ac1948595ced31329956c5a88251518aa2fe236755e02b56ba707895f84b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ce7404e03301680088366511265d708c58c15b7caeff4c277f49e6494a6de8d63cd91b0c3fbafb1ca2d4705ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181c1957f5841d3123fc4bccf640e2a12531b7dd7c8ee713a5097f73143ae9f101829c79f7d8253780f8e7ae80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24b64c121272a704193c8d7ac44644cd3f3c6257f61368da5f3248989104b7f8bf4372fb9834392fc606e0c351;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10553f980308dcb7f1f544be7721c61002be16f1ddba6177dcb37795a9ec3bb5383f6b3d009f5d28fdb7d936cba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19220888f5e143f4ebad42c6188cc3788404c8a6c1a56c41f2896c8353920b72ac48bbae734ee6b2c1e20743229;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14965b9a1b16b48b65ef28d980d18b4414ed812fcc7f69dadde77d633de389914c07713667d2f66cf43564db918;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81a38992a8b32f9316e100769bf7968f74a1a14c13c8114d928a99936828e8d7d4c38897b3dab0e437a1ef90cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9e48a813f67a792ce855e0831b6b6f092ca475ee03b2b2da242488478a7128a7b237ee6a27297cfc918d8ce50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10615f69ffb13d677a6148c3cfd0977a12f4b408aa739e1b88a7e21600a4e86074d4de491bb23402b00ea1289fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153edef6823038250f6964a379432f39eadc34b3c2944bb770fb8f76be47cf815c6b53d23ab9e228dfc9be21838;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da7ce8b26e49a80b46f18f5e0572a881cb3bafc2dc3a7ec11bb2dbc7402a5c830fce259fb5b2160ef91c371c50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7986116cefe8168d401e828d8d61b2d3dffaf8c555e19f54f739d3e2ef4fdfd94e18bbd051cd8d0df0ac6122db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb88713d254e38fd6a204ae675eff256508c231a92cefc3a50f66a7fdc4f11bc0538e212376cbf8371da767f37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5eaf4d3545a7863c903a39e8e1fbbf9da928b709901a5836753dd9db197c78aab39998f09915cb8e45b8b6052;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36dcff03c1ce07fbfc8f834e6b0409eac4ccbcfc7c9e2b19341832ab7b01f5ea9f8b5dc94e3314a001d6f933db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194870045c3e94eb3301aa5d047073bb83672ac48a67df6ec37d16729c20372c11ddc7cf3655a735aef82303a51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d2c5d774a157ddd2e11c5cae6676ca46317f859145e971bb09b55a5707bc3fac23804cf6a41321d1f0266289a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d8fe7e9f6b91d0874ff7d3be09d45db3d1b03d3b60ef68787fa40438639c28215a0c1f59416bcf728c25716a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2230c7b4f1d06c56654d2cc43b5236c2a4c46f8cbe46e3674e0922da47418867b6b3a61b7d8941439c76712835;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1639303f00183b90f2b6a0de00a0adf7addcd0dea02a1491e74673c2756db65fe49339adc23d56bad07decb2b53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17988d614f145f21e61cb0a80ca6d1ac76ad9a74bb5027da51b1bb7489037489a1fdf761d85eb183c2b6d4c060d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7558fe013fe140176ae06e447a81202c09454b7ffce14b4a66fd2c75ce0a9d38abb3c80fdb1001aa88a4c51d00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5b9b7ff05bf637f911bfc361e2dcc73a4c72a4043b2558749a134e8344b9d092ac75db134917d9317c3a8a532;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84674f78fe7b45c61d59b0bbbd7e0cb0579233ffed1728f3408dd0c60c22352f1e3cd6a542c84df713051892f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heec86723b1eef7b265c33f54fb8ef5784fee55d01a4a5b6a12babdecbc784a59ba5c3a4bd51150be1564ef2f74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c11d2431cc71b934b83ebb029b81be735bb103c4725fef808ec0e52e7f6848d5cc81c1fb772d96139effd56ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2b3e85e92beb125242b8244fb2b1c746e09eb36760702c94416010275126192f21055027a1b273642d66fa508;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h309e2945d432e52aa328389dcb4ec796811cfc08a92a8daade1bc80c7de4bd01ba69e68a5c18d247485deb8f56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fcb224ad430a4ef895c04e6b218d920cdaabfe450494090e9a55a68914ee0181f0e1db1ed5b39a84ab6b5c8dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4e1d6d4a2ebf99771529197321861b1a2666362add63fb3ffd954c9c70d404f3c7129c8c5db1d793554993dcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1539e6c6eb5cdcf40550b59912fd464d4838db33bfaa7be31dee6e29263fc81f551e9eecb2bc692fbd5c3f9e996;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ceb7b79093a848d068011fdaca804d72f6c8d34ef59132a5e7c5ce157fa812dbc3061bdc4a9a035888450ff8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30c99f4af7d3ce94e325254f9f09cc3ad9a042bfe8824f611fd4539f43e8ae0295d3b72a9ff6b961d1b29bcbc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha12e1d2245db866041e7c6a81fef31de88a0260273655bec1548b4b384d8dbe894aa8d3b194810c6b0e0f776a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85b26c78435197a18c4bf98f5e7bdb99480d9d7dec2dc2fad7edeea0921d4b5e61bf95c70b5ef270c370fc075d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ea0fbe5f12494c3ae196033de9c82d9a0f134dbf0f9aeafa17999c65f340c13c9e931154eb8da8489244f5818;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa9164d312b52de296c3da46850acd0ad1e1659ffb6573d7e67632f740f8820ebe0833acb8731543a8136ff05a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h217cb01599299957d9629f17972cf236e56d11239b9b7725fcd5fef486e10a99f8a0499305d34eea1e0e8c8403;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e4be56a237040568589c80a8c66bb6009a23a3aa548a67be4f559452aad3ac3166434682d8f7a189e16da659a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20b8b74718815ca0d067afb9ce0be8e971dc219e87823f66eefddd4944a008a89d888222075def5a1d69d71595;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141ffdc10013a19d2df9c3275baa441a6b223727d48283b6b2838e1d1af30a6cc784be81d1b6ea7f2f14f474537;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107bac78933a3fe835d92ffb14e54f86035012275d58cc64c5ec69f764aa2db6798aea0bcf65e8dcce24599e506;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105a999c48d40813b7fdd3b73f92d158f6d2f621c9e71a3b952b0a356349001119f8ef68a382bfc7584817d201d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3f4b1a3bf04399815bde4a2dd0a9a12b6c36f0e04c79c6b516a6d4ac74ceb3cfb01db411c0f11fd1ccac4913f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ecd797833d276177560e5e5c1583e575c7e72caf3797196ff0ad0421daba8c5e1d227d6116f42ca86e85511e03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5d0d842e12a9ca155bb870f1c588c30ad150b7caa1a1e671bb3d9e0a8d5261cb1b096ede7e478da049f9742a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1232df27265a9e3ccbd986883572a31d3204154ff01d619251f0c735672a645b856c547abf497cfd9dc351a2aa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a40bbea28fa75241ad0b14924f6891abdddacaa79533da9881f90d2d3bc3c0ad428547dc72d860caae6845c63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1650568e396b8ca0b4ef1f664e7cc3365a5554517a6fc3ee8581b0241bd2a73118fcadf2715a797bd3a76cb67ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1900511397fea4e364fabd9c64610024dcd6eb7c5d0849e5584458e29a5769cab8baa3e7cba6cb5557bd5595c1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e216c40088611809991d347f778e94000b3ebb3b531a75792ca58f776bef3c6a192bb9b566bd7d8921e01350ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa6d79337dcc3406cdd4c8ac56cc729f25c187ce19ec056638f7c1565b0309f5bdf8723484cfcf1e95a5ddb372;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f680a0982714da2b111400047fcdad6bb6ca0b0b39cd4a7509433e3fde9844ff78aa990c8815aa49f80910a271;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a48ba88a4ced1b4223694ca599f4f1f346cd5187edb59da6dfe194796a673e7f880d37297f332a1d84df2659f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h799b712de4239ba38e17b963ecc0cf77f6be2ef6758b9bab6d6e4dfc36cf41a45b5c24938026a32b6e0eebfd98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4dc315ed430d3edb65d2984f524a293a97f367920edae346d16d0c7fa4a57da8f3bc6143de2eaeb0b1256f1546;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1deccdb78fcfead3e3ec3a38ab105fed49424792998ed05aa32188472ffc71234c18d5b648986dab6e651cf13e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d31cb0e30cc5d6470f4211d03c80534a473661492475ba0b5908dfcde1fe9c0cc7f4e687bb48dde4108bc68b6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3af479726260c0164b751fa28453be6a2a12aac1e8ba4ffdce913fdc4aecbd30a252f3379b3e2fc2ae3afd91f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fbfa89ce25b2150ab056366e0ddeb7542e063356085db948315daea16548556db7c954875ef954f1578fc2217;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57f27c65a96a6667a4326126484cc9af20cb39b37d0f81b16218594a7da6a8e1f57982b3f49a6df08374efaaee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaafad8e23a725725971f187a70a5b9f24f36ec24b4c9ec8c9242da2902bf5fc3b3a278793d7f3884e6b558ffa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37cc5539dcb025506bdf78c7be5cb9f8af5f8f518095f67d9ea09b41b0ac06feb1272ff6d9799e8edab1d3fba4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2cc201ce458c05ef439ac0c5694bfabaed4fdb1c6deacd183fba48f9caed93485b8631c66ba3df137b5355aba0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fdf9a0b7cb47c1b23ba2cf365fd3ee2129cfcde7a0e5d57f1e990cfaa05d1923a820097994927073c6caf8683a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ce79ce634c3d5132430207ba3ee5218ca08a81b0fbc4d03dcd9e39d0d1e64406bf4f1ccf741941062196996d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91c9744841d00ef38f3e457cdc59f996f8316e7702b03bfdf6c0525fbc766226bc045f3fd4751dbd637bbf9749;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a79d2bfa116146f26788a5caf47ddada74d4ee60d20425e70815446496af5f891003ac46c0cd18ab8a23c315f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbce2e6a29028f58789db13bc3cda508944b151f4db3a8e6ac4baecc546be57df3fc589d8fd1d3d53636335d46b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c8293e39386c33e1bca6cd9942e8fc197bf541ab1aa5025b57b24de2fb7d66d03bd5781a0ce945228af92baa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cba278ffff4b13128ddc9b995d1b0722881ad71ec84d4761a79eec09701a24135f613bb5a3c6a878d538f1e72c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1429763bd0ce7ad9e1399e1fa864ab28e3aba5b556b3dac68a825c6f9b587a00bb678702d329d4d3f1ac6684c67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193d67e7b27c50040969539a6b32c3389022e4c4c5f06674b67beaf1814cc6cbb20b7d83810a47cddaa2d54d635;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heddfd2ec150966b8238be1f407e2963233e76c30152e836aa5e74a470152807e13c97a996268988eabdd8b28a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cd20f3880f5aa8b716a9acbbef2f136ca3c6f386f1b06a3d56b27d35b32c2f8add968d78bd8a07fde14e83d73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43d0b73efc858adc14c6403157e2951d36362a5970bae3560e74e737ff2d5e3aa2be3de14bbead81ae14210f4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h673350f2b288942483186f4194003a19724c11c66a0a8b79b3debc4482da35666f8905b2626cf3f54c732dae25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37ed88273a631a3cf720c50299dd468d4462f2dc6ce08fe5f2e77895964c704bc685410e5ebbed1a18a443c953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18acf85f9520faa2f41fa2a05a77e801f558fba5cf579f81c34f4418984fbf7107e7581d8509a449555ce2d66d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afe89f2fe6eba3a6c7f02b40116b9416fdda6aeffb131597df98fa72e95e6d384f3bce1d375d8093dd7c5be6d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19997e29d78ea38107aaaf2412f6b6e9f3204751e22d9ad3c9a73314a3a8cd8e5280b30a0707f8c256fcfa70027;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h84378f00e399fa9ad64c9bfab7e07c012f3e8ff7d036e55e4c530f9941ede25167d99ea90e8ccdfb2d0cfd702b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dcb2788ad35279745d50d114e39a0059a2039340f30421746b6978779bf54beb41f0c46ee7e9c864279736dd4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2fe0f6d3d191c7989a212c4a8c44aeaf66e4dacbeb9ae6f63aefb33c04bd7b62099b814223fb0cc382257c366;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h861ca2210d609400c0d9f89722c2284a1bc0ba9f0f8dbc6cfce0f9ea102ccb48b631adc99166137641487c4832;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4299c55d882acf64ecd73a4c2ea356219daf7ede955deb696bccbfcf5f2e968730f43496fad0e27166843a8669;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a977b830ec8dc9c987290979016378b848a19d5262b0d5c3c7ca8e01cab232098e6d2c99ddc248ae3a7cb1558;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9827b63fe42e41988b48e887d728ae4079b04d27485d86111a8c7e7ebad487b2dafed7ceb93085718579c3e6d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbebed2ad72683ee021c23225af6b7d4280bc4e1af6f9010f02d5a95ef57112a843fcd57ddc1e9612b7ace0076b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5b8b7d55d701995b90b1f73cbb57c3f03c991ef08488b387698d01600fc5a7f4499a35d7ec8230721f9dcf26c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c23f1bbec3979dd6986e543aac13fd4be297672fd830d8564210f58fadf1eace343463666f6d7072d103de4fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29ed4a260af5f649a70f88195a90ba2c14d69ee33649b24714701aa394a20b37e911567a6efc901f2ae81d84ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178e48f476d08b3cd015d84f45dfe44cd2f7502efb91dd3964ad4292b8ce6fe2b0d4a6b1e678b52d52c01345dd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h710ded40b17b2cd61e8dcb294322f0f36b5c04488bf246eb54bd3fa1751e9a5231e56b5dcb817048ef1d295515;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11845f9ad770f244048ead34df881a070ef33ed7bcfb6edf20c0ba4ccc7156a1c794d0893d53dee4ffbfc1c1adc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1c0a6a79a950fe2d92bc306c6f5016415ff9b86cb26d5f0202baf7f52d759fce384c75675ca4e6e9f57fa9334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h950ee1edd4fa60e1128c9e2e92eaf2eac472e91777da826ef8284cdb866d0242836fa2a218754b238b1c43f353;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bd58072fd71664a5844fe4a94c91579e7267afda583d9de8f8261df03430b91ac2a451d8fc6c5802ee7f464a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7eb6c03258747c55afb085926fc3f0c8dd284c157c695e88257248cdca9f79a55b9d7d72765165991cc72078a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb025a256c5a5fb37ff5fe72b0295a3a33da75ce70089e5d74f50dca736576b9e000419dfb2b31d00c6fa47d1c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81ee53cadff9d85d28e06e9da350d4c81da52a27eeb6f6b09a9abbed7bcede69a00c37f12cd09015fa9ac27b85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c6f00954e53c5b8955615fe05753abcc4ca248f935a1dba21782b1e78c932db83fe76ad8c51de3be78a122246;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4a2f04ded608c2af8a2ccac0eb725c19699dc808976b5c5cf4b10fd3cbfc06cd136f9696c8cd1059b0619b782;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8dd3df4bb4e620def24f9514af93200bb369e94ac8395d4fb5e327380a1874f49f5db1e663e94ebd7c64e22c5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d43f4edf28d15602f27ccbca25a0b2845285bce6bb28eb3a824c64e21edc95aa833076414aec569b8d3d96f1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc6037f1370d370949eb948cc63a197f958f7fd273e427828e4b3dbaec962383f72b52121ab3949a9e4ef0479f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a734b0c2e355462bcc071827c21eb04fd52768481b19e93530be0b61cb85de94fe192b815de85d66e2c5b0a88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaf78a30deebe0c1376986368416ddc6de19ebc2e6694fc17a7a0b784bd663c2a024b0369d32bb86ba495b072e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h821a3a9747e13c70e271d6697b8e6f02a28ecd6b7023cc10cdbcac60f97b114f187dce19fe8d9d6b76f47c5abd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4707897edc9ad5fca8c16c6d6056a118d5e574a7757e24db9ff93fcc244a8972d9ae1131b45299db158705690c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1847706a350f495eda835faaedf5d4ad1014b7b47fcc3b179ebc910cfd753de838b1bb849cfa796aacbb56cf7e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h557381b2a3c4d8c6536c5430c98e89fe4900d33e246c65408794e2dc99222051d0afa917c8012b8d8df79d9b76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a627327ecd62ef4c9562e7530a74ce6c7eb9695895722c6028f3f31d575034fe9dfca4e1454a20f87b2e136b0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc0601f0351c0ccb5b02af1a0a8843d7a4948d0681162e9463fad2aaa70672add6064ef17490ebe9ffae243160;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15de593132b2b6681b83500e3c75ad20af10d674b0c3bac2fe1ef5247c73df1bf9ff1ea7905583b2f2ef28d8148;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb8da6379648dac6c1a9c01fca7f698089736ba38c9b80498c410e7b905ad8b3c6974daba1aa7f535a85a670eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h216f9770ac7cabf57ec6cd94ebcf76c2eb9c7403308870a019b0bc41b9c3bfb17472ebafe35e79787badfb871f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c8867b7d1259e1cee57b1fa4ec5a3dfdcfb5c2ae2c5a5ff6d10d87a84075b20282cf56ccc3fa2e80da432b0fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a4ef44dab5fd99060ab75e29e4c16e1684eb05fdede44e9e9d3d87d34c3e2e5df6a7c3a5b1355121a14ba834b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c789ca59b1f028d9baafe6831d050122be92c9b202d984df891b5e5d3c5bd0bbf70f995ad69d471ac22cec28a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4aca7333c6bb733b4c6b5be43f64a91047bdfff34f9eba98e2eae10c5cd677067024b998846349f34a5f5763ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf54f9cc6abec8df783b93a448540fdf5273aaa222f2384d922183f2b1ebcca03722a27b3f829082ff68088486e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19993c31f2fd7c7f201b8a412dc661505304312840d66181cf14c4e244b71427a345e285e871bf88f2f2470b953;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5d5c95ceaa652e060ae241ccc6373a66a9d3357630d9e8474dba4341c9833a27f309598f5da554718f4673057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc128b6d2831b69fece491b5379d89a48546e9c016a46c0387a07347fcecccf2893a24cfbe76f4d10e0a0a5aef5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2b0746b257e4fcfa581c80af22693b8cff5dc0079ff03049eaa793011e49460de177453561a7c1aa80edc9526;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192d12f21f348b5185fef1ba46895c9cd72ffcabfa09db7ca9a65c997a7ade01472c3495abd6bd67ffcca33b7e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3602854977b1ef6998613f2897c57d3f99bff79d4005cffa51a7d8f8c3723958b113e917861df694c82fa3f3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a125e54d17d4e5b6d1dbdafc4a4ff325965d080642e20c323bf8a29ebffa3e68b9490a9c2015a6c9c970b195a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d356a4721fa170f9bf7baaabc7277e2fe79b235e1bb90596e57afe3dbdc37e64ad25ee4e3407301f317520a950;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dcb056432e58e2e159fa602363959cf9f7e622867d5df7c59a5c8fe0561b841a330ae61e99572075704550e436;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f8e19e1ef5376a6c8fcd93d7ebb6c102dc3b643a06b607cb918fb17b2724c8523209bd8750af55d284f195cb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1efe214b99dc582e9e045ac6f449546eaeb643633d98d2263a002ae0ba646f8377f6b38a35b438e7b4fc4cb418c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d328fde2b100c3b4c1b24fc2f2299fc3e0b131fca777b9c1b7b0a2a0eb0df66a4df568190004d90bf6a8c53fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16642e107a2d5c6a5491099edd83955cdbb85720e9e6efc5ab8b4634eab052d28dc1929d639061196e6be97bd33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10cfd2efd0f0d35fa4a56b15a972b79898ac2f36b8a525667a6cf4429def3e8db20a0f8f6d87b573f189239e217;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c3a8a2dd0f0a813c2b40915ba3d2bfd8d89ee07265fd0d1d44cbe89d72ebed0ed9be2f7edef5e7707569e3c85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c399cc9041eae65af2680285b6c86520abd5c6e42ed2245e85978f806a3b7c96c4c4dbe15b8a77e82cd71dae9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c4defda01e540956dd8d983fe21316064ffe738a44ac037476fd28c5cc0fdd6eb29b4277cc532edcc7532eb758;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7acb1c262fdb9b76760c1254a5c7a458a959cc62bc643f62e902c46a881b2de39fb77817466ea5c0c42039493;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4738bba96896e8f1f55d669035a72d82653ec9116dd5e50be72bc8a19d48b804e20e5790920f291ddc15b641e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a285b78d1c0a260868a68d45ad6af0b7edf644030a36f4d7498237495db0c387b2faad12a445616daba20f2b25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68ee2608ce9252869dfb3e5f0524ba01fd54fd202a88f187d215976c5ed0b3f770695c0dc87cb2660a84342f1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd4f38ea0b10eaaf8ebc0114f02d0fa4ee36070f5ac7f1869a2afb4400cd9ae7e390f727d0e8dfc459dd6171c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h884f82ba31eecd7727e66bca82bb53080f9d531770733383f206a4ed22ed017c1e2fc5c670f499d8f079c90cd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e93d4fc4b5146aa134b39dbd09fc8e7e2eeff034b5a3c4db1b813957984c3c68a6e82d8c7391aa9d9a6939366b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1983eae6ec6fee7e62cb57294d6527f39d5b92dab022d8650622019a56ebb538d25c972f8d0ba2e15a634bad9b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30e9dace0a1ed29e34fdf2a2513ab53348d6575b1117e20e3aa34593d1a51d4b58eae5a05341ae48ade375d3ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9f4722115949a2a6accc1ceccd26ac312773c02b7435d0be68ae4f62bb344586ca710373e115aec965c5d5714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1905d2c7b2940ecfcf0ed807fda6a5d98469c8b5224785bb9c41be73347e4d347ad7fc8ca1784beb5a7cb665ba0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb0f23bcf431a1624990b5bf22a87b1f8b5aded8e1dec5f016a3ad3f7a55bc56a70871aa39b93459a67aea3b44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b968529a8e5f1bc170b38b6a72ab73e607ba5db00655bd32a9269cc68375cd78dae1e0d75c475ee1ee3cedd8d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb59462a4371b38154565854f4c88b60a9a28df5b898779322c873d692aa04fc9af53ec802acbca4d5e08f36c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110c24453dfe897b3b7d617a75e0a7f835ce89447ca53507ec6a92892c204c0e48c37106becca09dbd15b4c9967;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5107f3706def56c805444d705490c568f1bf06e09a2e0516d253f84b036c35f753666399d40b6ddb900dac7702;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h820645d46fe575edc0a721ee8fb77c12705f6a2bbff6ae63f22e3e72612c2acf3c9a495078512e417cc7f61340;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h388e95e033739ad6d502ef36f86cd31e91626172838a79ebf9ebfd5684f205c8246dd811e18fa0020e1d5a8d5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a98bbeaff8820af9ed53d64d2e8d500ebd8f27f955f16c620d82b0443f877e87792654db8cf8c6b3c6c27232b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e67c7f24f34ae957af0ea2c94e43ada63b37f824f741c9c2780011d3620e05fe2deb34ae1084849f2e99f31516;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fc1674f74cd7d7c31e9ba110c77f2a94e9b41385e0ce32de37932f6beffc318da34108cc6298890ab7fc620f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f61e8e363f015336fabf36fe47c220c95d3b11498319e951c67daacc3858576f2f906df9c30d35afd26899001b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23c4909f7aac7b882f5cf4177bd96ce9a708a43cb9c303e4d8b566ae15750ef4fdd92dd40a306bce5d7f03897d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha00c8e38f6c1870ef5908f9400b327ac3866335b6af84d9287a10aa59e8cdb31470e65d62e848ef677471ca994;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1903492bd9451fc048a6a1d83e612f3ad0bb057a56be094f6e7a2b6fc5e9c254748866547292ee701f6b7f1d031;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha787caf83235d1ed346a2727d94a0b10235827f27a8f9094bb02c6cc0e5e408ce63f3bb0d393daeb7e2e03d05d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7feed34bbb4c0930433e0234b595d3559a3735019ac0c742c70384d3e0d4206e0050703c7d2cc7b5b613d281a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186ca7bdc910bd6fbb40b1412cb03d5c87ef6099b4726e84df2c7ce985ac30152672f10a2c509c5be58a72b3218;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1492869c0488702b4956c539c03db387f628f2360dba90d2f40b30187281e8f2fb9b4e76a1bc6150780984e1e63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h221c1d09eeb6d1b5890d73e37a1247bf7d9dc2a65e48b64aab9e3a57a93b1e7554fda8f5511dbd1f564bcfca8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114d9543297fff8392a5e39d7d8a124c853a69c87e3558fabae7b170bacbfa27cb071b85bde8382e569d927115c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbdb9f69bcb096ef1b58fac539b9b17fb7e6bcf28167d4cebed543cebe1c07d54b6e8f62d0d628edc273122d27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1bbd97d84f020f046d77e1b11b4341b3bfffddd617d06c7b7707dae0bfa202a2761a11cd686bb5e01b880a935;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c00c70ec1c20839ac36fecbe6a5d3b5135efcb90658997f70a5f0881c0efd4486ec51c7f6e690774a7fcfda5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4972858619131b44c58ba59438e162ed24ec99b6bcba8617d3ce645675a926bf41fae7360f4e21ea27b88ebfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b641c8cb88dbf6aaae28de22554eb218c249f23598faa08b7888994120c2e804fba45032d0e7e896f78dbd3352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd6be7c2967ee304b91223dcf7b6bead73e07bbe0594c6645fc30b81f5bf350d817e0ef2fd6dacf256a2aa2c01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he19cc58d3162e8eef629e9ee3985687de26b754c4974714682b1d37838b82bda3127c44684aea8510edeedaf67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56142ce0ac0088d8b8f32e2fb8ea692d1962663266d1f7381d19eac6ef29d6e3b5470d12f1e038f27b05b28f78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0e318e9e1a6321d5bf2fe74d2c13d69320bcf1f3d78fedc036a925ea5247229e33fcac82bf9fdb3303a52deef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he39ca454b95e76ace67db707aeab41ba643bc2b6a50ae7359090db9806d6e742f1f09476cc2b4771226ac2358;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f929dc8a92ab2c327cc253f7abcd06aa2a8e49ced9b0128d8df1c24b952e66d7e3d3b432861b156f0f2abb2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29bd9b58753d8685a3de09dd5128ea483588b2180aad29468781d853149e2475fbfb4873a830db9ba526c6e1c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86d0c5b7a60d511c35f24e106c220d92c48ebe22615ca299638c8caa27724e9c1cf1ca28a34f2be54aec5bfde1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65e35dbce39dc70059b0f6b9e8cc1c12423c90f7e17daf8d2877e2bf170ff90167e4e4744ceda7f53d4bf643e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5797be22e124339ab127c835614f5794a951f9a27320255476f15699f4cbe362e67b4a22116bf4deb8a0477f8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c92daacc73fc1a0a37ad056d5b84898a5a8389ace0ace2bcffdaf2ca2b566ff0229c7d76dc885fbde073b3303a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdcdc21381c4501406d246f049b64c182851b10185229fa58b58cee54f119a81f1cd7f2ab67c43ea781a47a53b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18cc63c6b81ebe5e0af56bc3f8fa4db062d764de29dbce3b3dfc4d4d4331184cb36380384bfd425a2af811990e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106b13bf0fafd3190bbe478538f1ec2e0a851afe23c79eab3e963a5f7b4f3d9bd449408e855eb8efa2f3dbca848;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99e2cda53b9f88a7aeb9ee206e1713517023a3dcf65385ae2d32a2fda45e0f147860cf86037c52b65a72b02240;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e07c643444cdbb810288cd2afd44dcff1cc9638fd3b7383e999f597595e66e499871388a75499db64f0bb096c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f663d065292a83540a3f61858af34ef2b92ebe9bdde143888545abc83af809d1e8c28fafcf844816813035363;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d49b07b916a2ed02e0df714b35de054afc587b92d01e15669d288520d4edf5a509bf7d202ec58929a7ba77288;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5da0f67a269be59badb721e813b71261c98b926b3f99aba732890426e8e40407a9b97513acb809296173679721;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90a802efb21250427cb6d442045cb383f27b052f21bec95795e77cdb4c6bb55636abc7fa9a3798206e57998321;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3820b71d3e2aaf96d338e6284ff536d1b5861a63eff1005de1013f35235d408504be92e361e0e3493c03cb7c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52ad4024255a0d6920452a7524427e043ffd69e3ce4ec599845cb655479890830d1ec1fb1b18c9546aae264c18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c4898186a4927ae97de3c64c876511e3c8280fdc3d804263cef5bb578ebcda552fa1f7cf0a18b9d9d9f5bdaff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d14e5acb5a1fbaeff47411556e829ee37a7485a4e0ade639dcca045bc23e849dd2f0ad2a2c49731ed23c1253d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3a10d0d901d8eaf864c3bf8e1952948e37acb3af4ff45649073cc16690d9409baec346207d2e36c8dd28bc22e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5e158cfac457a359090aa7d0d0d2a93df44f7cb93223fcd37ec65aa24b2a5357fb17e4b0808ea16d55377f3de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5760996a1f0ca81d529dacf784394cf148079b237130ca6a185bcce298dde92d1e394a9f4c71927dc114acff0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h663aace7ff64f55f0fc60e2c9b54bbe7564d7d2877d8cbf256235b83be2799901470a1b3077fd800ad2cac8e7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd13de5f93ea5e648ebe7c01bb8ab500d5a6b2fe5dde627d7770d64cc05383e7d2215130304b41d8f7cf945680;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e571423beb667d8d5a9740b92f398706b211e29d12e89313e8a93c385d5d5a25c0d68fdd3e0e96e34b25771b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69408711da478e50a203744cfb4864cd1b14bb01115e5f6e3a818cde5c1fbbd9b2b1bca7d80814502532bdc760;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3b90d85febf10324b6439b14f142665c7e336bbff5e7fe037eb9ec636ddccf2b8b4c936e151201db2edd23105;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36f29c5540981f033af936b9ed8fb98c5eafef418cd858247702959f9a678dc602b23075e0ead03dd28cee1126;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba85958cafca70736a2a821f3ad5a92d5ecbca751528efb3453cb8645cfdd3ed39bd9b058fcdf8ffe0d373d218;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117da8f7a8bc8d50b03eaff9982434f182469ff7947f40d1010f31d9e5571e96e0414970bfed104e4b014acc3fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f84d7f73f78ab84b5c0241bcee565446d2cd260b01db61c6f78677378d4648916c3c869f5a63008c69e504f665;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bab848fc4e680879e5569134c1ec823244726d92481e20a38c43ff4f5b4c2488918458d93d367983d4d027a00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aef63a8d6e4f77b54e364a90b8c74117a4e91b9558009bb795bdd3f6bda492bef6c10ce3049c3556c121103d0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebaef187011c2ff2bbcf2344ac97245fbe5e747917bd7839adf57eb1e0caefbd13fde979d4f329fbc31d1c92b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bffc87d85a31f9303fc6cd63d34eba926c668dcd2bcdcee2863109db555bc8c12b8ce69e69546cd57c7818d6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5522456fcb464f5f860c4ddfd6f68402e33f4a3fee9a761becc75482fe880ee1ee5992b09b39f1fdb45df09b83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af8026279938aaa92c6f205a2b634e89a7070fd298017639e4d3c9853d47ae106f9604f0a9d7df577a98b1d507;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55717846b1e851f61bac40bcdfde56cd393ead620c2b3783ba175749fa850f43cafc19274bc1d774ac421f5d92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h394e51dfd88a245de1af2be3b49b5d8a17d104a5a95af55b65eaf6491e29c650fea5041182b9d0f7b863bb3428;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7848f53f15b949e2ce2a0e7f37beb8075a2f7cb587aafd126088dd483774f357e7253d7ce4d01366b212ff6d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77b88b89131122a44f73a5d6b55e4eb4249aab39d81e6ae519cd9e1eb5ae1a4ae016e3e0a1070fe992c733d36a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb18276d1605e7431d08d8c7a280ffac4eac3d05e3b76c33705f35da1a8f99f251685a6e8fd126e61fdb4e90f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ae1207ff4cee655dff84e5e931e2a01a45d5902a228a451b869ff457bd0932c0cd10b305fc16617550e65a3ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf88a335e249788d0797c4600a50893c33754b16212bf005211b99a7341234bf5bfbc95f84a476a962a06bf431;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9467c19d6512cb3696f6071d3770aa6b3c8104fdbbc69c51a2208c0a9e43d6a1e03e30a115fe61192cda326d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b54546ccf99dcee117039592c07be8c64d62346b8a4ca3d84feea9bd9df991d41493cd407184fea381a2b64c61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18172e0eec2cd765e1f776402724e86455364cdfb9d8fdc0206805a3aed5203de1ead8999385393548ad2b2677c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15659b7f608d42f5416558a6d39e2a8069a2e1e41b68200503cd61b31ef24c489f800f06be0cb6df3999d107105;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha88a0aad5004e880ad4ed17d6787b6aee3d2cdc25365a31a0b09052764d1fdafa4d26384205fbc742e271bf76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h255252e780fffe4f0c2cc2e3d6bfcd3e231d3cf97408994aac10f3876b5028013a2b926ed7daf261a15f8129ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37926cb7bd3261b9900df31bf5f20ac86c1b42f2b1cabc875925dfeaa8e88128bd0e49b86e4fa568f00adc5a75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb9475990766e58513348d84cdd190123145317d40e0ee598443d7c75978d2a844fa74f9bdb82ee73f73da262;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e55011ba50c1176a66525964391a880a1a5311ca9f19e80f9ebdbf0b2152967f93c56412467e7cf7c542c01422;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4551d64eca66cbd82dc7a2ef564bde34d2ee7ddec8d2c21619418b6cbc6a3d1532082c6b775eaf308ba23f25d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86521563c9d1393c43e942098072db38cfdc18023aa9fb8efd170870c06d0fe60d87d86762f86e6b7581749c36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7029087777aa74221bbc6c364d6775ad96e4c18992fc8c7ff26ff57310a592a70dc0d069b77352db10f47d4b05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1214c1f78841bc4c065c5d57cfd21dc47a1b43374f4d74feb021dbab98b306b3aa0a060302ded8fd34b751aa6ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf36db943499c270944ab75f70c748d978bb5959dca29bd10279c6d7751e45a6cf526eddc60d07e2ca2458dc2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ce4b8f9871ae9cb4347a2de490f2b850827df48399981bf6f66fd7d2b59135bb28c373bd7c8139583955d4cfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cff196d53e3a040d9721535e182c59b55a6cb4fe171988f3ae2d999ddbe3b71a648b5ef1b2ed0c1dcebe5b9af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164b093792dd24db71548b6b8d1b29385b1ba74f4e35cfc9bb2ad31e323b1aac4fe863b948b18d64a243e9beade;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9326fe7dcabdcb329c307fdf478111c8435c43701c6f7e41a7f579167a2b3e2c81217b99ba8dd0482477af2e62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1647347186e8140667da9165876c105deb2b2ff661c7bc1a78d7010c397b08013d3802adf1a08eaab23885669a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1632a2703476638b551eb623c8360402e3c84cc17ad9c94f76966493d79f94518b4edf74e87203adeab6fa195f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h916525084c448468b8b08fe8983d7a9ea271e5a1cd697edd43bfb86d29e0be59d6b1a86dc710672c22f474503f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3b3ce1c93ddf8ab4e5c201a280c6c8c96b91fb8972ba614e518d2b86126651c827a004d00386863ba158464df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eb7cff51c63873a69f895471497f9066515d96f0889008b573781cd334ebbe690139bfc9bdf77de78a3107d6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e55f351a3acfc77a7360a802227b92c8dc2b423f84e97ba0a605e0f8d2990214332dad340632c7e854b3928845;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8af33b1e49372b3ee95593529d88eb74df1cea866ba84e0e10771cb0d9206ba0e6826f8b37f7b794f59ec8e086;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba1d6f6e0b050f488e6a3721123ede45a0631edf5cbc74f661fe4fc1a24694bec339d40a30c36812c23869933a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11da6b51f5b55c9e69db5d38ba1740cf271769398ed76f971910a7e12a67e1ca12034b25820327c0daf78ea8b43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1167223b76325fe7e84a9e50a78a55a93e32fa659780df6c2c5ee3e0c2f92c83fcd5b399e4efbf4077965d0bc44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165edf71188a8a8e4c671293ccead93606a848b203b47affc49b19e0fd124cc21ea845e3da6dd3a3b380a95becc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd23441e6b6146a68f420411dba6a6af46f35b937a3ad96f2c66632104901dd4a1189a32c58ab41b1e9f5acb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12122cc682ff32b794b7667fb020d474f00ff085c3abe9221a7e0e761c177c776ff2adbfacc29f1f5593bcc818e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc90acdeefbd1f39a8c5c25912f455b0bd0a472f981b8059f67aeac1c33009d53d9dbece2d04d26cda08c68b155;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f5b43d08fa0cf3cc65c05985a09761afbd5fc26627244ffa5498792b7719df6581706003c8174ea8650575351;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af98dae8ec99b6f9588555234a0ee63dd684d632afa16bfece34dfe5dd78f2ba6ef20cc4bc43208e543e80405e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90364351c8cb44bbd6c8b4b4e2b9c625be55c1baea4118e3458ece402863c6460ad7d8f61131cb76b0c5e66784;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127243b53b048a15a6cb47a045e7cb93dc213bd725c1350a4e9e0ec4cf18cfcc26809a34554cf7d94d0f59d0dd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bea3431e53a064fae9b0291eb533cd6fc7ae11ee921b442e3ab2bd50d90eab44054d482be74080076e91144c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97331f93f646f11f10206971871f8ff4f8fbe874f39e32799393b52e3185a56a574f70c2c1a5ff424e57819878;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fe2f4a551fbbf185e5dcaa0155051312adba898615505476ad4dfbf06a2af86141172b422069bcae91d8b421b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1210fa9eabe4c5f47d5fbc18b4c11717f7d12a8073db5b11c60706faf16f477c7cb4f20122db8fc1dcdeb37a9d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h826b4758e74873dd67843f72fd7e7b8c77bed0c8f1abdd0546d01bf72678afa6cf390cd9d3f1b4039129dd2911;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1195aa38b3c26ce986d454396d191783ba26968007fda8230844f82691812fdab24f5bfe1447abbc47214ee53de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3460988a9ce0752acc6072b5c2215a26af7e85f0428328b3e8ba60c8d5ad2d011817ab6f50bbead23e4ac5023;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5df86bde788db8def116ddaf91a1f182aeb0fdf701fae4f97c323e9d32837213b0de8bd560dbc822e5df9d263;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h760be3929ec12807a98be5ce13859178d22014ffc8d69353664b29ab83be86e0c54201ec46ed39c5531b7a763e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf06572f6c9afb0e4531c49f982a23a417d401a525f47a4ab21f68f6f9035efdb5b514e4e19987c0cbb9c5f5041;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h483fca0af03b5c7f6d0826079afe9794cc224490f693993d3219db6bf609fd2bbeebdb03a8a9b73f57e5113f4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ca601140d4178e404ad915f78bc7f0ce63803707d1bc4cdfb4aa15e1b48ebd3b9522e6c77df6d3b1d0b39ae96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6e3729564351997a06f753a61993a809167969cb43ec66b8bf819459465cc8e22aba553e5e6e853d9ac598135;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e7979e0dfd7826cb80b03bcf364b9d9f9a5ae3a59023396f9e2e3c2d4850130ee9658b78f4d3feb6c5f9303c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1043ea68e1b0cba73d13b4a29c5137181774711ca115ec5905a8182eae535073cf0d6bff2a7f1fa163c972e2410;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176ddf4056a4a1f3bf41228144dc1b205ea1e0f400a7bfc2c85d9d6df5c5223dd0b72c64c0056b9121ca7d26989;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf847d84b59ac7d1e715e5d165afccc84d7311799ae681aeb3c517d7d50eaeff0c3dd5852becb45a88d91a8575c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h283092a5c83dff6ceb99432916bb1bba0fd473002f3b8188b6ede2b6c6c3dbb86722582e7d8bf27600bfdfed96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e98237fb23117021fc13301e977eafda6470ee7212deac5d0d55e63780042c3c06d8fa6e04f05f04942778023e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf41e97427389e0991e41da3fbcc8dd067439eb6a146e22638ed0875b56277b197a06ab01b0c7e26681e9241c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7de9d6fd0678e9b4edfff7cbe1fde24fb4aab8472275f2b4b6c4de5b479ef0e08511a8eeda09e75521dded3c5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1751c96a897494e394fcf65abe5ff8aba9135055820c101d85cfcf6954d8d234166b1c628c0cbc41a22536714f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c26ba46f2eeec67f1c7cc4b6637718f15211b9909e9f8f52d5a048726f63ef42d32f1c29d47f7260bf3eafaf20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a596b40466a1f3c92b3dc059a5de751b67fe492fc4f948eac1b175d2e8ecd4d5e4e85c2b0576119205c5d7c9b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1537b39aedc7f4301694e5d8bd5e80755270308fd34a2eb1d3ebd10b4a18e358212062223da75203096d002de86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h354ddbb51e753afe6c2c4ab4e66bfbab93b2bce240551b8b8edf9a7c7aa819215f63a5757ef85c6cbf4ba55c9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc409ee4f4a8f7b75491c28b64632a5ce678471e79a5f0ded57015f3149b17de4b2c28bbbead3c1f14bf102aaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a86e41139475cdeff88a2795706b757218d53fb92850c158a1f27180c64bdd0c63a9b8ac143a3612d406f78871;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h207c17a44722c2ce124162f042c711eec007996412ab3efa2123c5ca61a688af4acac3a602e130782595b6ee08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fb65c836652e086e637d7506af889e38aa62b84052e2b474ebb300e169644f84c01a5fae40ead236b2e4d03aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ab104bfc4c2895e74f846006f855c2b6e3a7e52650855ca843bf43091f461b0b7852213d80b650eb47af2355d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha152bbbf2df2f02f9de40078e611a3357a6ec8840e129dd9b02defccde24940ffd4800fdf617111e1648b46af3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e94426a911d16605e0dc8f6a79b4e4c1b903ae3585b94e9fda5dd0a49dbd3db49f5370d28ccc65764e9152488f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a6de84a4dab74268158f097a3d987f9c1912305b4c96b65982fe6cd48b9da48a1dd919885acd7a3ea87ccbc57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce1c2814f767eb7ea7b1c179fbbf4bfb9ac5f77ee321882f91d59e485c129e81d38a78332fedbbc1ae4313d22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e240a5bdb7721711417015b8f4a1c7c25299b5fe0830dbc7f72743ce2565e5bf39546e6aa43b69623f4cf621ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f980ff15d2908629e2ab579203b4baf471f34527a1cc4f5e985e4dae46cfd06dae7a30329af5c72e414203217a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1659f3c00987932a703bc5e16ec79ccf3e7cfad2a0222b08abb014a867647815582754c673ef7f599f90312fed0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2406dc889470daa3e0782131cdd7198f7f579b0a9797f299a96884134004ca6853d21bf81da4367e28e84dacd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189fef65842735f29dfd51970f19311717e8e1680be624aa27efc8b41c383731027b670db2fde06b15dbf59ad1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97c21e7fe26c0cffeeb1e316fa4c7e02ba8d01026de22995240ccac4dca7c44ea7f0fdf7b19dd867ec3cb12334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4387e00753c930e72c09fc74f39d369f3f88095e851e41ec71aa5661843f2e110f96df3ca631328330581a0258;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h398a2135e5b96190f55258bd4b7f15ed0d182d4c72b8c02306e62dde724927f5cf0bc48f699bfe10bc9b5e1c2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2e54d47fa0e58af16b6f5d1aaa57e0a6c34087eb54190976dfc18b392968728c7537b7a61563973fbf0d05037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db0f09cec71da2b58fcf2cfea4fdccb1c58c9fc06226c2861310673ef487bacf234fb9ba7253b4320aed917d64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17aa5324ef12fad15f56347c6858eda3ceeae11eb5c71d7319641b674a48a237aeb5eb02388c99971d99d942a8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bb9be4d14b3eea0f830c3ba0b0d6b26ff1e73cbfe3bd6910f4e9102f4fbbbb8abee77cf914f8a3557733b5238;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95f2d4f8e68cce1edc43d0b5c0312e59e498bd4ac6b66004b5b7c6f0a185e41c83edededa749162e0ff1af8ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31ca1e3ff99150b92fcefa60410d7c682a399c94a0084e6f5923aa3c317877d492eb1e0155d6cb0f027b4eeeda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed9e05dce01a037c5686b4a96767b52dda12d81054be0a6bd00a85a05d7a957f6b119968806d5d49da8528c59d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfc7d2382db16062520435a7c2da11efe8f7df1207023d4b23a26c5eebfc5730dd7b76b58f2c825eefb62f4233;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188ac76761f8e62a36a0ca062cb0ae2eca4d525d42201e8b3662449613f45acd6937ee1394b86ea159daa6d9920;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1efeab6b930242dc950f6b01bd2e0ab441d6f31dac59f308167b2f2209fd9a2b6306399ab54d97d36c77fa5a477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df64a7548827e967ac2ff6dac452f21270e52ffc5a2d34d847c5f284b0e4c3241c1e0b57a771f5ad137d668341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b5358544175e3dd4f6c22dcedb005549034bab1b88df6f60ff10b62b1c3adcae784f7cc9da7871724e114ca40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b51fb4e6a3425cae7130da34e4b89fa3738e46daf2f15606dae905353e9ab83999e2553068c68092b7f16e9d99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138c6447e782271afede799435ab49f7a003f6f100a9c884fe636e7d272a12b8aabf92c66296aa3801175226360;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5f25f4dcc8100686e1bbb8bda2bb24c1e43232c678629e01a1df5f68fdb26ffc627d87e51c6512f6da1dad5c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7caba70541ca3201c6109ee1f3b8afdad9ece86ebcdf09189c143622685d4a8eba3a882a0fcf86af3c214479f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1684ca4165b4630ae303043d9c0194e56094796086add40e2ac7c199ade56a900a2d4909971d7ff6c0c9d00809a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6dfe874872185cafcf1e94f3559d4868a7d06a9996d95df2a658e33e00023b203abb7aeb40a8e41de2cf96df93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7567c84b93605d7f7cb328cabdc0a19113fa6c471929b4de6ca3d1215640ece93ccec465a671406ec2afabfdb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7c198c741b53f01a2f9e39da2715ad5b0ed1b352fdea0722207b8c0389abf75ce21523ac493aa7da72f792a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c195158a5a94da4d6032ca7dd5aeba50bcb38267ea6c7f9db2f1a71fb623ed788cd2e6d1522547a6b6b28c9dfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd514f1f917431ffde91d1c45472b33dbf7ac0b9d42ea1ba9222f7fb889c71f4424cec9d9594a2633447aa419ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5fffab2597dcfe24664dc22547255bee2c719b71657ed484bbca45b916b727635c301ca6698fee8004b5835d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99ef17871b03f5d20d313999e6fb2844f2b21fbe7f75daf2355ecabfc6ed72a75ec77480bc37cb54bb733f5b14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe4206024a014814804721f6dbae668e411045cfb184833dc3d7628964cc267f98c4e70803f02742e7334100fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h56f0109f967a21a7c8cf302a5773bff29b9e887d278c13961a6ef896ef660dcd1f3492455ef9f4368e327fa97f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e763df91666e94b26c2a0b6a36b72708ba84c7a0c4f063304e5498b5cdd3b03e089b0da507f8429e31bcd581;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h458be4510931d9ea5a053f53c675f009308d37a3b4ca3f9009975cf9f537cfa5236567d1a1e3e9e71e9102211a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156532005593aff5e7b4d4d30f659cbfcaa624aafbbbd17e8a4089e3a4b9b072de3e124b1b8289dbc4c04524eec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c0773b8a0890362981a5c5f9197f97d0b725d51f97e64278595562a0279c9c709e84a53b78bf361fff613b48a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c4f87949574e15f52df8008f98fa9e976214534b9cf99bb3a03a0acc6329eb3481b2d4eb0daa25c4e3263b1c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4396b076a1a1372a38bf10ff5b111244fbbb102749e6336ad4c629cdea76b006309eacdcb35bbe6d778ea4914d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3734064e48ae8305ecdbddda988c7fde8ff6600eb7dba684bf46fa7e21f351e465e9c3a357dd994ae29b1f3c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bd0cecf355883e1ced43a28368b40f237362a72c89d0ed62b41a2ae6f62401998b5e837dc460a2f0b5928f058;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6cc98d79b9bd9e772f8ace0a35ba69eed8fccc379486b4ce62ea9f7d06fc9b381aaae5d189397e0f9621c7d17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71da2d0c7d63ab5f1fd501bfaac8a3bcd965bdc62e36a2ad65a25a6a6712a30d4729b2a3dcb76b8ce410f5a8ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61f58209ebe870130ed3e382813276ef528aa6b517ade1b359a0691dfc560282da4ecc98b4a3f445dcc62b1b1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d43982f4c34a3f3b167c52aa78f1ea240688f5199981de8d11d9a0c5923b40ff00d17381d81eb2676c32d5e0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h307bbd6dfad50c4980c07379e6d4ecc1909bfa5e94717333ba7029d92faa2af273e23a6e81accae0155052d986;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h410ce2dce680f7e4837e5cdd98f69d2514777e2b8c01070e1fabc4774d0304645d4ab14a810304620c5fd26b20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h208b6e921f2997ab906635585319b4e14e652596b7ef23ae269863c3921567e7157092f27367ccc4556b3c01b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9122e32f69ac4e8f9ba4db6fb62e5e3c690341fa7c56f5bee9191156cc13852f2ddcc45888d5049bad9df61d9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c20b8b4ec4e02ba9a4c99e1dfe14535b418cd48518c320de32f73c64d660e6cc04329e06b1782a4dd75e88400;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f38ee346a7bffe2e9f4a41266385ebf440a825a8245549022e0f722cf93db4227d06901c8b4526767ee6d7143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28dd3cb7ccf755cebbf53231a00857ebea391e7cdc4b13f094c40cf582775661bd8a5294f40edb98735190b151;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1958887a5a4e5a69cd43e9f07ff91f759ff4b8830780258cdabbe9fc71c8b585f069052c0e81ab800807dcb3334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197b28bf19c95e302dce92385952aa0fe321f88267a15b9a122f74e5a068dd86a905dbd086cf5f4c94112e9bdb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193ece8639c6671eaea603a21de3f7baefc7e35beeaab45cda4fb125fd9e8d88402bf7d813135dc5f21c8630427;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f089b1744a8085510b270154ca90c876d88b782ab2b9046fd99c6fd488b275422c9a05200c99d4d190f176b203;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b54e9be7b6642a1348bb0d4ef77182715bc81b168260b21b5651218f990b799cc5bb4543864076596fa59295f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99216ba3104399911cfa4a3cee8fb0c9c7fe882b8b781317d7e39680a3cd8bd7af7a24e1069d0b6bae7ad8e228;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122718b4d7993bed3f1d67f159cfafb16cfdda56bc0a9d3b02bc47f66bac97158913c9efc3c6436b2b97831b6ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a6a93b6b79d0e02be73ff77ed47f8b1372afccf1a621c768a03589d1419eb04bea5476c06e48a32a1035337f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd3e9fc4b3bc9b92b8767854f4efb58a99d2e04f601d643afba0f87dfcbfcc7c3baf301c368c3075681e8777a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he763340f883cc2c945dd0c61103394f7eda10de0f192e98d614ceae7cf84b78996aec88681668889404b685694;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h976f8c8d91d9509432754c7ed2fe033b905ac034e7f054622026bca5fb73e4ebe4ed64fe82e18254274d39660a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1272d4d42408f40ac15a039d62c4e86c9bf37ad4df759f2ea77b7a30ebeeadbc13e7d2369a11a1f3c604adbbe03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137729ee3d8317aba78a42001cb0a60c2d6413f7dd67f90eec356e0cb2f6cb20f1ef9e94acce605d2f8a948c50e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h666302e5ebe6f051995e5054ad372debf80877719559e99cf239f5db05b41a212bf129c5c7d684653c357cdd31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a87ae95e3497bdcb5de8db94933865a56150de3073609fd0327c4a334baa42f4472865dbf52b86f85bed6b340d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175fe2851c8134670dd18b171dfb8c7f579c5cd8bbe91597dcfeb099262e919296e25cfe0c0fcd6f5155bdae88a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74125fad09849df182e6048fbaff0a72c2ac30b2474dd0b0eacfeeb0aa8e9cd320236c2722750093c905076bb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ddd5d65dfe38eff4373ae63229355f2b6e315d2cd0f5c89812a8e2fc55f2a38bb7584bc59e7c71d1f57a81d8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d82313b947d4bac0a5f9680fc853d832c803527cd0681fd09bde60ab7ed1767258c686c41a3945f40b812c26c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb61d7ff4fd989b6cbcca9ca48e42ac7e51ca4c094d34ddc50ab1e91496ff8252bc33c771691e612b3534a88e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15dc1ecf52d63a833ac0bdd93bc6908dbc4d0fa6bccb15d5e8d2ede82d8e7c0b3c6fa0003f6cdd86fdf23b05243;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde873fc8240948a883e9bc86f5ed06baddfdd883f2514f5ee5d2c8934ce9723c67d30c092239b4cd2c6ade3a2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d1a9aaebd76f323fa2710a8441c01e040bec0f4ade004b1401dbb298edbb17de5a38b60ed64b1732073f47155;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104a27297255caa1066bfd631324a4a84dc703370df701f880db3d89cf644f47d1decb1c7c79d04f9dee8845d20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12059be558605c591e31f7e8084856baca3553cf59c1140507bec01549d9cc800865000000b8be9cfbf1a4a1011;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c96d0b27779671e560e5db646941eca666b22faf93a7fd0acbb907ebe1fa172f917a01db688cc24e224a3a4e1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1f829e95e2597d18d8dfa7aa82c48d0a5cfefcdfd4985e7c3c533eb073274f452226c95c615caadab13e10029;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d29e556ee062c5a3a63a1823589baff1a72cf6fbc8e562f8c2009e96cbd30ddf785711c1f379ce8239d501856;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfde1b1df2daf15547cba59ebb0aaf878b6e4958d477b650e3c18bde367a5ce7ea8f69207c6b1ac3bac9beb8d41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d7ecc420c901d41bf57d78ac264f7a53a68acefcc1a832199cad104a00110961ee3e5998d5a901e0319fb3a23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bba14a0464f35c339523d29ab0c12db9c114bf2060501c4be4a76626c1f468f6177e98ff91b45d3e6b62d6c155;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1631b2299c04b7771ef383764b96d90e2a2f6957d02c79b3864ddc7a2c5e24bc1d7526f78f0d9347105d90f55ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hddc8ba6b477ad14f4f77f45e1808ba28e42e909b2b609445c6c42ce87fd40eb1813d4df91def6cfe86820745cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e148f984e6f0caadc05d1013d17f714bcc875a86cafbf83af1685a14676a204932b3ae5e1bdb7af662a35585b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196ab4ab77118168654ec14e45f93f779dd218f031e8a4e1836c59be5a5041b20eb739ef9b0641b57184100b3cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccd3ffa449167570112149e7e1af4d926c3a478d72c616ce0eea8a04ebc24a13861a96a3c01a31a46811adaf34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h666576acf493bcea132e5b84d4f0f2902a5f8f3493e8df47f449f0270e2f6e2553fc539e62c367225ab3f2d1a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1547badb0cb9d9b8eb2ee56197bab70595b1284d5666f8610f1c75a8c4df0259c876c2620554b00f54659ac32d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4d05e3af78bd32a2d274989744fd3198a28f10e2e7e2587f2744c3b032d0f803dd2b88bb7db4b5f96ccdf6037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d83b573193018b748893b1d7f754a554508c60eea821979201618bd5a448227ab5261d1d85ae7b7225b2bd4f3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e767954764ae8ebd1ae5b7b9b823082512577abd5b41f8b132602958f08c6933e78b57e951da2a3fbadaa392c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94396002ea8924c771db5469eab884057a80408ddbc9ccc7b4f38a5a4736f70dcde38cacf9a492f762fe7e47f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75df222ce93d7dad5910239b69d4f0c76fdfb17d71b9b9abf7105cd69e0f80291632ae99a9a62daec29fe81456;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h903ba23913ddde020d5afef5254ce85f7e478b11d199d638487cd6752ee83465311431f790c4bc5454402fb4e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97b35e5e940a3f2f279039d0f77c9bec2df8c459f151b5081f9d579ad8510c838b825c0c5d35c49a1adebbcc80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34e6343cfb392ed942f70437ce245ec7f2db30023cc99b12ca67884c4188899c4df100f9bfd609d5b0673a5eb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4175f5fa0513b7ae992dadd2eb804fb9b5d95eeddb5d932b91fc9fce71c6544963364d1233a014e478d0c1c756;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99fd1ef3d616a2f691455809d68e6362fb2343fe876e45ed902142be73f9fd64e48e523f932c4a072c92014e34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc79ee818d23b3866ad6a240602b60c242f09732bbebdc4e2da680f1a119115ff2c70f10ab0fd12bce56eb6c67f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d40ddab8436cc70fa0a3f07dec9727fb5d1e7167dd4bd3cfca7d041a20f3a5f8c2018b368e3b88c042e2b8abc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb38e289848ee47853c524f158461c0fe9743bbcba2418d8981a33135fcb1e52b4d2514f48a2233cc2ea17e3208;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdef3819e1e1b1addbd426fb36e4f7ebd5295e3b1fd991562b619eb4de4124d4ebaa82cee501b5f528f0b1dceed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f83d707954dfb2cfdc325a3c8274c35a0ef64b3a6ff5d399d0882417310b39ea84f07a2d3f357f972e9578446;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10cb38aff13c96bc8e85cd53320c0e67e32bcf3f3af18cc21372273a75ba396eb7390407895d02a1b0f7415cb9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8e39e0d013b49bcca526525d518d9d52b1bf70dbdef4c689bbad99c694bf1a9bc7c9672f2b31256792ef995d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4786a7194dba7864360c20ee78763b3de930d30630e1f915dd3934678b12957f45e4448fa39d3a05ea47578ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c50f8e17abce97b232160b6759f7b6ef69fdc8e19b953d572fa13cb61ee7dd9e11870622692f6d7c5f8088d5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1877aff311ca550ab9072b25c4c5fd86b7c471209f4abe06af83e19f3708d79e409c0e7344b9877968fbff72cbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87a9bfbe2af95b5416c198ff8703dc162517f87ce2b226cfc36689cc6edf888330a2e2f6c9fab6ccfaa130bc66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had314a577ff3fa18f6d6a9f0d5a92c85fdf661074e1a5639dbe8003a3a32141ec269343e4e16861138d4780b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h501597a3bbd923b16a94b4f4bf2c07f29b5ea2ba1f917759778abfaaf795c0a236dadb67fd5f203837669de6be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecce3036dd403f7b9347b358fb9470946c64a3356109726239df6b590908b9e6cf5655797494b10c4e66898ded;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3bd6e890fa4fed1d3bc19a64d1846c58e54153306b54f54f86a872d43fbc1a72be8e16906d6e9ebc15853544;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e044a7395dcba06c996ce256b88df901029ffff483c870de877b4e51fb6f21bced008716ab62df0a5634ecd11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1322d279df3f1695edbb687e8c16a4556cf71aa8c7261bd060d08c50005260cafca84fb57eec9ff6221e38e6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fe2151111532e00e70bbaa222f01a8f326778045eb0b03d071c59ce330e503f23c50410da601b1cf10cee70f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a5c542eb3b4a80ee9318d964dc8a4412acbf84e7cadab83b4ff4ca837745b5ebc168833c72f30ee902549ead23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc10b2605e36e5bc278f8d1c6854a8dce4f16697976738d2a263fcd9231c4ca2901eeee5571cbd76f0521fc8b45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5be9cc5293e65362f7361131e077c8b72d38205043fba09ee021f86a75849ba3f10ce40354703bca22b9180914;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172cce9eb1460c53b95debd4d685f7dac71fd96f0a1c1121f360462cc8f437b4c4b7fb2c8dbd96aba9b7c3a5c2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a7d6d456d05bcfa6b125dd99f9f8ff80e5ba2e3b5cf80dca314822c57fb9dd9ab49a8edae228326dc5c77a20c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6eb3b5c70c5174c0db4b5f79e9afcc0de0ba7e3afe2f1b94b3d94969a63c7cf34fbd4e6bc4f926b932ddec5841;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19253cae754cf000112162d2821632d023f84130de30f6a10117811b2221b72946ff925391fe2da14886b2e5648;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd8b9b75f4e3c282cc6acaccca0088156af72dfcb800322dc4afe75c3cdd95a45c086072b8bd21867fe99506941;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fa2dd6ae4c3d8fd2d5473fa15457475b01805d65ace98d66d6e5ebbedb91ec381e055049ba3b15a0a50cf76b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc793ddd9b618761a43b5ace53c190e376f0a5e9d95ca0604a9bb84a28113df84e603f507aa75a1f032979e016;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59ceacef67497e47ff7de3fa1a18ad774c63896e3ff0761e1110bdfb3ebb4bf3e6d9b740fd6c92a65f2e2f7c23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e5cc8b7375498c67abdbb4e7b27abd21b8d588c435e61374df284f7c9763057d220436eed7c57f2754636ff0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc51f3919ac06674e8880deec271f391141a72b207be485d2c5ed7034ac719ca7a147f66010270a0333990415c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf0de26cfc9a358c714c3b12cc3eedd74a2b8ba103d4fa6410306dcf0f3f3caec9585a3ae67060a65d39aa2904;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c0aeff8b1e5304f55a944ae334e2c5366cea76ec6e87ac8e360d9fed261eafa519b594843028b9cc680d68843;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1622028238dfa5b96a2a24c4784367894207409710e55fae7391e45ddad87cc4673bb18d28b30eaed01ccb98c80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fc9323af0f1c5e1c6d63c79baafb5d6f448dbbfe8b0fe3024a3221143df7496feea64a599b65d42c948f470f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1995fc0afdfbcfdcd8402047535daa845d4ab4f7e7fccd5d57e1d27b34146817cc4f3cb7a94ddc97f7a80ecf329;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f702481929a82dc561430fce72ac62177ae760d0f28f809b6fd11fe05ea6dbd3c23355168bdd1a99b30df22171;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14391a7cd034c9dae3b2cb42de12883cf9271bc836320505f56ddb696189a9d7a7e59ef81eb4c4d5c78698f05d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f47f7105fefd72ad0195de2f36c9a0619a1153b5cc295dd385b68a31e6cf8b7b9ad35779cbf07957ee368988d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13916910a7ed0f72f1d4ff79ebdf82b1e912c8ab3627dbd8e76b6e87311358c7132c9f4f6c84ef37b2a486ace83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d41e55ee959bb92ebf88d18ef9b44e5d8f13315ba72bc70414cf32a8e52e0a81aa8cd00eacb31a0e3f17fcfc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b52f6f029c041e033adb24c8ca138bbb252d6d9d1975700bbd16baf0565f825cb4ae0a28a74b24de7deada1e1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ea6431bf20f762967360982464901eeb31251661192810496a2a5c8994aed02a715f42386d96bf9cde89f3cca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6f1637d8bf26a4ad602513a8d2c217f25bcbe0e3ddcf75004ecdc99ab8c9763b83764444a67463965ecda0029;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h367e1b26208b8566d525a61492d09e7f8f2cf036816448fe1e05e7f01e3a2e6207e6a9a9ab4e50fdf5e8430bd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db543660f3cdffe0b2e147cf7d5e70153522f5e5ab07dfe39e34acb43de82d9b707da53049651880c59c07dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7bcabd68a2b73e57a2ec9c27471b05970fe9bccc0cd1d742fe872b5f3cb323f9db769cbf737e3cb5855456be0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172e7dcd441e394fe289d8598d27703e19277209e4820192913e2547edc9f3cb9c23b435698dd8bccb8a38bcfe8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55406140dde11b6ae89b5c8983207926b74627fa9dc4e88a2f676f2b76583ca93eabf725196d57d3a7f8c09774;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ea89d7db2b27b35a27339c268da3abe58a6975b3df35b2fa97d102d05aa294cc5d48ad5f4c322d5ef0fcc32da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13edf44ebca73bf69b35501d437716e88e8845a0c36ddf4a9c1c4f31376a52ee43419b5ab0d7cd8c45a4ed1852e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfdc09e72e92c17a7350d068118ae9fa23f6e54eca9e4e549fa676c91f850f122be70a15b0bf1ad334e09bb196;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7a5c894e3f34da07d59ac267b6328a4449d9766ddc79cae013164389dcde65f75a5ce65446bcc7358e40aa00c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75173160d5d3d70f73bd2d3fa5fa99ad9a6b5d1b7d7e0e82d53026c608123ab063ade48ef5ad9333724dbda978;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14571ab0669f97bd1cab98a2ee6e71d78bb5665d94a87ac031bfa5bcc5f4e9cd1270bc69139e5ac6c84c54ff917;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d291d84d63b99b6140e27b7934b803482d922e08afde0ed6a786f9a777930e1838af9847fbfc708ac5c6519784;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172a5d5d116d28a265879fc38d021dfe5fac198b7dbad527bf7ed0fd4dada98911a7fa273677026b01dd365b688;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d48e7e847c6c95ea6c85a9f92dc66f9fd998d96988fb4f3ce6843a1b9ea5b5a20bbe4c044b03ec87335c091006;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h87cc26d4d8b32885efbcb33705e85a00deac8b058c517871ee012276c899212516455f33ba6220023b569a0257;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c8c9c59c75e70f722b947fdf61f716e5fea48ca4ee0cf4feda7583e47fab23e659f4d4c15bfcd5192489ec15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h913e858bdbf7c22235e825685e255cb19a92aac18a2bed94a0a04e5c0dc9b0b63375a5610b6497a0694e5bb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116dcffef592a3136fbfdfafb034bd5fc4a42bc4017a5c4514d5d2176e925332bc21b985592529ed3cd89dd372a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h519387eb04e047086cbbd2e53c714017084cb45000cd460b2391d151a7ad927f0614592c406d9560f7ed45ac6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1becde7731f70157f7a4a8db3f0417ee7f42d07112df10f2b5fc74bbd4a0faa0990f673907944a52d2994577ac6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c7765ec1eec6b67f6fde25f487a7d7d9726bd05453a69ff3e4dc4ff6cbfd4e5ed6448da20c72e4582be5447e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2ada983b1c13ce52d1dd5b3c01ab93c9ca78dc0925b7535c9cfd5ec34f53c177539310028ca269995d0ac05c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156bf82821e7e6382fcce25e3743608949fd6191da569b781559e4e315f2a14b29d90c1b2a8edc4cb0ebf5e3f7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2950c92e58552f0ac60d584a7ff5ad5dbdef1d227bb60a328e6b7438359df198559dae667c0996d7616c7627e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfdd60b3d8d01542e5e545088edc1f9d95b690679e05ebe39f25e1faed4466313dbaade69c2e29c2060739b0b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179cf2da39ff22ee4c26887f1cc0e047aefe7468f36f4d1b461a155be8fb941127cb0592e4932a1ddbcd1b3d322;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa1ba1e5a4c010c58bd8d437f51792723fcd55534843d1ff40ff3908373cc3580dd14415aa91166df4fd66634e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c712bcef0230f204b9a25cb40fca11f1ad536210659ace0acfd4c9522fdb564e0f0d6d0442f5c7f880558476;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c695f469a7e6005656622c9e727ffb71bc4ec56769ef85430d8cadccb6998a5372c76cec5924461c89876f3dcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6f7188eac1dae13fec7ff0766763c03991b02a961e7f8380f2b0884c67a9440a7fef13522a092890a162b5f83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ab3e1a9b3a736478ee3218b8ad1981c64b999debe191a543ced137df740e2a8c912a4d5ce702f84c057715523;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he991a687f82cd86bd521e979f9e29ac53f1dba6118e8728077eb35de4771d4c46b76adaaa04cfa497b3627188c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1114d5882dbe25e5c096a06c49f7f634d5e0e48064dd67cf3f4d3762b08f8c88c2e26d2fe383a7ef228c2b5f1b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152528a2fd42c395dbe97404b89bf2971436c30190d06c72153e24918ada84c00fcfdd0f13253063b201ada191f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he769f915c73f9264955d7a7dfcc5cb49047aba432ab6b64120880c4ba0ddb708d310f0f47b9cd0a6e65bd7a6ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b348f72eab25966b005c553d79d7692ac5b53c10d7ebf51c6f1b449fc661aab13db1032318520d9056a3692cdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h157a7570b9e1022b68d7e88d050dd0c42bf261bee6d2127d0cf22967fca96d0af107c85fe80c94e135cbff9c152;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b74656af895a2c5a1fd97e3e0e6a45cd74ffbe0bb1c8b8f6aa8a60bff77886f5b665f0d9cafaf39d63c871a52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h896f2ff5ffe7fac5ba33560b3fba266be5428f9982972cb42e74b43566f5ff19d136e585ada3b6acea6a9b41ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1289f7cbe6b3e152f6f3995bb6e494194870659ee2b9c379ce00bef2da619fec0b53502c4f1607e4f3c1e52a3e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7341a59005a54188d253510b4abf49aac19651ce5e1b499a99e10ad4be616a90c06d489841b60e98c0d35c84e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc5d7659c493576b1740782460f9f3a0569f384e68e744919a759ebecc5d52a1140abfc2604828af831f994f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19710f302675d3d505474eb67755933a41ddcb2318a06cef5782ffae040f8e817707dc27c641557131a1834d684;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d01e9c956d3a2467c6df2e4f9119467b5cca08883806cc63867bb3c5489e8e6ba48688944a282430b45923cb12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f062496f1a54fa96668789e34a00e39c39417c0055d891c23eab2091f32f875aed40e6c88eb672f9b76556761;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42ede42975a0cef93a14ab84e85e272cd4c468e128cc5f0e634c275961ceb98fe2483245376bdb3907f9b9793;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1058d8fe382e2558d4effbfcef707f7122be1021fadde0dabae6b2b419ab9bb904f884bb4950577656c9d626011;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc79f3b40a01485cd9d834f159d5dfddc7a1c0590e2cb0078b653847a086ab53449b571dd1265dfd404bf0e6e91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5123800578f5fcbe355613cfabfa25f285863f78240d018f77d7fecaf1a8e325d4d57def04ac6d5387d42911cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha209ba36a961c131906db1751208e54d9012d7dfb9339323766f8e7ab9896da50eaa303936c8fdfb1c4a9da99a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104ed153ec08578e52c788c7d4e8d43d420623ee636112ab33828de77484e76cd7acd6a513f174a3c3fdc07665;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7ed185e9b3f87443999b4494844e0391cd41374b519387f8145a17695e57a96b5a85d9ffe792273cd593df73b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1431bfb75c71f7475ef34c32d881f7ba76e010d911217f84f6e45314f8c1fc6d779c97371e4f3bcbba17be0857;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1974986d137cb9295f301669699c4a23cc67c0a9f02eabca44ebc4527e7a75d671e4d9b15dabe98456dae210656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155313c51ac592a535b9e2a5a553a3b24380308f84f9a43212427051dd6ea4292de0999ff03be4b38c5b6f72d53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h375862b9438a1c007f44fcb7b039cfdeb41d9bfe7dcfb4bee25aee4bb780a84f6f403a4edfee49d733c13aee4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a8b8e0d1de144a53f719b6041c81d505040042a6f7497a65f85e48e5e17fab35e2f52b637aca11e17e35be8d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34d0a867800883c81c2593c8457d099a51420a7b2ff579ea997fe816bb022898439ab257c87c161e56defa21ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54f3e63081a3a5837aa84a93923056b3f8c3f694a2e676968864840188b6d4e38a5897f24bde604a3a6698bdfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd51104ad59d55e00a5bcb309c67e7d3ba40b2392a35a43074514d4a35647bee3fe5cea6aa76da07d54b75dfde3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef49eb11d85827e3042f37055eccb214716aa857b0f9a74b2cb0ec15849e588115df6ff32d1c8a8514b753bf87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1f30329b17b95f979fbea59b6c344bca9b490f30405452ad4ad076d2953ee01e86090845bd90f39305acbc062;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114c4476107379d427ed5c8971bcd04c0e26f71a63754be09066200606f77d44585c31b7e9c7be33d5aa863a740;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b739a139f25d53fc0420fc674a888f9ed9eb13b0ea001affe53944a2db688c63d27c2a34c1279affbc059f9325;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138fb2e6920324ff0950bb21fffce28552c8e079b80f1d56fcd8c1be971bc10ac2d58ae077e5ccb52c7e43d5f1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb08b8e86ff183906a3970ad78e86c026e2ef97220441f986c04408bbcafaecb579e5f4340a6607656806148230;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf07d12d19f02a91e5ff11b1bb0389a71626ccf072909146db43363a2e107796aab4d88a556f209e0dcb9d2f2af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h702326d9219e3525403a8f0465a421d198d06c15ca87234d680093de41a2ba3bdfe18c55f815f2204fade32b63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he767eb615d945f4b8a316a8cdf52fc31175e4b89277ed54393422d09186871a3317da937d71a8838b704b4029c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ff64ca6b10250e3b334a3bfc2bc9d35c4cace1fa6ee550eff0690128298ef7b39a7c231fafc4a4ea20ba451ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf84d37ca5343e5cd54d61e1789ab0d5bd8bac5c3c018511f0bc65a2387ad237dbf8fe5f47a1f7410f8c504882b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h157aab9380819dcd9eed1f2de88509be3dab6bb70692ac21d1cd6a782ae30df22293fc4bc30b36123bfb8339b1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1feeeb02f1388df422535ff4037a9b775f71409b7062da2d630d4e218a60b280ab4fc2b709f4ed7422f1555c414;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125cb70aba57ff4bae95df8568b6a6f8668d38eca7b7bd5c929ee818e256fb1e88ff28e33b2b75b2ed22788bf71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7409e1c26d37366032c52348950662b80ca513fb1887848001b06b519c0c43d96f28e44713abac396e26150aa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42c1fc2a34d5208f36383b548dc9168deeff87854ee69baaa1dbf3d974223e9dc8913ba6dfa32bb69414033673;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha21b213572ee9738c6f64e6e17917cf4ed16bde4b426fb0b5ace4162c5be372a0fb87f9db74bfc1aa14c10a209;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103daafd56cc33597b5c25df3a12a214082e7a39f1478d04b8e3079f0b99ad276842f417f6103f5dc8077d7fbb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf263bfbbc07ae17d809fa8c60c801bb73cb1d8dd2536985ef5cf689e622d3210d8649930bf740e75d1c2554a47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa4640a51c5ad999fa4f3f75e28d43a6b7f8b6b85e6f5907581cba6e73fc42fb4d36e36d66915ebf4ff9f2b4fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14570acc8f279b82371bd6d9ae9c54b3923740634b299e55d379f2197f48895ecc7b74148cd9a61df9072d369d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0da1f550f564b492e74afde46aec614f84b0d30ed2578d27a00c6df0e3393d290ad5d5035224c7c0c989e1b3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19410666d2ce9ae4bbc62e53669f9b936e396edc07036f9b3786d3ad54b1c1b260dcd297b19de0cc4c0d6af15a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165aec9e1a632a31ca383cf601712bde0c4adf8a1f067504a96887af478825acaf7601c73ccc640f1c749ade14c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb4bfaaccc35db941c4a9c6d45f0b2c7647fae9a597a5f8ed1a222fb512218510ecd9f6ec181703ee36ca9f5ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1270d5712cd2e0a0b598f05dc5a477d13199b4cdefa0eb0fc5b492825473cf82aee24d5c03736973e4fcad5de2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5945f45f1060d2269019417e1b95adb95d1416a25c02b74a15f4b9271afd793b24ad3d335bedb0bb0c59877b27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a9ebb94d3d0cb12eaebfa56d14392c9ea126ccda0d25eba1ab4f5883526b4eb3e66aea9f6907dfab344855d01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0d103beb340a31dae5ad99c4fe2053947500bcfa70a801b78719f40fe9e6908b92a287c623d8a8171305315f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c482b262d50d7d15970a707e60040f84ff98fbac12eaca3087b5b7b033b5efffdedbff8a8c7b41c957fa84593;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f55ddf4a98c1b76e6c7928931f139a5ab1879aac7dbde44fd2c813ddb244b8a7e07dcc1c521e8108105954f540;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8f18e5bb6d4d14fa6598994b447be5190dab3f495e7d0cf0ab6be7c811980472450c5b930733cd43f0658217;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ab4b0ec20c532d644aa9525b07a05ce92a708fae92df4bbca85e8c350a9b1abf1c7912fa6e820dc5b2debfdb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d6c80e64efc559972bdf794ecc3eacff440f22819756b8bbab17a2aa56f193ada895cfd9fdd3ce06cf4bb135d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4f3bea461d92de042e07a8682d4f7cd0c8cc7990ae0a89c7f195d7a2e8f4d8b352c8f9bc70712ceee09a63c73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d76d28d86186e702c50388ca0534b441a17ab30675950234198135530abbc85ed90e5c31cd58eeb2bf082aa0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104b347ad8f0095b32248e014a8fe4e22f4e432060ce5459387436c5027d837ef335d641db283693f000ece9e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a155051c07b85dc50a2c9f9345fc0a91f2947506f9fc59bcbcd66de0ae03b666e91fa6c0bb9d924139ebecf733;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed33d8d28f09fa74b2a6fae987c8ad07cc665306f57ca8f5719ed541ecb626c039ad4386c5d57f4f0c193e6205;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197a98211ff82adb4af15614f88c86b50873b9586766154a7c0a5a0c7963c3c9d49ce3433f61ebca739f3f617b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134cb68bb8643190ab7788a5ff03588fcced312522254082e3caaf406184593f6c00ad0e92c05b58630f6e80a4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb94e5dc956dfe1c5ecedb6cead91f8483fb6388ef8cde8347017f48a3625477bc260d407e2354ee87f48f8f74a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f7bc8f8aa19ed42fb64a9afe7456a6e6b84d341ff0038bb178e80b36d3557aa2960482f8fbf254ea06436ebf3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h865d5373f2258d8f428742a2c78fc3d2daf52b4c26c9194c3e3db59e2485e563626263a9e8b8fbaabc35f4768e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1455d3d8556cc34ce02b423f39e56f62b4471c889652245269e4c00bf4f545785d7258b73b24507896760518d4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b03aa6b30e34602ef53f93ede40a2603b71e5650bbbdc5402f4cfcf85f2db55742982026982b4a11c028d318ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19446e7aeeeb726dd288adf0b647b98e17423074e8d1902389112093c2a6a6656734709368a00225f9f7ce55fab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3613766d0911fc0c1e72333d3a955541d9f8cb67a8df267e0eeec6abcd108aa0f22c94c2d4e0ccfc40cc746e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e00c15e3394150939e6a18d8cae9033a448453b28715a60bea7628729bd611baa6dc0e9df595203f061a04f9a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf442e57fdf658b2711e9e431393abc57e46f04319a0c6badf51bc740c2ae86ea020c36768444a80cd3fc3a10b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45a283f8396619f8612b68af6685156c05b4577e949b4253c3108d1ac3744ffc5c8dbebd6b89b6ac179a676f60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1652e5eb44d39f0616502d9e99201e2ebb28997ec276d00e7d6206169fc3c0ee9411e5f29bbcc1f0e12ccaaef1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h378597fe817e7f4032cea2a53785c7ad78745be65b452e1b8367d43fd3aee3076191ae7bf49940ba02bc01c32f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haad04c3ebe8420c1dd508d3fb7dfd84fbf937e2efca2310e3d770c5a4e0e6187ddf0f23b852ccaf65e46ae80a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61a2afac0be8a6174e5ea0b033d4d4da54f54c54b016fb97d040cd2276cb44f74f2e30e7044a46794f87dd18ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b9b097d8116836df6f0275d6b202052233d2fda4b442a11bd30670a8df85bd01a491c7a44cec854ffa3c0cfbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75d9d755d1f9b934a64b63d954a6b5456ef8344961829d3cc3188684b8ab1a41c4eb3a62b0d9603d2b5776656c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd7d2246960d3fc65b207dd66e4868e7e9068a692660b8508a699a677ef84dfdb264fcd3a26966d44f975116a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8a1ef31e4473d0f545d48d2b2dec139dc752abc0cc741c98fee746e3fef6115d5a7e3c1906d98251dbc0420ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba16afa05f87f977037edef0231774720c622fbb4efbe6866097fe45d1ce680b53b7a750cc8beb121e2571b08f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1952fde7a2d712ad510a23d076ea202f3a185c47fb6c8aefc21dfce2e2bdb2e55735a6f710b6209bb76f124a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13401b06cac0ef5520ffd181f3d5cabd466a9e3f48495e1f42005797944e3666b3c459a40a2461a7c901a2c8fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7c8ea479b0d3c430f342355d327c96c5e23cbb53dea94e223e8d295d9580c4bc6c7f20738a579b3f68b0d60b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac3a8816d3723eaa4d4144a0126b5437a760ed5c6f7157122db6057358eb8cc500daff0711853bd3f50a41ff31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ff9ef105b13f3c387f466d0ceb5c81ad435b99700aef75e100ae022bb0a4cde7c436fc8056f1fe5590e05225f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163170c4ac54fca715ab6016b38eab19b8c3f2b9fa0f12d8e43a7d8683b35d906281efa623e61de9204366fb87c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15faf7a3809d4e022a91c27d3b45d8332d2a6d8d8f60f29d5e3d5ccb426cfb70ae5daf155821631f36edce61a60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha68af05de2d60946c040113b2aa9ff3dc05dd0ff2e52192c6a62b28930051dc6ad2c9ab42c1df34a979ac1144a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e8d7f35d12d9afefa29f31683459b2babc6616c80f40c3b4acdf015f540ecd4b94f0b907c03fd476706b2bbfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h723c1df407e7ac652f62cc38190afc50921cdb3e9c73f89317b883fc9798699b1e68284394ee795e594bc997a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1907930c8047980c1bf167f2c5205bb76692b12e3157db8e4113febaeac73bceb328e8c2caf69173bdaffa6cf68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4871eb4e624a140791ceb6f32d3c053c82fabbb53368583f2cd327c9fc8095c0baca85ffa3caf43d7db7716ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4168867c814c6fff197bae9c601708185d5cd9eae399a1740e83b6952922b047b56f8e1e7b8ba207997c305d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc292627b0f86a08bf2f2107664c4fb0216a3630e3b809ac5dbb94f13505518a57555a8024d1a186fd1a723ddd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h393e9dde19d2827ed3a9d255218192f873d89f83d4f8de7ba2a85ce8bd255a265e65686f364adb13519549333d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f85017062d52a1984066879780c33c0bc2f54f4dea804b770612acb9d64b3301b5c58295181eb15003e6a6c5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc005b56f9e92505b1a8787c18ed01aa36ba07f08877df473fcb2d8bc5875336d5d423969ce5aa99dc2c061245;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164e1917c73ddd60a7efdb896a2cab303a61b3ff3a48e48d5d625248e53d2b80ab4e35a05f6233a9cb09124050b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3260974579a6538bd8835070622538c1edb09bd56c58e70b4b121d07003f35a159f7a8d2b123e092eb9732bf60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5769170ecb42d36e3fc5cfd1877ecdc8896acbbc8ac32dd2d425110e29e136b77508d9a7c2e2749ce827373a0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7424d0169f9a61f5133b3ca27bf223fcab505c28d99d2a02ac063c3e404787539d6e8c119255395995e643da8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133a6f198730deb4df50b451b66eaa5b2576992964520368098da672323af3ecc7858029f40f3a40cb8bde424d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aea4c417f60c1c6ace53f5d2a926f7e9980412141c6de814b73599ef16b5234eea59c99128a137be36878de318;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f8bb528cb503f312be6fef0920f6f8eb800ea89f325f5af3cb0ef91ca84f6f0e0b206909672f0dc49dd5cff72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a3b061db757052dfb57c85f6dd2801a62f2d9a8ec7d981603da67783aa7d1f9e1fa1b93b65cd295d538f6efbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3aaff395f1c33baecf4d0abc216154ee90b5d7f4dcbd704cd2c69129104aa80c4532b201005a3f2d23c05d2579;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143aea45092a4c3808e6dbe861585c46ab89ac9d6fbf62abc1b70d2a4fa8f83bb372c48c30b91eed1743bed0f75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc26aa6fccfb630503b896166ab2b3ea4ebc9d7526f371eb5efd32383dba00eac342bdffdc3d65cb72e7f2718c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143cf1cd83e70f0d2980e150dbf6720b9ff823ab7f5d3bcfbfe113cd6d12c0a3cf4e268ba7e4bd67f832634f352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb4ec81b05b669447962c2f2e63187110da5bd035f7ef07a763ac8293968dc71fb923ca99ce4309f1ad0479df1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h895d993e22b621e5f9a154e592b3be0251b2042626aa49958e57e9186db30c6cf09c217f4143a3474bc1feb0d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107f53ddd985da234bd42eebbcc65ceaac2b2c2b757cf5feff814e4941e48fb9b8c9536dc432c245ceba42c70d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117e5a4b39ab87cc885141bc655662a2d34beda2f1d4c83ebd0a68abee736f5af8911157e709dd226d481ab6241;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8e05a6953db60acdcbebd973377677bee35a3ef8473f7243b0395f1cab10d1d91c999d196d3d89df48f9f8dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc96dcbe1c5cc72b05860f4a7d86e7835ade3c59e820d29776acbd682a9273481d63630d59c0cb4966cc337e680;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e40b05ff0880ff4bb800fcc5cf547472652af37b1a758ba54b5980be8d233a159843d13f3e017ad7fc8bad150;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12275c7839386e452f640900cf6f49695973b97dd5f35d87703fad9bd385f974999cc86c7e4353c993603284932;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93e87f47a59e8b1f2ad2b64654f9e7f983fb6b01f487be2e6e1edf22b52b1f6a4e082754a7b01ac844821b234a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c0e43704268b97369f383be942646975f5b01ebe3b0d7d6e47bfa199a4030612656fd46c4aca766c9a56bc9d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a31d7d95f34a9bdeb292530650d17379130e8f640ab41370eb81a40ea5082ccd220dcd6011e0c09f25b3f4d57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dccadc60ee49e620b2b36e62a6aa8b52493530e21b9c73d8ae7864d40e61ab25dfb7a49d183885d28674e395b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbaf6c022071ae0524e86ecaf6dff7e68c5256f227e28cd1bfde76e82847e0385b2a0f3df07fc1194d7f7032d99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d108974a51f131d62741cb9a44e357dd0767a6b3c659a7519b3156a1d959ea9107cba6e6ef7d01e4ec312b6f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h972182e9db028cb0a6faf3589c175d1cde5dcf061929bfa0b92365a09584be62a2de1a9bb0c334c7650f252b30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7318b745005ed4e5e0f0f7183be6d5cc4f158e62a1007c72eab3ddea5b5c31b697a9bfd20f19e536840c8e85c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb74dda885b49a2e1225188e4ba3d49776186ab3b4af351eb604da0f319dd12dc9c0b58e716a56e3c1141d8e3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f50b8eec75a9eb098eea7edc2a06665d38c9b514172365da82c52e7b2d6d40d67a44dce3ca74f838814a7c6ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he45ac8c6fffc5fc6e11a6fdd0c6dcca7bcd1b82130a4e61e9123394ea6722408ab3d3e653e691ee8208fb26c5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f65fa4a220537f603a1b104d95addaf8ac003d776b8b654704d5f021585769ee4e24a4e50704195b37f7f2262;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb574c1bcb6353a5838e0dc55ed27341788629dcd2308cae6ab518031df57b3e35c2786f0d44d650e26d3353ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170afc59ca87596e7f985fdf50c38315e5f21cecf72b19203565cb7e84a72489acafa91988f1c8ed74bd6c09b09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fccd64865f1a9dce15bd0b6a98dc8f9f6cbff4f82a48678450f4d461897cf63f6079603106d89ac0550d6065d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0cb2081208f7d196987058a08c338b61da27d835f79c132db4fe38b9dd6f28693e9c2af3dcc9f43e213873236;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha0fc57d84b59ef089eb32d8f26f9e809dd62c21f0c4590b693ab735da90b21d6c863e8d795eb3d04096d80a424;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98474c68a262eca546dc51d68110712c3a5a5891d956f1d780dcac59832a3d604e46b0ef549cf28680c9c630c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104e88ab966466c983486c494451e2e25525bb234f8767f15fee579765ce00d3a75e34115d28169129abf90c982;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f9c8c9b9369c45c94f90aeccb73f9fb02796d76f82c7d3a607f53e22516c8909e05c629780ece52af94c0b9bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16eb1b096f608d14db09cebee82544623ac47b5e407b6f07773ace627e5ae4d1525b9ae34c58b798f15c76da5f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h329ae39130dc004d30b281135f3491056dda5ecd6a71244d197967d843a35c584b6f08ed8f79a36d3e60771685;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1daa8cad7f3df24542a26fb2bc63a1f4e828ce3d0bfdfe32ce50bf4bd0cb1fb9d7dd74d2e1281305e00ee0206ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9f3c4894485c02f5d2cb87ef3fb5f9e1d7dd84d73425af66455b1f976000260de89b2185416a199cb99eabcbe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19fcd4567e2171a63557409e0fe4133ea08c0aeb9611cac09b997ce094b8ab79066a1565627ac0d1dcaf9ab86e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccfdfe8079ac8f3a4777fcfcdb32e48f826bc21ebd606f71b296cdcd390f96acaf69fcfae9f2559b063ca3815e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a445a245e6348dcc7c9579bb0af77a2f8839da96ebcf01384fce60c29edba684cd62750e3bd8dc8c6836b06b0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1dd8913389fc547bd59281368352e02ca92c79968de3ad7abe81efe8856247156b3da93e74d7c0a3c663d6ef0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1761e4027b100bb227031f94b8e5ca5725fa8b6702eb518df03becaddf2646eb7d75abae7038aef8782d63b65bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2aa6196778679ef3a0dd93c9a7be6a66028533cece0729452c8d54662c47a5da89348e9e14adeaf983c2bab40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1042f1b1ded1825dc3e2f488c8c6e669932c22469d1ae66392054914c763437913238372e042aaa8805ae808f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd30596522780cfb8b55bb4cb022d72da2c58ac39fa92f8e026059356ed995b4c1e338cdd60d5c8636ef09de75a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1530d9f7b5618c1a71f47831b6fe62fadc872d77d34aaddd43c03e1c0f4f2bc0b08479410c47d3c063f3e8e0ec8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdef2dba21e628a146170111f1a13c13ac76bee3347a051eea979a1779383cfdfa5608aae8a264c0c5a1eed83da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc0d90fb1a277bfca3ad9d3b4c96439f335b4cceaa61ab6a9780a198f653e6666a24e927e77196dce16aeaf02c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c53b455742a1b9d0d47a2f27482715ff9cdd6501b1e0562178b025f72766ebda77b28fc8bfbe65d07b77b4444c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de20e70b164f9b8fdf95ccd6a821fb38b1f40457b90d26523f68fa2b33b76b77d0d46516779b8cf1c73d3e5034;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h497acc8e2da8a6552efc1e34e4a1b0c7012faa80a4bfeb5ef1f1a7634f9818596a7a34a4586f33a74b4ea54020;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h867108bc9e4c654d6b9863619aa3b5b7084e70126b0474942fff01a716f9623eeed17c69a57ee61067ac9b8ff3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf9657e088e7291e9c2104162f9e33c48068bed65c5972d4607ad34abc32ccebd19541b8faa190fc7cee7d829e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d8014f9032725a9a01d8bb78bda01b8f06e009b348fef0b9442a188a7d718f3b08f7470c496139c43baf8050f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86302d71b7cdbf206cf135aaa78243c985812dd1721f1c32ff2be228e6566de7bf5aedf8685feff454de21fa93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d374a8291a763fd842218dec5b7d969d5e1d298112ef2c807ab2583fff38e73ad1eda08c47cc766bec61408b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ae48382e733ca339a65aea8b4ce4ecd6671bf9bd36f16446fdd72b19982015ad9722261c094d9406d6c11e2ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c54c80b3450ecb990119d88af884e6ff1a02cfefba20e854d4d11bd7b0ca9df41af3725f24aa54d030cd1e36d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fedb92e721d6895167c50667dad8f632a07cb800ac70947280d3032ef7aab020f316beeca955bd33787b0a594;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196732d0abeb45680db8afa8b0ecf2c23e0c6a0bef7eeee20135640d00170c693f9f83ba670854344c31bd8bd2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d660656dd586150806228377b480ffa6458c61a6be3717dbe643943cc7110c4447a0a3106d402bd1f18706698;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18951b0d419feb61cb5ade634f92153780265771896cc552b10245d1f14250f9fa22a6e33effde1bf654414682b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c1f178fe4c09290efecf988dc5beffb8784106c23930df34bcee4277125fa7756b6de8c53c45046dab1e5139b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92876b64e1d6c4f3c90236f7dfa485a8bdd41168755d95c6e21a924f34ef3a2b141deee81142d7614953e31b7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e26efa69a0a8d652278e864459b4a7a7477a26e2b57e242d98e345d8ce8dc84d677ed1e9217ba69987792c876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19726f6791c88ad5c0dfe4110693168a712686335ad029079558dca4b4849a69dda1990280e14741dea8771fbf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a2f9b115399114a577ab407390ed629b44e2798c7fe929e409c80cf08820c15e25673104a54d15a82b9f3f80e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d2043906319e7671d9ac3b060c26ba9f7b848be1ffbd511873ef8aa59fb4852bcdea640850e95c50a479d8ab7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b8f0638124c0e9733657db12e3db7662bd7a0423a0441c1a268e3c3af25499e1dd16fca681a85d74b0608c955;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1177f19f9f42882c2dbecead6d29b615542d0c3edf998cae06343921a02e19611be90bcfbf54c7029b184c5f904;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ab5d6c797d0d44493a62063ef1cf908e7b6ddf764d594dd1d5159760f995bfa5650f878284f9afd98d3ba5e99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1696d65959b30cf86d074bf988577cea7bac7583217275270b3f1327ae0db05644e4c28d1c8db248cbb38c7b121;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6375f46626c1c96fe411bf4f4b4edc679af8e93b437972e90f83312cbc8e000ea445ca180a5137e2f787814d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfa066eb46eca3827c40950bb7d3f8c90023c19957479886ccd0256a40012cfdccab38190b96f034c92a8771fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15340d3992a5a77aca1d4a2560b33bc7b0237cf871de4c7d88128a7e6f668dd338b46e2c5bb67941e1c47c9e1d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h868fb875d28e380e61a81f403a33aa68fd82280ddeb448b4eeafac989a7b25c2b6cd5aaee4b0c9f5ac61913ab4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1081d8bd0b325605aeb86440f19847a7be0d1675cd182db20f0649a5e159615ab1bb402923a8d3d6d9620b2b187;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cab0ea353e61538f7380406da73643ffec0f07f7d3fc9e6c13d3a7b7df197fade14a25471a480a921865ac1959;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b1fe1bbd72f05c65e84b61104d89516ec9a4b083b91532b0f74e763f2e524376c6a68e2831006147d6aef4d17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106c10a3f5a56b86bac079da074bce0834fd89283d2a6427f1a5b20d4072c709631cccf7c49e43bce63e444b5ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h551615cb4144229af5c212a63c949840b6bd92520893623c7feef725a9350d34ff211e9263433e5276deb507ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25a796c568e2d8627338b0cd339ef9ae984fb75fcf471f43669e5d1cbf378e9651a11fd99c7fbff4cda1816138;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5cc5c3b1d7bb1ad130329b00ed85612936a5cffa4320c0cc71f245c029b10e7c43911422de7eac4a1a34627d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1c296ec3ef7f13c538ee5975a6a94619aac7973d3fa57cf6b6cd9e68c3700cec3df8ec7910f7df6e483eebd31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d33851ca1b7dc58a76e7e341b282f2e95f4c4051566aba4914cd97eee4c6d1273a38a3d374b3a6ca0d8b17c918;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1533f050516ee64438c725160ae254ce85f5ad76faead52eae39faffa0d982fc9aaa527b2d7076e0fc9a852aa93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130d8ce343669d6318221e3633c309e3735663791fb5ba684ad61d10dbbce1557f9a7a2cc40601df23e1cd09bce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76b158a1ac9156ce52c893de521c3fdfbc8bacd464d6725a4540c04b721f7bed9d987e147e8547f11fbdf082f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb90fe29f7ff989ed524bfc3b4683ccab2d694d408d5135c2e24fd9c0c696cbceb161853ccaf316d71997448f4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecb19f3c970c5a1b49486accc662f1a7890d37cdd7b91efa335ca841d01e6a10b8067cdd5a3033667ec530bce5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e015f74326c0c2e83e859d1b0396ef7faa0e77f574648af8b5f55269d64889eb1a9fdfdc1f5b6fe12772a2523e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc10f927efad97398e7e85eb78f094b51effbc8ec8d5c7703eefcd944d2ac6bcb05c02fd3f2b3adaf85c7b50b13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1009ef85c6a3301a43feda4c227bf3010ae8c0c4287af378c960335793f6456463bb95d0a338a711b248ccdb591;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d41096a12f816dc4018e38d0d457050474921eabbf5f17bda5e115668c72667d36c777c7c9c7e75462f2a38b94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61c919c703f859a9dd0d6b07220d8f8998241ea4c310cf1e90b479d16fd532deed75481ad4a6814e9c50b35e8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc8d32da48328e196a2310565f445603a0ee45efd30fd61c9bdd8659ff988e1ed073ee691ab17c488ee3cb179f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143ef3abfbe04053a8b793bf978d52fd873f545390288081349f012ba3c144b825dc000278bc38f22560196bf7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b77ec84cc7a4337e5afe1086ba288608afd1f8ef651258cd8e6ce175c7cf3c8f5d569cc662a66e3b588185d54a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c79044e2bc3ea2b69f6c74f4d68e09f553a2ddc3d6e4580a8e5c990ab04a7b1fd42b3cce7b36475bac720d1dc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h21690a93a4d6e65d090488c4b48d49a402217959d01b5b758265a79c327f90fe1c8cb85d5ef37c4de7670f37c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1092a1eda783407b4c3a2ca5d4879f5ffa4263b8ed29c846d6c6443afef0f606ba9313360103cc7efb4b574ceb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h129060bcb7877b43341a5f95d3420ba1f61dd4f179647c9108335753615de4dde438ceeab88e107b3ec44d3f5c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h312a6cb63c34457239294fcfbf30f8c36542ed984f67f7ed0d9a6707aaccd6284f163e7140f036c39b6d321ac9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7aaec30127920467c009d387ae733dfccd1429bf0fb2c9b556bdf50acbea19a668b79587d5f3c17ef71c2d9eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cc8d75c0c1decbef1d023303b7e1cbfe0d13a74a8c578dd9724ff941d7f77ad2ed933dd9b7d147e246fa42d92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h783f64ae564610358137f139b8a436564fa8e2593bfabd9829d0f80286cc065b2e13a849d262eea46ec8090825;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ec4f2e85e19a8597766615d2943bd61ec057ef5380ffd6e833469e84da8524af242b2b8ad48c48f73f67154a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3805c92ad8549cf0ecbd8072cb3aa9ae66aa28f8b01f6f90344b32f6ff9e77d0824fbdf0f420b53d31d508b6c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1661209cb59fad400dbbd946620e78aa0cf6c2cd97af9c7eb2db9fbe0e640cf402b3bada814c5d5c6a8cbc62e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50c120eea390c05a6f3a2fe45d59a5a533ae1f484e33e91cb174f46fa3c2fb87b62987dbc2703a3c4eda34f9e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187d307badcd3962bc61e7f85e7fe0a6e1d3cd936d4057aa2e2db9a4e770166f5a5a7043aa68101a50dcc571592;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdd861132bfc8f3672b37265c1b03244eb369c20aa2227dc3a7ae3696f03287212714c9cfe3f182d962be08d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e710ada350c066ad1f624124c020fd6df855f5f89540a7582be26a418447b22658e5c9683061deb7c22ce8b6c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59bac7c875f05c8974e81f2bbc05fe5c1a9952939f2b05e2043cf7a58b02c9859e52041d0f4aed4139bc5f9b08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d658e3c3d75801633ed5ba079c195465e76eb75cbd17489831c827b60705c87d2ecf320e14b2ddc0bdcedd2e47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2a7ea58fc332d73ab7ddecb1c58647f500e53f0fe120b699c89d9469220a952d068c7ab8c4c4f093b14f36591;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82cc371b143a0307cdc04744a6568523a23cfca7c330d2bd51f1ae8281824a8f8b087cf64a2ce62fc3b896547;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf95d298468ab1aefe3285f1e63131405a73ac9eebc77a2b1d31c1c6bdd2b8e7b30d7536c12320109fe20338b83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20dc5028d1d1687b7ea10f7a92fe900ce332b5a55b3f8f3d1da315704e135987e34ecc0fdbac6032363e61d3e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4ee547621c0e3bb0accda9a9b2b4c89446ecbad8beafddfb1c73fd3b403c335c5149a2f52f0add88679d0ab36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1673a3be260a166c6c6581dcd6274ea6fb22e34803bda2fabcb0b2dac6e126f45c47da8d835d88127eddedf5b89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h252747fff440a16085f4bf98ed95093811d22ab6079e9e1091aca17893432473ec9d23458fab0456de458da914;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b44d5a155851c307ce20ce0be6254173463e47cc762b69b7b30a82d3387866a6f19296b74e10344911d09894fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ccfa3bb1fc2bd3215ab28220a7c30f2425f9c0c3efde11b472b2c486437ab46be58bfc6151f6067c6a40589d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1176167f972af905505c48bfcff74f40ea2588b48f5cf38c84ba5df8987aafe9f8f1caaac0691260502577767b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a06c2e265949d03dd958d62739de70a8827ff27a41eacfee3bd886deaea85c59c21f35b5ee741acef8e61add30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18842c1d7b8d5979ad9e5669e3a2f2abfebbdf513e77a5fdf4e43e32a36ea5acfe114d57fcadc62f156c2a9adec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b61208cd92362fc0b756dd40846e11172782940a25f61cc6eb730101c4e802a577e5b7e4846bf0a6285bf3b02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd35c214eb81d18620a8c998a3d2f25be66673d14818aae002d4961d76e9670ed1dda814c617c7a3c4da5ca6440;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4f6a7ffad50d6cb513585f84f070692f736b526c78a6215725996f4221bc3b806aa0e30ea5359ef4bcbbc48ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb35dd0374934125d4983433a970067625540f3d76dde4736c2a2adaf7dff2d334899efee1ddede9f373ac5030;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e43105a54a6220578cfe22132bd6ff7b78621a776a3e8e944d5f479e95dfbd09e4010cd08bec9b915f56d54bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b00b5ce9380f8ceab9cd5c0197afb60432cae66a349af05b7d7e55bf4e5b00044528644facf51906ca639a439a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1947fe12ee6d6c0daa45d819af9a1433c6f9ff0a7f2799d4760e1b6beca4009a15ccd8c585b31f83685e03d21cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4ac9120192dd650d17e48eef294ea530de3401ba07c07533353498c8f004cccebbfe118588b7400369c6b5657;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a5080ef00430dfee7526de857ae33c1202eaf56c68d1d33701c41467f7a38e0cd0e2f402fbd37544e3bbc2b095;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dac70ec80769c5e8fefec4b41d83b05652be50e271f655919176849d9e2832c28f1d212c80a7ade07b71e68676;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he480668fb3d42b7d6c2a1b1d10a2ad66fdc8b4248decdacb78a63e6a2f23be394393b9a24fa3dc614daa619032;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fd7a5105ef6a05b99ef91a43d04cf8f2168067f45ce047b084f2f47518d786c701e2a0aabbda12e33d0e30eee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161bfe166ffac94d560c043107e3b0544fa49e0816fdb9bb7dd990e4aebb651dab352398a03b957a8792b5aef62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19348b551c90caf576e13c42c1df594e03d38332f6ca6951b158938a3f35663978e23c93fe0caf6b51840333dfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bc8b55113f714538bc5c5dcec058aa6b9b0a12eb3eaf365aa012711e509536b6103f92ff54e774923e2fc4636;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec8c4bc6f8a921aa5b8ca96915ad42bf3feca51e8adc978f08ce41fb37b48957dac0a3586cbd7b0bc80f89fbf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h904ca50ad38ac3d5206358d42527379f2be6c19cecbf889cd25323037dbaba6c4d7b70474dd365bc7edafa61b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdae4ea7842fab64f4191c310b392d05288a4fabe32c4cea1c5ed530a33bddff063e00c530d6405e36708568bb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h457046271bb547e99be6ba1085a86d4f89373762be84052a2a432d1710304b9f14a1be31f806c7f537581ded4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17400ddb61a59cdc322ddb10ce6d202afaeb65b1772e69b3c48e2e06ad730968ccfd037e0889234d3a6822aefa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb65c9377f4d18c6635e211464a9739ad08cda5c0d78195a0d36efed502d0b3ec5a54d9bcb582c5f9ad5bc0ecca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ce432f4b303d6e50e1f73ad9feb6911e5965a5715824dde10222791176963a88f38ac25c8731a137b4617e83a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd571892a3c5023b7b7356f46510059fba3a3f3b614eaa2fce3746f706f6f3bd32be57bda6d013ddca29cc414cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbcb1bb34bc891ae7d768215b24730efe2e415634ec8d0361e85676e4a97245702e0d7e559c31220fb58e3c2585;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h96a00c5a3ad6eeee0ae4c29f0c278147eb911c6059211646c75685ceda5c4b7ad7442f50ccbfa0d12598221481;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ceddad3550ea6ab625c09a56268ae74a7dc6f3a7114ff492cefceab1498bdb8d4322e4d8969ee50dba9b9eb533;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4c855d96b1ac88b87e8774734bb38b446edad34a7a3459af806c5ed51d3ecd2a1988d633592db12ff740c0d4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d62ab0546001f927206e8d84c7597aa037793acdab987aaad19761981e0498d2dfe83a88c21376d2b02c5a31a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1864916cfbb7bc4ce9ff70fbbed4d502bc1a03ecc174af4bfb2dfe2f7dc1b334eb3acf7d50845b301a87c4ab352;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb102b6947228e888702ecc2863ef0d0b9ef79281bdd84b8a0e297c6101f05092b3eaa1c33e483967b13f44ddf7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd743792bad894513c0f8102010f31cfe0ab829ff6a735c19df64a348348abf45d4f1e9700850d9c70a6b48e936;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4bb88f3c574ed03e09c70ee28a7dc006244f0f3ce7d0d55eca268c9455a59a25529dcaa2172631171b20a9bf19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1303aafebe6b36cdd2867f17efc025734261d8feb8fa02ba27b399b0b7c3905c058955431a1bc78eb053a84880;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f59883c032ff2e11936b51089a711ba3d48576c0ab9c0202c9fbed90c75e6bf2dea6c1a1b152426b6e7a8cf15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ed17526d5e4cd65dda53e7d9f10b75bac0d47651c1488ad0dc371048a4c67eab09ab4d0d7ef3188b609a4cab5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1579b58eddd9c6010faf29584316e60a6b47ac641c6abcb38f3c3f7211c57ca494f4ecaff52f12b096f59a49bb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185727adb249b42a855402c7c36f0bdba629dc51edaed5ea1b33ebabb4b7b21024fd047b9d9de70336336c96627;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41af7effc2cfb0bedea408c3266b2eb4788b64c4338375fdfff25645f4a3035f42223170b44435a3a23513e12f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd9ec6cbc69ab5732881c608e3bb47c067c9a072671f89d528edcf332c597e1c43192c32e921d89138ac64cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133eae895a336953b6dac0c54b9085ee43c8e770eb506b0187c01bd6576d332684ec9f444c460de5e05e8bc36c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h717eb74ce776f74cd9aaf0acee614f8d03f0f5634eb67f9daad6642f0ef486b44cc5992fe0ecb6a4eace235217;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1d112dbd2b5f5b862f34e6a22a576cc28fa87d02d8bf9b9e4ec3f89bf07a9320fa0833e24ffd0cc65820fedd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaed1e65d5236eb5f1475124311b1bc93de28ccbef32c6065b484b580aaa4bc2edb9f208ba674078a666291b22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h703bf6cba2da6141fc6d91236429326b3d4a4b5722e30a8da49c90c42dc244195fe3b5c7f372cba0700d8efb5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b98020d765c9db709f15d909f5b849702ecf6f2f7de4f2e40f04bf9621debbd6c6d884235e889f802c5a8287ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e59326220d5ac19f31264bd054bc57e7c17efb096d6dff4b8a522cb1c9416bc12158e5f04e8ebb4b4838dca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f76eca4a1c1e2b3e66d0e241c9a4f075a905c1aa2b3087d942f422586d9e7e3a35b1ca291702e415096bc581d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7f36972cd5a007cff47e1cf4445147e08ef9c7a8aeec44d04dcf5ed26f9f0d9bdac720424a74ecf4f4d411b3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfcf47c53414abd5feae68b9bffeb801f5e5ea500b1f1514e815ca1db2752fc31648c0ced96a6c9fbaecc158d62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e0d05ff9a60cc82aeca9f67a4027674fa08a817b4fad78d1a4ac79be5103c7c183185784a4543f194b794fa43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h327f8025b0030f97c1c607ef01cd935695ca3187d222e8f1695977a11e372311c829c3a30ff5906ab7966fb682;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ed4290a8e1af2bcfe3a73ecb33414cc5861fd68192d5c16f5348d37074b5ba4b4cbbe5fd7d85713b3ad03f432;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc9fe668e3f1b856d4075cbd2f446dfa9d24df15e3a989029ffb6daa3b4c5964643abb422c74e07b4e4d5715fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e752d80c29f8665dc7284dbe4e50c3cee99598446bb0feecd8dc5df248e69d30890f224e7d941724096fbb0da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5976fd2fb8fe6088fde43fc98f6b6a57767232b26e7524232d85445c8cd9ed0cc804d63b696fa72a13d40d66f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'habb93bb0e39c25fd9bf649989a7cd4c7955131c89f872c267380c434a3fa185dfb8f24ad0073ea0d414a8797bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed0c4e126062f83df84d9d8ccc8b8b6dbc970703010e3c554b539d586ca674fb47adbcf585e054bf9a0bf7867a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36be1b151a8ca7d489675562b83970645b0872c4b164fbe99486b8a1f2f79c8a09967608aab9b49cc69863d9d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193fd9eef46143c4790b3febf5ffa2cd62a9b728f657a2758bf82bcd1724a5b34c23a8ce0f4bbdadd85b2bdf103;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d0261be40565e02b7836ddbebc7c9fda9211ff80ad942cc88240fe2fe2ee50e02a4e2a45bd7cdaccc4f670835;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f5b4d17071b710daf86ba172fbf35c25ad609cd80a3a58340f4cad60f0ae5370372d9d447591eafd12e72ddb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b61ce277865e9fdef75500d8f3cd22cae385844d48f7492894b59341fe88f3d868d72271effc29418908fdbfa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd19e2b19efaaba86ac960caa49ddf0e79e06ac38ee7d7cbf5af6b4baf3bef6e3d90f226cad0983ea308a3a2b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5e6450a2548a5dec610cbc9a7a2bc59ff3100f9e990c2629ccdcbf57b3c5cac38dc2e94484710b52f2b1639e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140eda16d3f1b982e11c917b049a0f706b744aafa3701de3bffbd1ae4a249f88bbc1f53ef85990b08e6b618ccf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc21e0cdd264b2088938035b5b652b811fba79ed919b9aca9c5d3c14419a1956de27e5e493c01491f55fd6ba3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51a8a5e1682b5ceea2df2ebdaa04c938a93441c0a686f242b6b05a84cbc536b1eb6915e0af58535c7e3a5f9bf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd62e2d2506c5576ff0e9e77610d58d11206a8eae5c0ad4bffde02b39a574c41d8e581acb777ad84fd5343fa9f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132c60ff452bcb048a4b050d27d43ca371a8940b1117d92c58705a6f38beb9126fdafe87571f8931e2e01e5daa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe079aa492312f2902b4c765af978be3609b3ae962163e18a3b34cf66251f46aa5581c74267143ac1f5b9ac99f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'habbed3830e3177a5ea61e038a30038b277994b73b8f29e0232ce2eca60edf8140e9423909d96d8c79395ed87ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a22fe6097dd0e3e25318b361224f34a3cda30e674a4dd299ec48ad6e92527c75a55408880c8e5949512d369657;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd95383f5d0696ad4fb395641aaf63d749f53d63046ff6ce71418b274ae477fc6c4f3023955f7b622aa05b087a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f993492c1a9ae820d6a92c87738156377d3d6cff447911593a463056debadb3c6de59f6c4929b6bbabe63f7519;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c889cefe9f134abc8cf60801917c83cf4addd8e6460931491a2820aaf63c023cd5d45b96e95979bcd398feb571;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12acd00f2b45da768d9dca1bbdca8210e38384b581c5fc3fe8feb328836f557f6157699055a3304645cce8fa945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h426f74364d44108cfe259fee442f26d4735582bb4acff6b9855e30222cfbd543fa82e0b3d2100e29b04d5a40a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26e19cb054d9d2a02aa311aadf53448d5b65253020d8ab2baff4bcafaa282645e561df62dafdb29625544a885e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bfe7c7c6b4c9520eb6b6792e0e9f67f341164973bb8e8e1b145edc9d4e2ed4c1364052ed24d007d1ea9c801b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10fff3cd05ea57d9d755747ffb4df37a52828d5cd751f3a4f8af0d50d2b8d3608246efad49cbfedb184821e4554;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97dabf6ca1fe0bab27806184465d7cef761e9af48d70baedc320b61b92939112558236eef42b3f3da49b7d2fc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ff4310e7cfb85a01ba334e4d7240aac7583dda5f4e4fbee62fae8370b9b0a4da96761961ef3767579c9706b9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ff317523bd560c5d328450ea9c764892623e9baf2a21e145a3a4e5931b2f227f25ad2ef16d1a8ff25570bab51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1a9db3cf4f47678fb8726b24735b3dab0816a949e7f597aae5949d57804bb147b9d2b70865ed4d640f8fc3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134665d322f55d22e6a9c1534a4967b89c9dc1c42dc290841be2f00d625f1b30a44a382c338edd06a98313bec47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33e86b9f2194877cc879b215fc0e8cb6dce8abc2f67526c54abf5e6a84ca1b74ea34a32dca5b7cd240fafac443;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haaaa9f4dba0082d574cb2cc5e89514b4b20a3789a2732efadafba98cd1332a971037e28f7a9de0d1ba3f0ed4dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c8319c0b2202638744c9ec3e04f2f806f782046080c129532351ec017fec5f81a1f2ebf19e8acee94f928c696;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7dd084d109f8f1a81b1a47ccc5adb80a68db9dbc16307a698d59d3cab889927993bf02b835cfcc6a8af93e593;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19226fc276ce9a80c8fb64b667e25cb3236a84c96d9ad939edc6ae2f5f4403289ae280326a64d05bc082ceace3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b93ab207869cefa1c0fe3c583450c9cfd0fe710e8aaed9b012e8de55a4f6e1a29a02a4f43fde87f415303d53f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b168efea730990eefab5f1b3f50691e2c61e0051c54e91f3e26e7cea3a7b51945f9a53853935847aacc788d1d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cac4c79bb11bfa0129e486c5eca8d1ba87f9bf71d21b60af4a6648c93576c3c0888bdaa56c18f90f8bff7c464;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191bac83b72da54e63b71b9f8a4a3a65c1a3d5886c20bae927372a25ca64002b2d20f10ed24ddf0c70af054b8ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1735881cb7d76799a6c9e3eee015a8c7cbe6000b165dccf71593ed455381c8260ec637d4d0256c012ca9cd7b48c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f80eba69ad9a96793dcc3182c1e68c1dbc3d4feeefa19040d5ef0c9c8fc531b4250f16e8d8dd12f921fb027dfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b8f095dcfc875f4d7baa07cda10f82ea46f44b800932117b741ead384adbbee2a49c2988274dc7fc20df4ac89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3405dbf9405431028f5f5d34f7e1825b9a31abf9818f051efcaf5a4a5198d95e9a298eefe28415baf9fbfa3974;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc4ad7215b74b0be3ff590ef76da5bbef5b559a3b5d153ad9990b0ccaac33a79ae67581a2aa6a58a9c319ec30c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2a749e6d6790b87e0a8980dd96a8fc7704a06b8e301bc3924f66226584360289b5415e0a757c0dc25f4553e9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e97a0ce716aa5de1867dc01f4683d849653809d8ca27d0cb86cbbe73fe0cf84e084b2dc9c56f5ffb0a436d152;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b472a841b16a6d9b14497ad42a9db52c1bc8a3fe61ada150ba4f5f912848ae4c569cf2bbd2c64b2267f43bc951;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d6f0e5d6fa6808ffafdfa997caa9103c44ed77accac2b90604371931e68a9fe7d7dde229d225f131f3c234938;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5ab32afe9c1f826f77bd1f5b6a266af2bf48b0e7259c526dd6408192f54c4ecd2da50d1eb4cd49f890d9a531d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf41d9fb9b268125ef25ee52bc4f0ea5775e395f2104b74cc81c562a3523e560bd0f5f2ca52f177edd886f98361;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbed18d48df48dda7d3973d39f9ca1bcd525e104a47c8fb0f3fef4e69c4122a05b09a18c62da015643ab27900da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80df2bd228e2d4e8cdb8c00d638dc2707eadc1a5b10fc628246cf1e043ecf833a8794df1f42b648713e87752f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e498ee537573ea86ec781be42c89bae2ae80652abfe4fe52eee407b06a5210cd779ab8927bf85adae75f48e1b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68fdedc4167185c77f1318a2513f6c8da4634ce74be34452fc678826293501d2db158496190be266d25b6cddf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bb2595823af401b98334f4f4970d214f98c5ec362f591488ce494d765e0b45faae928b5aed4ba2c7c9f7caefc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c75f9cf4ca3c42f61f5706022115331eb10633236963dc3e01d2b28bab79ec2ea2b0dd3752105f434f4c1872b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e983255bf03fbbfa4a9c51e16d28101fa8a906b46de14adf33e5118c72c451511ad374720a50c315360b2d25e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3082a012be411e9df42dd6899b3affbd6583ff5aaac383776d3d2ada4666dba759bfaedcbd55666b1de5d92885;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bed23f5e3ceccb2016c83389d0a8c8e74bfbcfe836501ba6db521252ec0420e398c43dc0b4c1225dcfbc9d295;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5f16880251dee2565669405969ce23314b7dfec0024729866b1ecdb55dbec6b8bee4ce87c3710c847a68d6b1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e3c4004e4aab54b1e2f2ac80b9a156f3ceee18b76521d902fe74f30503de3d03cab53d9dc6fbed885541e9acd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1493218d91c7fc66a40765c5165b94eea53e340c520958c2165fc65e7dc4f30d05966ef2e0943d4b2a88f1a1bb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha22e18001716c885ee1b4fa04f4ade2f93cf4dd6466800671d38c6d85c7abbb95f650bd76776b59279c7a18595;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1363d4534bd8ff6551a151f9d63210afbd7aad426d7ef868aeb37340589b1cd83be87dbdc5411420f563bea4def;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a09ea3529d3d65a0e1fe4f6bc66801ec9652d5e1828e6b18ab6ba020e29b2edd1cc0bec11337d9e89cd569ff2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2362a1d646b6d18bffd479e2c42a46a3a1e603325b90e26c61356a3a5c8b4e928766c2f0568fa755270d8f08b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133fab60db389a89a63803a507aaf0dee983f0492bf4cc8acf3c09ca0ca19ae91c4f018798c3fc97707526fb5d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc9151d321e77bca18c04be26fb479c1a7ffbc1a09d42a2b4d563857000391ec597da8e4c6d07486d970e14046;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f2753504a24f0278b7c8ccb27056a29032309338e9ce8abf687feb2645a002ad8fc5126c82023cb9af6ed93fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81e0509495b197b9b2eeba6817dc43a435b043f5b0e17c0d2bfc52733f63fed2edd6d721e636a36f3d61796ef9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75637acf0741b8a54edbeeaf6aeabccdaee098cf28b2771947f7494e95ce89c70b8caa0ed3242cde2d69d85f98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he66e3a62217938ff3bf71df4a2d57e98fb6d16f9e265658fd15193ef3f049d021de06ca3014933125295e7faeb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h468384718b4591f0fbefa81955ef6246425169805f12737eb97daa04b7df5e3a9032fa4316cf1830068cc01c8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55e0304f3f6b9dbb7eaa438a7b679016092f08f2e62e6f283310f6551d239ae8e06ca1792f34463a9da1200183;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a36986edc518e60fd7f83013875cd9606a0496c2c5637df09174f1b22d1bb2b87d59a1dee4b5edd8a809960eb6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ced77bdd0601eaea2f063693c3c6b8fa9732902e1eb44e91658cdd04a75b5aa78f3930bc263e499e17dbe84613;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9f5aa0606c2bf40e9d9aaf0f9c90f76f9573ee6fde8b20312de45e0515086edd21a46dd94f8a63ba8e281ee5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h464eea88b2204f9442c341c2cffe5d1f11c590a0179b2cb8b5c09c1aedc171978f039adc32e716accd300eadec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea407e32cf823c6d4a22c0dfb823393ecfd87f9fcea7e8fe15229c0e7747b2f711ad3a63c382036bc972671d37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbba889300a6d1653f1798346bde7da924dc000b959c24ab34640f0805e6e28f519a819efbbab49f49e566c677c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1719da5ee62d48053ffb8995f366902797cb86e0edf9dde93cf3308808ebf5c059bb4e86f271dacb915191920a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f5c698a59ee9b18190bdd47ef1e97507b3890ce8fef3717a9122a368ba85b979120995f478f7c2034a8e0959e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33b3527cc155ee78e6183f2e4676019bfc6be588044e5f16fff4e9530336b788d11a8188fe0ed1cad3a85bc2fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ea6ed41cf9c3c859ed97f256b6c7a6d661072bcca4b0bcdaf5f3615c6a7bd4d0a8d2a6d6fe3dba5e4d6a2a1ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134c565d04e7b00f39755ba272e8408c879dc94b2cb4cd3eefba364b5113c6bd236b94df854a4c11a78217db5be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150ec845aeeed1794e86e69ebbb989816fbd2eb2792331a9d37a4bd4bdf0e878617db57409ebd603a0f3de3b813;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b356184b56ee71cc7f224ae4b1326dc9d6c3c579422cf311860161f52f6f1e284074b4077f6f1d03ae84df7fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he58b45a0d960e8caf798e7d14851d0665075938c118d4775a65234cfc816beb51b15d168ab5e9b938d1f69c9f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3699ebb6857ec8b828765b334d219f630779f62ba98e2c578494ca0fb908c61c21748faccbac5083f8490a586;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aacc38ad2da10bf2bd7b087afc9906f6203d9faf683974d925a6e17da9d8c9c76becb1a21cb5f6106c7c04cf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147e47de9a5083397089c663d82ec196f2cfc7f1f07b214ca371eb8bcb68d47fe2b4142380b9113f155537f0b9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb9ae8bb054cb6c31985196d274d61693467eb1f720e5ba88eef4abfcbf12a08d0826be0294bd5adb678118ba1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169cc08d5a636e4160069e7b1a5625589f39ebd8a6d48a86cbb4cf101bb80c8c7bddb1ba516f0467fa62057639c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1111b24c6f5a5e2ee0357b46067e1a36ca9578bbb040144861fb71eccc0b35a0eebeb06b44fd55008e5a52f2180;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cae200dc30c30f71151023a302b542acab87e8b68ef627ad78c6c6b2145a21ddabf8d73e168f2fb39dcbedfe0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he11f6687768227ecb8829412dd3228e7709fe118e595a86bd9fc5a26c31c4fecc449604852d7e1ab7663c04634;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d8de7c6d15a632a64c1923803c809a9d8208b08d81df62c6cc36300f26c9b0de7f8efbdc2de0c3da6c8cba7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1720a0e1756698b059ce0553baf6ba676b867ba483caddca6647af5ac568dee9a56cee9e3519cac5d0d0db55c46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafa290142c79fc9e48ce02bc5032760bd0f98d3af8c516e138e107914ea2fdc8a043f7d2a2493e472f444380d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c43984b345559c481178d3943bb01801cf858ec147f540e97b9b20200a08ba484766704a6a98b856cac7cdc67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1331dc1dd44da7b2dc6ba8fd1c3831535163e82e274ed56e60b3d8f56185b272b58ef474ab9bc893d330ebbfcdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d63a3e41d952cf9583d2a0e2cf63a3c43acd8b6c381371578f7ce738ef1f31a3c86f9668ee3ce1b79068cebaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25990651f2278eebd7b0426a0ebdfed164842f705c0f190370a7484206cd4994358b9ac598719e195c14ecdd18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11089c020ec5e6fc896039eb45d8d983bf4eb471e4b356c9536163b34b799bfd65d8a98184c8b4f991755b23cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1baab7e9726cf09741ce5a8218464d4f57c4cdf374970236d37ffb9faa9ff0219275ea2fca435c4b224b8c3ec16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45b9727e7ea3fad15d2c0afc55582a3f5dbf38c7b8fb5d9ea47fcff61d446409d6d0d02b6bf62ccbb993d7edf0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h370302443a860bfe9e26546b36ea358fd0976a47f419376fa4dad1e79eb602bd1b451bdee8d645fa3a09ea40b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49a3d2ff62cb416570b554717d556fa94eab4f26b8a69d45a94e9999a01e1d42815f1b68da1724c12f5c77ce01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14bbc59ac509ebc7137c21992df9c00bfc4492c62a97d38cc3b1e641926f35f5eae977536c54bdf0c2e3f17e8f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb39b3c0a8e051c815fbf96c11490f983b5c387ef6ef005f4f223b767ce18c69b526cc4fea5cce8131d90c049f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0ad6579b1a4ffc3f7e16e1116f8aee5319be8bca7a0643acfa3ae865191e7d1b55af9d65008c117187dca9903;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcde8055f5796f1619e5467c36bf4726664ea241fd99a5595b6bd92c6314fb33db4e4c28869b08ce8316901c996;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15caa0729127c6d555fe4975976ab9cb948080114faca75df0c7470357222d0cf09037f0935ef9f81edce89fc0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c828e156ed21c3d18d19f4dd3abdcfdd578e7e1077d8ddefd1b2e8e724a258479cc059724d1e13c9bfbde63e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10733f1da05b2134f7a707c53449f95e603e39023a42ec43a5528d86972b4715a2ae1143f31f705399021bc32c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173d7a0af7bd245e00a9498526d20ccdec983fee33c28a0747f9ef5caf7be161d13fd7e55abf4305fb84d38b91d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23b90b40883748555f37151bf918a72fa6e7b3c18392438e9ab760af971417d2c99bb784a5f29d2b1aa06d55af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdec47d08e44330c6c7986703eb15b4fff2622f20c1c0a6c19d31f05892905749c62bfd21d0089ca6e70de47667;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3b956b1ab2eaa65be23d73ff39ec5736edac3709f7de7636e47bf2c1734941ec04e789f8c4bccf6f59f2e1b22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1558446f39d2efed246d20ade68c0978a6db5543f3b9ea67e07c0fbf6d0d9db45170f9d7b7af142546fc0bbf8ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f53f0efbbab437f7604e4d92fb15eb9e80f950c224fe1b7217baabc9d0a0950f24a937eda618f4e1c0ea60f823;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c45b07187dfe0ce70474c9fa99729f6840b2850cfa35c2200a96067abac109bfb314b82218628bd56e7b8c672;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1385859675df761c0eefd0be79138ade135f2e384a12d08cc5cc626aa196f73f74512055685ffb75d30f29b909c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf359157e4841e8bf1af79f361c650279dc8a138aa13ab3411ba81f679824fb69117f0112b4cb57616a53f2f5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116aca192d92acfc044b258f561f33250b2f88cbeed6556af1d31c9aeddb473ccc1086a4f6f4e04a5112a045d61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99b07e6d2d444ac324eb46b38d9b2d0377c918d22e9f1f363f7a9d4d1f6618d3c8ddafb20e4fac23d379aac098;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150de39202ba19d262d63b4add3ee6003978d6c2a41aeae98ba5b8da6b4dfd2284d8bb3de5f88fcacfe5bb87fac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99ee789a142b9a37c09f09a970984f1f4a40c9b1592dc91c89ca9da593b36d9fffd1b07f6e8d355423170e3ad6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa08806d710c9fe7d8f206afb1a05e9bce4423fae6ca373359cf3748f04a0c1b5a0f3d26c7906a6656ea5d23ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144ad17eb1d147ac67af9173880f9af62463248cb860c3225986c65d1deee61b28b350f3097001104ba68ceb744;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eba62755ac8e3be47dc356a9bdf3c37b39bcfef9488e12500b0484bffc0aa1e57ec3f5c957e9f0bca7f1b8e334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1869c9d56df3e937a5b910f021815cb435bc492bb3a3b09d2bd9389beb9b20bb270de5b3fbd6edcb48ec651d44b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a24fddc24df621e753aee73246e28cb47f5477a9647632fca07d1ba1fe9a88d702811b9a0f3aa1cb286144dd9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f6d8dac78dfd85c1b0cd3178048ce1c48a54f5924d4964e545820be0824a5f896e99b6a209a0964c1961d437f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef811b5d9d612c8f1b7a4214e67354f0778e9b0a6f852289dc61e63a06ee6eebda432c52a7c2c5a2b88ebc8d5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db5146fe752a6fa0c3b8ba7ef3e91ef8d783d1933a61c0912ad11b871a674c6f5954eee735dde73b4d14d04fb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ad8c4fb2798f1adc2b68c7a81fd77e84231aea61ea5cc5c78282e7c9988e375aa2ef8a09ce2a32b67638b80ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1389057089f3670a06671749e916ef318d0775f6f32482f4015d21f052068246a6a40e0e6023df127f4a4a012a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d819f653bf7168772430a59127870289350fdcf392d83cc06e0c10c3779d6b3516adbc516cce90d05c1f18cff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e57e22d1b3f61d7a6f0cd92f84018ec528b2cb475fc0498ba6c290fd3c606dc434dfeeb99cecce6550851a950;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea06f872690f3066a9f34ac35bcc4c8839d3ed62c66039b023b322a3b5e56b4d907d5f3066fdc85d4ea57e9c7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e66be8260c55c85507e2677fa6315cee1b25e577ab7317aaae164edcd3ea25a8725e8cfd27dff5012debed175;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h177182d443b28401782038970fe664c28665d095a7caa94f5b3ebf03119e1bef2b5abf47d0902131cfbce399847;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198364ce9ef45a88bdc43af4c330a666af229f19bb0b23ae3b4beca42cdbb39df49b9c5a6196c7f62d7caca22c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9ac85d9710f9e7a9cfdc06a31550fa6b4bd22d2d26bd7ccbe92b3e8dff9250230ff173f4151cd6cfabd78add7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150db9fca81966ce35fe8c448b2d30a6a671eaa35686fed7fb796573db6e5c69929104c0aa4cc3cf34da509808c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5420ab48988d37481fc00379045a39bda1f1d87603fa6649d155eb8745e166cb21da5542fc41ff96d29518310;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcedf29726a70b9ac96bd1cd16381c35629721047a433c785ebd2608662ec7889aead17b3e9d23a0e10af321011;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e57110ce478ecfa448d323bc5652687931231034b8d06391e6420a5bac594b6d8cdfba36249567e18256220d22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d45ed118af774676e8bcdad8732d6c0a1f800237d9b0d57ac936d2d3f34c701d36d899441971bb934d93431d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123a0e5b56a6714b85c1c919ba599229eb7c411feb24fae8effb291a424301072a30ef772fbbe232f95780eed5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12959dcc21661ce240c6a6df7276a4f67ffd0472df0be49cdfeaa1e4d27db15771193e4f082b48d4d8b5ec14b10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1b220929f2d2c4e1488984af218152e78bb973b0e72dcd6e18dbea3dc06eb5c9912b7ee26dad73ec14cc1e444;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd109dd47155960c5fb21be04bedf51b1d6684b241f0ff6c7f76d56166e3db667effffcc57f434c4aac6a059623;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a8d2d43a077fa5c0207bb4e5a4cd2375648fc86b035fe3cec8d311267cde30b9b345eff065dab4064f80080cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168e20d545e75cbcdf331a5466957363f409a45a46aac29ef11fe49eac181919db804156ef58c0e0c2b739bb207;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161dc326db729850c7f83c0671649bf800db79e5d73e809eda63349b0f9deb0f9741fa3c5c3cc5b78d40dae36cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71cced5d7555845456cafa5b901e9bdf29d85535716acab299c873889040b548403588f071ffc0dc71fef0ed10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bfc27735618bf6cd238cf2a7814b2c94514ec720a4c1c70b2e79e1ec098a81569f2505da136872e7e7e97782e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6922e9f1585ac7472b79b205d8c0f12968cd3fb3c61a7534650546f4801ede9fa358582184e7dfc83b5f575ed2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13778b90680743f6efd4ea5fdd54a4af98978186438d4b777b4acd10406bbfb7a5fcb677351aa7de4ae74d5decf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5771791c13a289f04f208fe176b5ec40c115d613d08af58f6c38080e1aadcd71c7cbf35be4e958983502e4d7b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb24693c75fd734dc6065eec25e9d038a69ea14c68c96a81ccd9a8654bd9234f030f9149940c8583b4e7e48198;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b4e2ff605d25ae2d364bccdfa4f2e7d6c9c36390f5b530e6eeeceb223bf6e0ad59a9985e26c4e782e031522b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15337bb5f9d1e2bf856a791c94acd40694b5c1d3bb11df604b29c883075b5491135f832f6cb94c8d3730f0f561b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a17caf02017f3dfb2ea4db360321419bb354f93e97e554956f17f693a86d4fd73b79a5b092230806ac7544768;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e6eba5e7dd60690320e1ca8c51e704565b38de47c70d9fa7b0be034d0fbf6e46455963ea7c7e9155ee1e51cee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132345062891e71fe30bef03c76e9ba0267df7dda20ed20b2a4161c2e4b391641229afb801d05197031b0053692;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h558e1967c56e7ef6b52292549fa050537ee3c07388fee3ee6e912c0db7690a390e5febd2085ebede1d769acc86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f1ea668f2bf7ad5533d68b332f3396798fe4122e116fbe436a9a3ad8149f5b8b1829370de40b77e7271be5714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he35966139e1655408b1e34943e55dd87777b17caef122c07c4da4df3e8db6cadf349d505ced48622bea668fd94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e70310f68cef61efe1a207096d608beb60a2f5298e67bca36d7bb648920b46266b7178fd3072403db7c6c2cb9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5be362af3e398470c48c801bbfad4ae3d1c01b0f34b1dea7ee0764140306f05703c27892b8b81945a80fe15086;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ed76db51b50784a5d07bef50df2463d77170d3f3d56ca742e968dc46a96ca02d699f29d2933cb9b032bc2db00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha59d1a54f2a5af79e637925c3542801c6b71e5392b6142fb32fc0a223809cc5d9e83db51707df55a5828aaa33f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c17eb387e8d9a2451ebe0681ff48f70044b2776be4a95d842babaec3a02bd4a60c5d3108d8c7787c35d97e19b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c28f1cea3b2054dd87cc59182aa105446877d7a242676bea162f075646895e7943a67b419390f6f8e1e6e5adb1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd37d78b089e657b61b0eda1f200b613e2d46c62ee58fc305896f4e8b6c478a4d797386997c7764eee970297b81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h661660bc0be3c4f60a4d17a6ed58df1756d80e120d350df782941289b4b7c983fb559434241680684b7e30ca29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f0dbb68e1c0878c82fa3fc5581584162829c87c462758e492fb0d7c3e6a6d674568daad486024c1b7b0635607;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cc0df7c66a66cd9e9f2ffa065da5868a648b447d03d5f5d07b31decb0521ed2a87282f6c2a73e09c2fc7649e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbbd918389afd680271e0dd340c4dcee18ce18584813ec8c673f679e169eb9b3396f1cd961c850527c6ac460853;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca50d31ee3bbb89bc9fb294057cf2cb9eacab94bd2070649e4d583582ecb7dfb82b3a6669a0fdb2b6e13847575;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd423f87776f2ade61de3b7e0f8b297217990412df65cc274cede26bcc7099b104e0c93e306dc9f7af34c322bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff73e93c41430aeac9803cfc6a82ddd53f3b53a64cf626d54223db19c1039eadb7c8e2064423ec9362862f2f40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h398bc0ae9f767bcb911c98b876c3a806a48a2f39a2914b49831f3d03b9a62a73577e2934ad8394d988d6c346f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h278232d1b0222b495284b032e29992ff48c25d9ea9baa4032940dd0909c61c6ceabadd4a7c7cd2bf29df04a22b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de004da6a54d363b6f096bc89d13cf77642d46d38bfeef9c61afb31dce06024effff3c1cfa76f5e11a378a9740;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdce2e0fc2991d22dc20531a0f2e9ae1817140ec640363b2ebfa3fb3b2e6cf09715ddb2f6012ca019b53cb4b35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cccab71eb3f78e434d2ceca9268f48fd54e7a0e6e375c41febd4b03d13889614c74eb305b1001d6c2ab660ea1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1193615511ba50b4feb9bce3d1192f901b698949871979ba7b2395cac1520780d2345ef6d0a2f0c24ef8920aa41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b84b036318b6254b6b8cba5ed9efc02f7e2bb818fb771d82d61e8f01bfe0f834b166553bde29418fdc3cb16dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d6a2f2bdabe09729cb91e10d88090852ca4ffff98b1078f16f0e80b4c14405cdb1a5a34591d3080aafeddbc09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b769bbab3cf18ae2d83a918f04e2ec28450abc0e812b31527f3bb60f52e490429c2e95d1d523d5fc2b4c973a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h190b4e966ca3573ba6e47af0a51b9f34298086130ee701368f22b6452cda9bbc6d11df5dc5e91b0c0052478f5dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5149d2a255b9c3c87620acaae7ef75fd84cfb69cfe5d37744c626a3e2e713d814ff162019d30698fc5b8b199eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5727d469a2a8ad13723c6c96525097ac945fb3ccd896968f4e7b216628cebc43498766d6f8c6f0d635152c1cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7dc432fef2322263fb30a80e82e472dd35371cfe235901eefa41398210bbe9bd71d7e832371426a7a9b781c322;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc688779c5494672d75c56a685603b8ffc4c886e2718991eaac7985baa423677ab2d0ed103eb975979e20435b17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cb3919027eae400af5f16be9a9d481c4b2c9b6666bc020acb87eca752a37989bbf2b6c075371777b8756bd9a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e676cc49e96b7574304f6d9629bf7ef8fb138645682bc0b2f46afa99661692d98b0eeaf5518225d122df6bc4a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1643a6747d9dd5e73fe23c10e1eaa99cf7891ef3a82634fd80ce8357a68d44dd3e52b00ed6a467654444d371e57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fdd346a42ae4aa60c959f039e54bfc8cf80aa3e769a6aa8ea833518bcd4fcf8279efb49ebfb3b4a9cd2d39816;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e9445edd0eb1a731d9d14e379f9aadb523b6ce1055b8d6ebfe26ee3116299d064b2173ffe12bbd803fba93a52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c90839e362490f26e38d9d481f55829a24ce77d6496bb19df2fc088193cf92751eee9b5c93744b3856ac7f727;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c36ab0125e421e330a78f2594728280def5d2aeb88d5b3df01405883c9a30a3d6300cf297a23e948bc5ce5cd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd3e233e45d1811b8cca8766e7f972d296a97f23d8be87b16ca4a8d23c1101b97d29e8549198147559bce7ffb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55e582af48f089c1b24c5bdf792907777d6cd74eead7cc2067b97fe245a35a49335b3d88b584e21f4b07c521d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28bafdd6684bc4bfda57a55acc73d4d6f938b114ca720b5e2147fe4fb02c49b14a5f6176ed98169c81b4bac600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42a3f33644f54b2d5fc351c2ac2b3de4012574679af118b2a1d09640231f8946ebb7f4412da06c0e3ddf63c7b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97dc6fd78d5b6bf524e38ab68c743cc5000a04edf8f36ac7f75e5c35e02ce6d4e7f770364d394f15aa769f5d88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8d994528a00d1b825b92201ecf3195abd6fc93e9d888f3c4f97a0270803475c2971ba31922174cbb678ce1df1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117088c274e1a1ca1e871d00ccae82ede3fa7e7149c66f9dd2b96a912a2b9fd4d6f8ded800ec311030c503ce3bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c6ad10ce903a1a2adf963c0572fc4102cb3cd904da6b3eb5fa5a8834f03c0d092f906609dc940f3f36e295dc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64aa85187fd286b3400f1d13ec46c8c1d1e5f653de3043375afe5252dd9946165fb36b2171b051cf85bd4bfe84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85981f0f1b2ef1fc249edb9b928aa0f2333158d70e74ac96dd74e9e5312470772e019c62fe316f088a8c03aa7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1063d5018334b89ecdee194f17fa281b3e4760dc4dc65146b7239f5d63a875fd87a13dccbc443c839d069e8d25e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1451a1d015765292edd9c02bcb3dab933d76ab84fdcd269d36f4a7d29d09b942fbb71f75c269d856cb7f5540a26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193679533f827274a99f53b679b6307c7cbf03561ec2656a7a3a138191cccb7f45b82d474892fd51d9b2f58b57e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf887537c92465979c89a13dcc5ab0be43b86dc1df7ed84baf58cf46fe3c60d1a6967d26bdae1bd458b40134cd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1375fad6a6bb0dd790a30938c810d08a6d395b016342ac2049c0b75c2c1ad2922189fd61f2c52fff868c8ff4091;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1482f4f898b83625a210c2d434f9f1b05eb091ba0861425c2b0b6966afda28be62e50fefe8e72e989836f5df1e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9b46f9debe8e8353dcb6ef526115d3f2086c0051381a93c149efaa4bc5baa642d47851974b63180ec3865c510;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd33543b0753774beec54041614e0f01ee44672418e6f1aa124f4ab5663752153619bd13401b2ed38e374b9fd29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc351402838fafa70d243cc130c03f2cc2c997d441e7b1e1d810b54297c72d7b2b5d444abf2b7399bc41271a682;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c739b897f7aaa0a953ec5515a3ce4eab06a1af4aa8402bd2f73bfdba86116973c857f7be988755b70209e6ec73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198184b904d3ffc806fc8ea1d8d5aa337aaeef001c0d8675f3bcc28afb9f10f7bf0beb8b81aed35e47b38d15a72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1557b53c966916b8d3ce5b5f457c0aca574e862ca7d94b2ce4a2dcaf68132969877380bf109aa9278be10e44b82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5ba84e982364c7b4d62c0cfcaa48d2bc3cd162b7bafe9ef31a51a90911f93eb0f6805b6f2e960eca91d70edbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h634fed4362f044355a643a6000e3f41be4b1b54294db5db338d8208af4f19f0b5d7a898e7be43e7607ce635e4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cdddee25b91a00a8afc1267830c4973a5f71d66307cbf9f71ea5a00cb3c0077d1d850ec5dbad0c87ff4bf31e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he05319af8f9c86b238d15f929bbc0e9214b2cc1be4bf02f10b93e311f776da4efe5a5f6f7f198bf6ec46a7be21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b55a31c8a7193fc2e50c032e6d0e92bf8c87ed5fae83926d14737f3157bb2b9dcf35c6ee90df343e91ad51659;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77d3418c4c20e1a2777a4bc1b3431e6906ac25f679769362d4e8448210529caa3c06075f2bd07d6b1bc23f517c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f6a53063fde9948a9bcc4461d364162ef684df8cd259bd90bfdced387909c0a05ba19f9a282d4a4357b78a667e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h638fec915ee83040940d3de8b9cb34b27e34bc09cc9ca728f32d9c0b79b2026a853f224caa41e9d65372c93cdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d67696152840374baf4fedf82c09bb1426e301326668bc04b3ffaba317d13c3209d47944cedbccc58c575f7fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40c84166b0e044eb64ff1f096df17b267640a0e9fadaf8ff7754bbc633e143cc2fabf88db574f1d73b4516003e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba80242327121c22b4b6d4d4ad2b9923c2bd12641749caed2dd99c06f0e7f091794e56c6e2e374ada005e28e3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha99355ad2fcb395a10d30e0875fd120ef9d1d5a8e03376db9559c4f37fc33368c525973d159fb071b4a08cd968;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e8989585a20660c78eed8d5c2e7cb023da4efda7e52655c76884a1381aa4c3694cf15577cd6e42b9595d06700;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15da0bda91336fa305bc8012abccdd94b8c9ae0f5e5ca8a0196468cffd3c69efb94194baf415f557a487dbed39e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13dd6c3caec87800d0cfc6e04ba5365c23874e92a8952390c1cbea8c797949be227110003ff89511471df8feddf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c5d9a010c05f3c2c099f39e104eae30eb4e85a54c33694cf765db9da57d860d8a2864cd031fafec68870991ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2605c85483ab25da2f4997a072fdf6d91af84bc6476c60d59d534b417ab61881e6ddb1aab0359a9f52ca513e69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5cd824c3161e8a925d2a45830b49824bc75b43011c2a253947e60c55737e9b67d72f12d3f808215fdce35d294b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e5a5a0d1b1b6f166ea72152e6ad4c81b802ee5ed5284f1b914585053e99c359305228fccab41895e7e3d0e8b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b1078f92412a7b83fda628e832a64e8a30af1d6948527d88a1eb7681eba84f98c2460807b7616d09274d35bdb;
        #1
        $finish();
    end
endmodule
