module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    compressor2_1_32_12 compressor2_1_32_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_32_12(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [0:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    rowadder2_1_17 rowadder2_1inst(
        .src0({comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [17:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [13:0] stage1_4;
   wire [14:0] stage1_5;
   wire [16:0] stage1_6;
   wire [10:0] stage1_7;
   wire [21:0] stage1_8;
   wire [28:0] stage1_9;
   wire [24:0] stage1_10;
   wire [29:0] stage1_11;
   wire [2:0] stage1_12;
   wire [0:0] stage1_13;
   wire [7:0] stage2_0;
   wire [10:0] stage2_1;
   wire [1:0] stage2_2;
   wire [5:0] stage2_3;
   wire [6:0] stage2_4;
   wire [3:0] stage2_5;
   wire [5:0] stage2_6;
   wire [12:0] stage2_7;
   wire [5:0] stage2_8;
   wire [12:0] stage2_9;
   wire [11:0] stage2_10;
   wire [11:0] stage2_11;
   wire [8:0] stage2_12;
   wire [5:0] stage2_13;
   wire [7:0] stage3_0;
   wire [5:0] stage3_1;
   wire [2:0] stage3_2;
   wire [0:0] stage3_3;
   wire [2:0] stage3_4;
   wire [5:0] stage3_5;
   wire [0:0] stage3_6;
   wire [8:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [1:0] stage3_14;
   wire [0:0] stage3_15;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [0:0] stage4_15;
   wire [0:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc615_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[0]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc606_5 gpc9 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[0],stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[1]},
      {stage0_7[2]},
      {stage1_8[1],stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage1_8[2],stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12], stage0_6[13]},
      {stage1_8[3],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[0],stage1_8[4],stage1_7[4],stage1_6[6],stage1_5[11]}
   );
   gpc606_5 gpc15 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[1],stage1_8[5],stage1_7[5],stage1_6[7],stage1_5[12]}
   );
   gpc606_5 gpc16 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[2],stage1_8[6],stage1_7[6],stage1_6[8],stage1_5[13]}
   );
   gpc615_5 gpc17 (
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_6[14]},
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage1_9[3],stage1_8[7],stage1_7[7],stage1_6[9],stage1_5[14]}
   );
   gpc606_5 gpc18 (
      {stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[8],stage1_7[8],stage1_6[10]}
   );
   gpc606_5 gpc19 (
      {stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[5],stage1_8[9],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc20 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[6],stage1_8[10],stage1_7[10]}
   );
   gpc615_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_9[6]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[7],stage1_8[11]}
   );
   gpc615_5 gpc22 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_9[7]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[8],stage1_8[12]}
   );
   gpc615_5 gpc23 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage0_10[12]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[9]}
   );
   gpc1_1 gpc24 (
      {stage0_0[17]},
      {stage1_0[3]}
   );
   gpc1_1 gpc25 (
      {stage0_0[18]},
      {stage1_0[4]}
   );
   gpc1_1 gpc26 (
      {stage0_0[19]},
      {stage1_0[5]}
   );
   gpc1_1 gpc27 (
      {stage0_0[20]},
      {stage1_0[6]}
   );
   gpc1_1 gpc28 (
      {stage0_0[21]},
      {stage1_0[7]}
   );
   gpc1_1 gpc29 (
      {stage0_0[22]},
      {stage1_0[8]}
   );
   gpc1_1 gpc30 (
      {stage0_0[23]},
      {stage1_0[9]}
   );
   gpc1_1 gpc31 (
      {stage0_0[24]},
      {stage1_0[10]}
   );
   gpc1_1 gpc32 (
      {stage0_0[25]},
      {stage1_0[11]}
   );
   gpc1_1 gpc33 (
      {stage0_0[26]},
      {stage1_0[12]}
   );
   gpc1_1 gpc34 (
      {stage0_0[27]},
      {stage1_0[13]}
   );
   gpc1_1 gpc35 (
      {stage0_0[28]},
      {stage1_0[14]}
   );
   gpc1_1 gpc36 (
      {stage0_0[29]},
      {stage1_0[15]}
   );
   gpc1_1 gpc37 (
      {stage0_0[30]},
      {stage1_0[16]}
   );
   gpc1_1 gpc38 (
      {stage0_0[31]},
      {stage1_0[17]}
   );
   gpc1_1 gpc39 (
      {stage0_1[31]},
      {stage1_1[8]}
   );
   gpc1_1 gpc40 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc41 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc42 (
      {stage0_3[30]},
      {stage1_3[10]}
   );
   gpc1_1 gpc43 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc44 (
      {stage0_6[27]},
      {stage1_6[12]}
   );
   gpc1_1 gpc45 (
      {stage0_6[28]},
      {stage1_6[13]}
   );
   gpc1_1 gpc46 (
      {stage0_6[29]},
      {stage1_6[14]}
   );
   gpc1_1 gpc47 (
      {stage0_6[30]},
      {stage1_6[15]}
   );
   gpc1_1 gpc48 (
      {stage0_6[31]},
      {stage1_6[16]}
   );
   gpc1_1 gpc49 (
      {stage0_8[23]},
      {stage1_8[13]}
   );
   gpc1_1 gpc50 (
      {stage0_8[24]},
      {stage1_8[14]}
   );
   gpc1_1 gpc51 (
      {stage0_8[25]},
      {stage1_8[15]}
   );
   gpc1_1 gpc52 (
      {stage0_8[26]},
      {stage1_8[16]}
   );
   gpc1_1 gpc53 (
      {stage0_8[27]},
      {stage1_8[17]}
   );
   gpc1_1 gpc54 (
      {stage0_8[28]},
      {stage1_8[18]}
   );
   gpc1_1 gpc55 (
      {stage0_8[29]},
      {stage1_8[19]}
   );
   gpc1_1 gpc56 (
      {stage0_8[30]},
      {stage1_8[20]}
   );
   gpc1_1 gpc57 (
      {stage0_8[31]},
      {stage1_8[21]}
   );
   gpc1_1 gpc58 (
      {stage0_9[13]},
      {stage1_9[10]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[11]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[12]}
   );
   gpc1_1 gpc61 (
      {stage0_9[16]},
      {stage1_9[13]}
   );
   gpc1_1 gpc62 (
      {stage0_9[17]},
      {stage1_9[14]}
   );
   gpc1_1 gpc63 (
      {stage0_9[18]},
      {stage1_9[15]}
   );
   gpc1_1 gpc64 (
      {stage0_9[19]},
      {stage1_9[16]}
   );
   gpc1_1 gpc65 (
      {stage0_9[20]},
      {stage1_9[17]}
   );
   gpc1_1 gpc66 (
      {stage0_9[21]},
      {stage1_9[18]}
   );
   gpc1_1 gpc67 (
      {stage0_9[22]},
      {stage1_9[19]}
   );
   gpc1_1 gpc68 (
      {stage0_9[23]},
      {stage1_9[20]}
   );
   gpc1_1 gpc69 (
      {stage0_9[24]},
      {stage1_9[21]}
   );
   gpc1_1 gpc70 (
      {stage0_9[25]},
      {stage1_9[22]}
   );
   gpc1_1 gpc71 (
      {stage0_9[26]},
      {stage1_9[23]}
   );
   gpc1_1 gpc72 (
      {stage0_9[27]},
      {stage1_9[24]}
   );
   gpc1_1 gpc73 (
      {stage0_9[28]},
      {stage1_9[25]}
   );
   gpc1_1 gpc74 (
      {stage0_9[29]},
      {stage1_9[26]}
   );
   gpc1_1 gpc75 (
      {stage0_9[30]},
      {stage1_9[27]}
   );
   gpc1_1 gpc76 (
      {stage0_9[31]},
      {stage1_9[28]}
   );
   gpc1_1 gpc77 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc78 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc79 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc80 (
      {stage0_10[16]},
      {stage1_10[9]}
   );
   gpc1_1 gpc81 (
      {stage0_10[17]},
      {stage1_10[10]}
   );
   gpc1_1 gpc82 (
      {stage0_10[18]},
      {stage1_10[11]}
   );
   gpc1_1 gpc83 (
      {stage0_10[19]},
      {stage1_10[12]}
   );
   gpc1_1 gpc84 (
      {stage0_10[20]},
      {stage1_10[13]}
   );
   gpc1_1 gpc85 (
      {stage0_10[21]},
      {stage1_10[14]}
   );
   gpc1_1 gpc86 (
      {stage0_10[22]},
      {stage1_10[15]}
   );
   gpc1_1 gpc87 (
      {stage0_10[23]},
      {stage1_10[16]}
   );
   gpc1_1 gpc88 (
      {stage0_10[24]},
      {stage1_10[17]}
   );
   gpc1_1 gpc89 (
      {stage0_10[25]},
      {stage1_10[18]}
   );
   gpc1_1 gpc90 (
      {stage0_10[26]},
      {stage1_10[19]}
   );
   gpc1_1 gpc91 (
      {stage0_10[27]},
      {stage1_10[20]}
   );
   gpc1_1 gpc92 (
      {stage0_10[28]},
      {stage1_10[21]}
   );
   gpc1_1 gpc93 (
      {stage0_10[29]},
      {stage1_10[22]}
   );
   gpc1_1 gpc94 (
      {stage0_10[30]},
      {stage1_10[23]}
   );
   gpc1_1 gpc95 (
      {stage0_10[31]},
      {stage1_10[24]}
   );
   gpc1_1 gpc96 (
      {stage0_11[6]},
      {stage1_11[4]}
   );
   gpc1_1 gpc97 (
      {stage0_11[7]},
      {stage1_11[5]}
   );
   gpc1_1 gpc98 (
      {stage0_11[8]},
      {stage1_11[6]}
   );
   gpc1_1 gpc99 (
      {stage0_11[9]},
      {stage1_11[7]}
   );
   gpc1_1 gpc100 (
      {stage0_11[10]},
      {stage1_11[8]}
   );
   gpc1_1 gpc101 (
      {stage0_11[11]},
      {stage1_11[9]}
   );
   gpc1_1 gpc102 (
      {stage0_11[12]},
      {stage1_11[10]}
   );
   gpc1_1 gpc103 (
      {stage0_11[13]},
      {stage1_11[11]}
   );
   gpc1_1 gpc104 (
      {stage0_11[14]},
      {stage1_11[12]}
   );
   gpc1_1 gpc105 (
      {stage0_11[15]},
      {stage1_11[13]}
   );
   gpc1_1 gpc106 (
      {stage0_11[16]},
      {stage1_11[14]}
   );
   gpc1_1 gpc107 (
      {stage0_11[17]},
      {stage1_11[15]}
   );
   gpc1_1 gpc108 (
      {stage0_11[18]},
      {stage1_11[16]}
   );
   gpc1_1 gpc109 (
      {stage0_11[19]},
      {stage1_11[17]}
   );
   gpc1_1 gpc110 (
      {stage0_11[20]},
      {stage1_11[18]}
   );
   gpc1_1 gpc111 (
      {stage0_11[21]},
      {stage1_11[19]}
   );
   gpc1_1 gpc112 (
      {stage0_11[22]},
      {stage1_11[20]}
   );
   gpc1_1 gpc113 (
      {stage0_11[23]},
      {stage1_11[21]}
   );
   gpc1_1 gpc114 (
      {stage0_11[24]},
      {stage1_11[22]}
   );
   gpc1_1 gpc115 (
      {stage0_11[25]},
      {stage1_11[23]}
   );
   gpc1_1 gpc116 (
      {stage0_11[26]},
      {stage1_11[24]}
   );
   gpc1_1 gpc117 (
      {stage0_11[27]},
      {stage1_11[25]}
   );
   gpc1_1 gpc118 (
      {stage0_11[28]},
      {stage1_11[26]}
   );
   gpc1_1 gpc119 (
      {stage0_11[29]},
      {stage1_11[27]}
   );
   gpc1_1 gpc120 (
      {stage0_11[30]},
      {stage1_11[28]}
   );
   gpc1_1 gpc121 (
      {stage0_11[31]},
      {stage1_11[29]}
   );
   gpc606_5 gpc122 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc123 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc124 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc125 (
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc2135_5 gpc126 (
      {stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_5[12], stage1_5[13], stage1_5[14]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc127 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc615_5 gpc128 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc129 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[3]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[5],stage2_6[5]}
   );
   gpc615_5 gpc130 (
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[4]}
   );
   gpc615_5 gpc131 (
      {stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_9[1]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[5]}
   );
   gpc1163_5 gpc132 (
      {stage1_9[2], stage1_9[3], stage1_9[4]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_11[0]},
      {stage1_12[0]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[4],stage2_9[4]}
   );
   gpc615_5 gpc133 (
      {stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[18]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[5],stage2_9[5]}
   );
   gpc615_5 gpc134 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14]},
      {stage1_10[19]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc135 (
      {stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage1_10[20]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[7],stage2_9[7]}
   );
   gpc615_5 gpc136 (
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_10[21]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[8],stage2_9[8]}
   );
   gpc1_1 gpc137 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc138 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc139 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc140 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc141 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc142 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc143 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc144 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc145 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc146 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc147 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc148 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc149 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc150 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc151 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc152 (
      {stage1_3[10]},
      {stage2_3[4]}
   );
   gpc1_1 gpc153 (
      {stage1_3[11]},
      {stage2_3[5]}
   );
   gpc1_1 gpc154 (
      {stage1_4[13]},
      {stage2_4[6]}
   );
   gpc1_1 gpc155 (
      {stage1_7[4]},
      {stage2_7[6]}
   );
   gpc1_1 gpc156 (
      {stage1_7[5]},
      {stage2_7[7]}
   );
   gpc1_1 gpc157 (
      {stage1_7[6]},
      {stage2_7[8]}
   );
   gpc1_1 gpc158 (
      {stage1_7[7]},
      {stage2_7[9]}
   );
   gpc1_1 gpc159 (
      {stage1_7[8]},
      {stage2_7[10]}
   );
   gpc1_1 gpc160 (
      {stage1_7[9]},
      {stage2_7[11]}
   );
   gpc1_1 gpc161 (
      {stage1_7[10]},
      {stage2_7[12]}
   );
   gpc1_1 gpc162 (
      {stage1_9[25]},
      {stage2_9[9]}
   );
   gpc1_1 gpc163 (
      {stage1_9[26]},
      {stage2_9[10]}
   );
   gpc1_1 gpc164 (
      {stage1_9[27]},
      {stage2_9[11]}
   );
   gpc1_1 gpc165 (
      {stage1_9[28]},
      {stage2_9[12]}
   );
   gpc1_1 gpc166 (
      {stage1_10[22]},
      {stage2_10[9]}
   );
   gpc1_1 gpc167 (
      {stage1_10[23]},
      {stage2_10[10]}
   );
   gpc1_1 gpc168 (
      {stage1_10[24]},
      {stage2_10[11]}
   );
   gpc1_1 gpc169 (
      {stage1_11[25]},
      {stage2_11[7]}
   );
   gpc1_1 gpc170 (
      {stage1_11[26]},
      {stage2_11[8]}
   );
   gpc1_1 gpc171 (
      {stage1_11[27]},
      {stage2_11[9]}
   );
   gpc1_1 gpc172 (
      {stage1_11[28]},
      {stage2_11[10]}
   );
   gpc1_1 gpc173 (
      {stage1_11[29]},
      {stage2_11[11]}
   );
   gpc1_1 gpc174 (
      {stage1_12[1]},
      {stage2_12[7]}
   );
   gpc1_1 gpc175 (
      {stage1_12[2]},
      {stage2_12[8]}
   );
   gpc1_1 gpc176 (
      {stage1_13[0]},
      {stage2_13[5]}
   );
   gpc606_5 gpc177 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc178 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1]}
   );
   gpc606_5 gpc179 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[1]}
   );
   gpc615_5 gpc180 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc181 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[2],stage3_9[2]}
   );
   gpc606_5 gpc182 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[3]}
   );
   gpc615_5 gpc183 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3],stage3_11[4]}
   );
   gpc1_1 gpc184 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc185 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc186 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc187 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc188 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc189 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc190 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc191 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc192 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc193 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc194 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc195 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc196 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc197 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
   gpc1_1 gpc198 (
      {stage2_2[1]},
      {stage3_2[2]}
   );
   gpc1_1 gpc199 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc200 (
      {stage2_5[0]},
      {stage3_5[2]}
   );
   gpc1_1 gpc201 (
      {stage2_5[1]},
      {stage3_5[3]}
   );
   gpc1_1 gpc202 (
      {stage2_5[2]},
      {stage3_5[4]}
   );
   gpc1_1 gpc203 (
      {stage2_5[3]},
      {stage3_5[5]}
   );
   gpc1_1 gpc204 (
      {stage2_7[6]},
      {stage3_7[2]}
   );
   gpc1_1 gpc205 (
      {stage2_7[7]},
      {stage3_7[3]}
   );
   gpc1_1 gpc206 (
      {stage2_7[8]},
      {stage3_7[4]}
   );
   gpc1_1 gpc207 (
      {stage2_7[9]},
      {stage3_7[5]}
   );
   gpc1_1 gpc208 (
      {stage2_7[10]},
      {stage3_7[6]}
   );
   gpc1_1 gpc209 (
      {stage2_7[11]},
      {stage3_7[7]}
   );
   gpc1_1 gpc210 (
      {stage2_7[12]},
      {stage3_7[8]}
   );
   gpc1_1 gpc211 (
      {stage2_8[5]},
      {stage3_8[3]}
   );
   gpc1_1 gpc212 (
      {stage2_11[11]},
      {stage3_11[5]}
   );
   gpc1_1 gpc213 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc214 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc207_4 gpc215 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5], stage3_0[6]},
      {stage3_2[0], stage3_2[1]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc2116_5 gpc216 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc217 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1]}
   );
   gpc1343_5 gpc218 (
      {stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc219 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc220 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], 1'b0},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc221 (
      {stage3_0[7]},
      {stage4_0[1]}
   );
   gpc1_1 gpc222 (
      {stage3_4[2]},
      {stage4_4[1]}
   );
   gpc1_1 gpc223 (
      {stage3_6[0]},
      {stage4_6[1]}
   );
endmodule
module rowadder2_1_17(input [16:0] src0, input [16:0] src1, output [17:0] dst0);
    wire [16:0] gene;
    wire [16:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[16:16]}),
        .S({3'h0, prop[16:16]})
    );
    assign dst0 = {carryout[16], out[16:0]};
endmodule


module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor2_1_32_12 compressor2_1_32_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3d9dd81be2499927b8f890f6f2ab3be07131903c1d77dd490f50c3937df1c2a14c03f8b92342f51e681202af4874e6b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1d89176106b5ada53bc02675abe6529aa5c434be63e1448a2091d698b9b6c12f08bb5ec3cc316877c5dcfd61e255df97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h469f450d3b32e9968a8261dfe167ddc90f144ed66b5ac2195976f6514e821f1fbbb8a951f5337f80b4171cd7d93bd6c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc1ab3d26a4f7c6e860a5e65f8b469c990575d1359cc3b7f9cd11c6c09914257bb0abe01b1455c6a02be58596c857af67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1442a0596baa004121847549d4530dd9b5f7c64728a9d7f1d1e09953babe30a27523cfe5546d0f21619a79a304297f56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc1a868843958de22c527f6a97bb71df1c3764dca530f465073539aad2f4978232736cf2b7187ef81b489a93e7595577f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7e86c0ea415523bf4e193808959a56af4ee851e2fca5b9a3abeb2f28cd112019a9e2b25103bba29dc2cb7806a8d19e40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h10e96a796594c91aaceee0630d34062a5f08d53ad3c7f58dd69fd56db3d0a5d5937dd31c03336ebe26cb08f2219a8d8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha418adad191ec89b9e5d360827889831722d5ad7d9457299fb971f9541fc6e240c78c308d59a10c18122254b9f8ff72f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd00bd8b0637b90d19b972d168beecb7c73d5ad97e66071131ec4eb1aaa059978774110acdc2b6c312cb7bed4c0435de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1a4e218742e0c9fd681e1d25240ff68371674d4cbc288531088b346bef645dafa1201a6c5bfeb0a65f5c0d4f5d304248;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4c8431c53cf0cd25c81667f43c1c79bc1271fe626e3e1f4a13731bf10c825f4b1f616437b5fee605514e4cfb1b0d97c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h822035befe21f1cf0043e750fcf39ad8720fb9faea890ad183c9aa0c925bd9570ec93464fa021f75ecd65db828d238be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h766c68cf7a3ffccc0930c52c5f82177162a5886b81ae1079a0f49fe98271a57c5ab89fc8624c4f1a76a49c828cb6b552;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5437eb615616e4aa756d8afffb0a4fd74bc13b4ecda6651b82d67b3873ec07fb1d7499cf7a7b22558f0a16a6bb6297a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1f016c5667af6b4b43f30563ebe0ab509056ef6b5b1868a35ab7be62c4f04b99dddf393179fbcd8741ee74642209f9e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4838bad2d58c2d36e62b45a29b7a904fd25b290c5a29a13560e5b0b39fd6ab8eabff678cf46709e6b78b68f0d114fc65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1f47a33b0e59202e6cbb32a53a6a4f1fa7e1d15095c4d7f69fc7292519045f82db343049e0aa7ffed58cf469cfd19a89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h44dbb042cb8331fcd1db871d0860c2bd5576494d08badaffdf07d7313176049b09ffddca960a68c34db7dddbe89ac310;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h63a217ea0aa48c6cdfd396169ca810ba05d74488a2ad4238c9cd2c54a88e2637893cffbde0a8837585246358d4041ca8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h70a3de7306a5d6f9bc02013deeb9bb4358347768a0bdb6c2f3e5c83cf7622f782ecd85bd49a8a4420f01fcbafcb34474;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2e81e4ad642666fdc251601418c319775f783cdc719a10d03197ab63e82d6dabcc8b1b8604e6f2abfcaedd03c93ae8da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h165ba8b858c5e195b3eb15e0b93f5ffb2e2a71908232c34aeb28e86510e4cc327f5d40d731a363284b16bacdbb9a1b7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h394dc1f9091f29387e44479e0ae34dea149d1203721890c0540fba3a6cda6418a82cecc4acf36aecf3e617561544c363;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hae8397d435ec0cb45221d549604895efb950c50742ce6840b6e57ca906bf4ebf50e1872e2d41af1075671642be7707d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1456919ce894a3e76479088c86179204d73e4c417a9c71842879e276a2fc64cb7c826b060e88582ad08e32d6906ca919;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8b43afda84011892fb1f151e6fc23a924861a2a4e906a74d62cedcc7827197b9ffa320fbbb2e55438f8af564acdbae7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd99d3f7e42a5bd9c2763df8d340881adb30af9fb7356109e0b039948cfe18f8e4add3e156493270b57f2f27d0a3b9fee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h471b42eb8c2daa72215784836e335d3731aefb4525dadc789ebcebef8ab41118c7f78968cca4f60ede793266052d5317;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h95508e8da8ad3c62df6a7688ef419fd8801218ffa222e0a03a20a858d5e6abc8464ef0c235b509090c364b846fb8b0e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he391f6dfcb8f0ad60a5712b936f53a842b068a9c3468b09dace8dd514b725793611af0407aff17253471f3356ab4554c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h390c5502003fdf3c489b69c97e9ba0a0c0a0c11eae23f5883ba02a40c22e248223f9900c0eca04ef16acdc57728f7f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h54e9dcbb9853d1f5fbc60994490656c6ee62d1f622133f6d42238b95bba754f88ce2b1c8a5febf2754c206d5303c8f42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h62e6fbab31959afac46af12cd66b22c9205dbd0d379606fc362249219b0d3c401ec717813a6e0ca69fbd04f8fa1463d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha54f860e72f46c09d697307bee8b2b827cea459fb338801aa3fdd006119760447ed51c8cc9d522376a4fc32ca8f4f4ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h113fdc1965a86ed6c2d789a26f839d29cbd8a861b4a7ecc15e077d4daea4c82271547133850da9e03316b506c97af5dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbb9d049002925627a2cdf9cd56b32acf42e943f03f5e93aa97107d6169d117da3c27e77515def97fe7cfc1f9ac1bffde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hcc816fb1afd518831655c9dffc3b0e4f6afd84f50d39d460e8313991cb7eb96a00f71d18d0fabe9679f150d9791eeba7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc14478ffa27d912ca0737d1d5ff926fe99d46bb1190dc673357d8fce3301dbca6550c1cbfe378d3bc27a5147891a68c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd08dda348c2e556b2743d6db34cf3c148076b2a8709c26e12b49b472b73e29c35ff6790b0d06f163d4381db155ed0b9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h23887af334f96c39216f7ec24d20aebbdf63243b4046f7bf0712b4d45a43a0c4dada346518eff7e2bf407df739813e8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h17cc896eb8a835180c1491f3a1e57c46a6b2853974ba1cefa19b8aebd16dd8431136cb4ea55d3151e2d5b0970745ebca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7e07867d99625ac42437f6b9a23e7821b8bb977e3a2625cf2f9adc70978aea28c17bd1668d23c91679573c9cea54e17d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb6fc377e254c2cc1af0f9c2571261ab06cfeab7545a7ed2f89503c8bb556cd4ad77aeb5ba10d96dbec74f88c19a3c2cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4979f2dca1c388f61a0afa63ca5b5fd746f6e3c1104b922e7c15d5f9be24be22da24161dfc8a9cfbfa6ed510d0f93b63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h443ff5de7d420ba84eef32ff84ba47cf0172d779bf62877fd346b9e0ff4f9329cd74bd9af3e4b7a1275778cc1f89aea7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h876eec2a2292967ebb38188d26b37849dae48f1230c0129f7f4a056d0cc4f5d316dc8413cc5a14158c0e4f86d36e351b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5fc12bd2a54daae5ac714d5e3070bff3617117d5ed8035f12f53677c11983b27ac773e4fe79d3c8632fcfd73e6b756cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h34ffb83a775d167cc90cd4b7615f871428149d3180b48fbc6da88faafac9e8fac245c97c718b2cd86ad95fbe44bce9fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha21a2ad0739a62d434a0e25a80ca1a14999c55320ed6214f158f82c34a9b99b3479240cfc326925ac8fba7e64eed8656;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h229cc18040a48f65dd52d0bb8853d015e28cffb493860177c9e19873bd2c1d8356b7361b6d0131bb9706e3607e0f8b63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h36facfecdf7d978fd63b363af6947005074e76033880c18d3478b39fc31495de3ce7543dd246df16e97ab7df0a8c2373;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5a9ff2c83fb41948c9f4540f9f7f6635368bbaec39407d64709b35bcf76e990b4b446ec32b6557a1095c754ba0057c9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he968132bf3a8fbaa96b8bb1bcf03a47ed55cbbc86775cceb87fabe0b2c80c5e922ea5ead0cfeacad9b38922c7c1f4687;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hab3f0bcb9f827d96737c8d11d7bfc269db002a97f158932c3d6036f663e841ce69346cb87ee60895d33807330073b24b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h64b3b80506b741b777041f819a05d80dbbab2f0b1a63891a656908b68a1ef686b7ee64c40eb08d005bc2b6518199a0d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h395cfb9bf192839732b1a2296733c08b18d67ef80a3bb55121bed63f9fc606e8b0534ca666083cb4e45888a586e1f174;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5c401782f712354c776b6d1de0375c361491783e25b59be31a583aef38f1e25725d8b72396443c33bc3c0f781e0dae74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2e671f419ce5ffe6c807389f0d9268cb2615222389596d0ced92ede6b4a34ef84d1b5e8e94a722c9b23c5cad912d2874;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hce2b21559a93f4181eb849f03967c7f8d8bf3bbe634a1d10cf290c4aa67c0084ed78eb0b52241eba496eadb226746f95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5e5d3dbc47841c88bee8b46e8b93643c06d96daee5159cc308920700e4bca3106fa34ef103035bd6ae5e66dc9830c11a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6277f763423a2937ee122bbb896d9d7d1a73136e755f85c654ccc3424e1222c1f17acd2d958bdd23cde6e56d711eb1f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hafa1f50958a9f57099001c7092e554871d605296b673250719d793c40c951a42f46781777dc8e3d3e03a32901917ce31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he587b9fbfa1136b507d957883efa00c0912556c06d3bcb38946a6fe58538eb1384ee972a115165610f9f24ef0b0ed21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hed21478e8e9f1fb2d67183e04538cf3f8dcaaa7f6f2d2f65612a40f22be10dea5ab147a62bcada6cf017689c2cb956c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8a2dee52041233908a3b7001c217ef0444f1660707e143cc27bb2ec42348cb3bcba36ca438822c2c58f713fbc31fd838;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf9c9a35387f7d9331fc0625f27fb26a5806a537273cbd3b99a7949c83005326e9dd2a934954f89e9e2101856434f2896;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbb6b0ef43de7066d6c6a41e8a20605bef81d1ed55496c302d4e177c3575337ec4bd7cf089004b586c7fefbc91ca453d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h94c74aede407d6e779bb93c370be5add66e6b79c76967bbd290c8e3e44e04833343d01a57ef923cc2d9aebab1c07119;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he2254c213001718cfcb759ff72ef63b4e5ba60469f3e7219d957c35a166fcb8dc97c384a85743ed66f9398a9dee87885;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4487d4eafb951d82e28a12d67c09ba22a633b5d4c39fe77023c39540bff25e34926ae9ad8d39bcc8c94b23f8b1834e63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8a4dfb76a3e8a9bccb58a4718d01f6a1f6218c71bf74a459cfce2be814be14f4ad1012a3763e55917f89f574725cee39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7722172df6212e314035a7d77e7b3170efb97be46deddf31dd965d4e386058b49b997c3c5225711ccba4f39ef180783f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hee840a7e026dce217a4d8b305b6dcba9d27ee819b9a31595f3227b122b3456877aaede93ba48b1fcdd49b5d701d9e26b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h38b43ff2dfd284b0077c5d7933f4349bb845122e273f64b2e56f15c267411162b7856fe3fc196a99587c974403515c14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h55e76fb5f9b1f5f7290493f8537c6265a7f5e0ae08bd842f419373b47a64d0cdfeb1fb9ef78cdd36f1c4ea5df9b400e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf9e98d3ebc815b4c7870e8654beaa2223d5d8006b5ca36017fada8c697b3aa77a732736f0878697af7cdf4a86539dd9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb27b3e4f4041a81a7e41d54efd68f6f19a2eaebbb10ad53889b29caf19bd365d4bc5702caca93228ea02012e1cced12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h456b6583a48c7550294e2ce079f944ff36e96481a70301f018f54253f8c47a7483ae70031399ec9452431c676728269f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd3a1664aa3efc03b0cbca05a21d9cd2c59097e6b98f99e320c3064209f7a6f63dd8bb18460a99ebaaee9c01061a40d24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h934c2e5b93a638c7aaa3769dab7eaf6dd256d744db8bed52a95cea5baf2db29554255758af3d33e8b4faa1486d96991a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'heaa56258a1e3270ec120f0cfdb4f6f38bdc66863f1a05a12d659b462f422f317169a6e1886d4e97cb629d9219143ff62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3c59ee8eae77efed81b87fbc7a0ca0d7561405aa3ef38d6028f7d67edbd75cb8962c53613e30d64d2e5c98cbf89a272f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd975334c62045da24075fac9a98a0855c25ec36b49aa549c886f4da550f6f4feac0e1f5dce59a0e4b3834d8d00ab5a62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc4e9cff90e934c21122efbc937c2486474e6cd3ad8292cbad0c74212b3271d970e98a8e251c6964d59b55d95a187621e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he02ddae8ba6d088fb34190641a071838503814472f736e474554b0e1041d340b8577a8d41812b1c74e67fd282473c75a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h345a3c75befa280610e21453fe6315a18910b88a9404826c60498e11c3c2dd03ecedbd7534099731744b39d4d665566;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb58b81a0e48056782a3b7bd655781bb1dd84782a06d0264beea8175246788326b9706f58d62796de3a441c09b8f2e569;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h363e9c9f75b5a5d0c2de9680c61203bf617714d08e8340ed7c5e8edf6bfa81051d47aa163f38aebe0656fd173ebd4369;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6d0cefe50e5b60b6278db008d37d742a6f4d69edaa1cc28f0e3fb09db644cc6ac176a68ee22f48a3e23db44484bb5e84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd138e1de8cc26c5fa17ab81132bdd7206540c8d33326dfc1678c5912a5ffdcc61616bb1aa34be444e8a2ff0fcd84bc45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9d5e1014c4308feb2c946b1a00a72a46e471d91c9306db265b4f68a6aa6a8930af09efb71b013cad3dc99ecc9063d058;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf0c622ba81639dde3c357c1dc8da54a1ef95f96acc715cd3318693fd3b27e66acaf78864bde8246f5498bf008bbd309e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4955275d6a15b698c07ac5cadf1560078b5738e7d7461e3977284741b1c2a51c26c58594dbc4da9d85479606f7144571;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5f05a7731d2bc563834846204148a1cad2d3b2bbeecdb374136c27a063565227c002daa23d81ee18132361953311313e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbacd874922b8040e32455c26607feeeed1d61a222c98afcfd80eb1be4c858c0bbe7290d950349aaccd723b21d257b0dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbe0908ac1af078c352f89bc642fb60f9cb21c5ecc22566404125eb9a206ad53eb17f4d057265e1a997e73845f2969428;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1a5f3d6705e3da60b4aebbf75e0b12d0d86a809dbe1edf5d478a6876547f9878b14c1396d39d2b72639c8c5787daebac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb235f341c5d5e4d0cb5bac145507e4b6d0672d8fc6224b005906b659808e35969960caf01f81249b99cba1e1e1b660cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9817c8b1c4f35d6a13c663f039404e8d150f2819b104c3f5154e3553fd6be40988d10588ba7e81d526bfa9035ad9b9a8;
        #1
        $finish();
    end
endmodule
