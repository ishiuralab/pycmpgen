module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    compressor_CLA16_64 compressor_CLA16_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
        src16 <= 16'h0;
        src17 <= 16'h0;
        src18 <= 16'h0;
        src19 <= 16'h0;
        src20 <= 16'h0;
        src21 <= 16'h0;
        src22 <= 16'h0;
        src23 <= 16'h0;
        src24 <= 16'h0;
        src25 <= 16'h0;
        src26 <= 16'h0;
        src27 <= 16'h0;
        src28 <= 16'h0;
        src29 <= 16'h0;
        src30 <= 16'h0;
        src31 <= 16'h0;
        src32 <= 16'h0;
        src33 <= 16'h0;
        src34 <= 16'h0;
        src35 <= 16'h0;
        src36 <= 16'h0;
        src37 <= 16'h0;
        src38 <= 16'h0;
        src39 <= 16'h0;
        src40 <= 16'h0;
        src41 <= 16'h0;
        src42 <= 16'h0;
        src43 <= 16'h0;
        src44 <= 16'h0;
        src45 <= 16'h0;
        src46 <= 16'h0;
        src47 <= 16'h0;
        src48 <= 16'h0;
        src49 <= 16'h0;
        src50 <= 16'h0;
        src51 <= 16'h0;
        src52 <= 16'h0;
        src53 <= 16'h0;
        src54 <= 16'h0;
        src55 <= 16'h0;
        src56 <= 16'h0;
        src57 <= 16'h0;
        src58 <= 16'h0;
        src59 <= 16'h0;
        src60 <= 16'h0;
        src61 <= 16'h0;
        src62 <= 16'h0;
        src63 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA16_64(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [0:0] comp_out67;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      input wire [15:0] src16,
      input wire [15:0] src17,
      input wire [15:0] src18,
      input wire [15:0] src19,
      input wire [15:0] src20,
      input wire [15:0] src21,
      input wire [15:0] src22,
      input wire [15:0] src23,
      input wire [15:0] src24,
      input wire [15:0] src25,
      input wire [15:0] src26,
      input wire [15:0] src27,
      input wire [15:0] src28,
      input wire [15:0] src29,
      input wire [15:0] src30,
      input wire [15:0] src31,
      input wire [15:0] src32,
      input wire [15:0] src33,
      input wire [15:0] src34,
      input wire [15:0] src35,
      input wire [15:0] src36,
      input wire [15:0] src37,
      input wire [15:0] src38,
      input wire [15:0] src39,
      input wire [15:0] src40,
      input wire [15:0] src41,
      input wire [15:0] src42,
      input wire [15:0] src43,
      input wire [15:0] src44,
      input wire [15:0] src45,
      input wire [15:0] src46,
      input wire [15:0] src47,
      input wire [15:0] src48,
      input wire [15:0] src49,
      input wire [15:0] src50,
      input wire [15:0] src51,
      input wire [15:0] src52,
      input wire [15:0] src53,
      input wire [15:0] src54,
      input wire [15:0] src55,
      input wire [15:0] src56,
      input wire [15:0] src57,
      input wire [15:0] src58,
      input wire [15:0] src59,
      input wire [15:0] src60,
      input wire [15:0] src61,
      input wire [15:0] src62,
      input wire [15:0] src63,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [0:0] dst67);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [15:0] stage0_16;
   wire [15:0] stage0_17;
   wire [15:0] stage0_18;
   wire [15:0] stage0_19;
   wire [15:0] stage0_20;
   wire [15:0] stage0_21;
   wire [15:0] stage0_22;
   wire [15:0] stage0_23;
   wire [15:0] stage0_24;
   wire [15:0] stage0_25;
   wire [15:0] stage0_26;
   wire [15:0] stage0_27;
   wire [15:0] stage0_28;
   wire [15:0] stage0_29;
   wire [15:0] stage0_30;
   wire [15:0] stage0_31;
   wire [15:0] stage0_32;
   wire [15:0] stage0_33;
   wire [15:0] stage0_34;
   wire [15:0] stage0_35;
   wire [15:0] stage0_36;
   wire [15:0] stage0_37;
   wire [15:0] stage0_38;
   wire [15:0] stage0_39;
   wire [15:0] stage0_40;
   wire [15:0] stage0_41;
   wire [15:0] stage0_42;
   wire [15:0] stage0_43;
   wire [15:0] stage0_44;
   wire [15:0] stage0_45;
   wire [15:0] stage0_46;
   wire [15:0] stage0_47;
   wire [15:0] stage0_48;
   wire [15:0] stage0_49;
   wire [15:0] stage0_50;
   wire [15:0] stage0_51;
   wire [15:0] stage0_52;
   wire [15:0] stage0_53;
   wire [15:0] stage0_54;
   wire [15:0] stage0_55;
   wire [15:0] stage0_56;
   wire [15:0] stage0_57;
   wire [15:0] stage0_58;
   wire [15:0] stage0_59;
   wire [15:0] stage0_60;
   wire [15:0] stage0_61;
   wire [15:0] stage0_62;
   wire [15:0] stage0_63;
   wire [10:0] stage1_0;
   wire [6:0] stage1_1;
   wire [8:0] stage1_2;
   wire [6:0] stage1_3;
   wire [5:0] stage1_4;
   wire [7:0] stage1_5;
   wire [6:0] stage1_6;
   wire [5:0] stage1_7;
   wire [9:0] stage1_8;
   wire [5:0] stage1_9;
   wire [9:0] stage1_10;
   wire [6:0] stage1_11;
   wire [5:0] stage1_12;
   wire [9:0] stage1_13;
   wire [6:0] stage1_14;
   wire [6:0] stage1_15;
   wire [5:0] stage1_16;
   wire [14:0] stage1_17;
   wire [5:0] stage1_18;
   wire [11:0] stage1_19;
   wire [7:0] stage1_20;
   wire [5:0] stage1_21;
   wire [6:0] stage1_22;
   wire [5:0] stage1_23;
   wire [7:0] stage1_24;
   wire [6:0] stage1_25;
   wire [8:0] stage1_26;
   wire [6:0] stage1_27;
   wire [5:0] stage1_28;
   wire [6:0] stage1_29;
   wire [9:0] stage1_30;
   wire [7:0] stage1_31;
   wire [8:0] stage1_32;
   wire [8:0] stage1_33;
   wire [5:0] stage1_34;
   wire [7:0] stage1_35;
   wire [6:0] stage1_36;
   wire [8:0] stage1_37;
   wire [5:0] stage1_38;
   wire [5:0] stage1_39;
   wire [6:0] stage1_40;
   wire [9:0] stage1_41;
   wire [6:0] stage1_42;
   wire [5:0] stage1_43;
   wire [7:0] stage1_44;
   wire [6:0] stage1_45;
   wire [5:0] stage1_46;
   wire [7:0] stage1_47;
   wire [7:0] stage1_48;
   wire [6:0] stage1_49;
   wire [6:0] stage1_50;
   wire [8:0] stage1_51;
   wire [5:0] stage1_52;
   wire [13:0] stage1_53;
   wire [5:0] stage1_54;
   wire [5:0] stage1_55;
   wire [6:0] stage1_56;
   wire [9:0] stage1_57;
   wire [7:0] stage1_58;
   wire [7:0] stage1_59;
   wire [6:0] stage1_60;
   wire [5:0] stage1_61;
   wire [6:0] stage1_62;
   wire [13:0] stage1_63;
   wire [3:0] stage1_64;
   wire [0:0] stage1_65;
   wire [5:0] stage2_0;
   wire [2:0] stage2_1;
   wire [4:0] stage2_2;
   wire [2:0] stage2_3;
   wire [2:0] stage2_4;
   wire [4:0] stage2_5;
   wire [2:0] stage2_6;
   wire [1:0] stage2_7;
   wire [5:0] stage2_8;
   wire [2:0] stage2_9;
   wire [7:0] stage2_10;
   wire [1:0] stage2_11;
   wire [1:0] stage2_12;
   wire [6:0] stage2_13;
   wire [3:0] stage2_14;
   wire [2:0] stage2_15;
   wire [1:0] stage2_16;
   wire [6:0] stage2_17;
   wire [4:0] stage2_18;
   wire [2:0] stage2_19;
   wire [4:0] stage2_20;
   wire [4:0] stage2_21;
   wire [2:0] stage2_22;
   wire [1:0] stage2_23;
   wire [5:0] stage2_24;
   wire [2:0] stage2_25;
   wire [6:0] stage2_26;
   wire [1:0] stage2_27;
   wire [1:0] stage2_28;
   wire [2:0] stage2_29;
   wire [3:0] stage2_30;
   wire [3:0] stage2_31;
   wire [5:0] stage2_32;
   wire [2:0] stage2_33;
   wire [2:0] stage2_34;
   wire [3:0] stage2_35;
   wire [2:0] stage2_36;
   wire [5:0] stage2_37;
   wire [5:0] stage2_38;
   wire [1:0] stage2_39;
   wire [1:0] stage2_40;
   wire [6:0] stage2_41;
   wire [2:0] stage2_42;
   wire [1:0] stage2_43;
   wire [5:0] stage2_44;
   wire [2:0] stage2_45;
   wire [3:0] stage2_46;
   wire [1:0] stage2_47;
   wire [2:0] stage2_48;
   wire [6:0] stage2_49;
   wire [3:0] stage2_50;
   wire [2:0] stage2_51;
   wire [5:0] stage2_52;
   wire [4:0] stage2_53;
   wire [2:0] stage2_54;
   wire [3:0] stage2_55;
   wire [1:0] stage2_56;
   wire [6:0] stage2_57;
   wire [4:0] stage2_58;
   wire [2:0] stage2_59;
   wire [3:0] stage2_60;
   wire [1:0] stage2_61;
   wire [2:0] stage2_62;
   wire [9:0] stage2_63;
   wire [3:0] stage2_64;
   wire [1:0] stage2_65;
   wire [0:0] stage2_66;
   wire [1:0] stage3_0;
   wire [0:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [1:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage3_21;
   wire [1:0] stage3_22;
   wire [1:0] stage3_23;
   wire [1:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [1:0] stage3_27;
   wire [1:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [1:0] stage3_31;
   wire [1:0] stage3_32;
   wire [1:0] stage3_33;
   wire [1:0] stage3_34;
   wire [1:0] stage3_35;
   wire [1:0] stage3_36;
   wire [1:0] stage3_37;
   wire [1:0] stage3_38;
   wire [1:0] stage3_39;
   wire [1:0] stage3_40;
   wire [1:0] stage3_41;
   wire [1:0] stage3_42;
   wire [1:0] stage3_43;
   wire [1:0] stage3_44;
   wire [1:0] stage3_45;
   wire [1:0] stage3_46;
   wire [1:0] stage3_47;
   wire [1:0] stage3_48;
   wire [1:0] stage3_49;
   wire [1:0] stage3_50;
   wire [1:0] stage3_51;
   wire [1:0] stage3_52;
   wire [1:0] stage3_53;
   wire [1:0] stage3_54;
   wire [1:0] stage3_55;
   wire [1:0] stage3_56;
   wire [1:0] stage3_57;
   wire [1:0] stage3_58;
   wire [1:0] stage3_59;
   wire [1:0] stage3_60;
   wire [1:0] stage3_61;
   wire [1:0] stage3_62;
   wire [1:0] stage3_63;
   wire [1:0] stage3_64;
   wire [1:0] stage3_65;
   wire [1:0] stage3_66;
   wire [0:0] stage3_67;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;
   assign dst20 = stage3_20;
   assign dst21 = stage3_21;
   assign dst22 = stage3_22;
   assign dst23 = stage3_23;
   assign dst24 = stage3_24;
   assign dst25 = stage3_25;
   assign dst26 = stage3_26;
   assign dst27 = stage3_27;
   assign dst28 = stage3_28;
   assign dst29 = stage3_29;
   assign dst30 = stage3_30;
   assign dst31 = stage3_31;
   assign dst32 = stage3_32;
   assign dst33 = stage3_33;
   assign dst34 = stage3_34;
   assign dst35 = stage3_35;
   assign dst36 = stage3_36;
   assign dst37 = stage3_37;
   assign dst38 = stage3_38;
   assign dst39 = stage3_39;
   assign dst40 = stage3_40;
   assign dst41 = stage3_41;
   assign dst42 = stage3_42;
   assign dst43 = stage3_43;
   assign dst44 = stage3_44;
   assign dst45 = stage3_45;
   assign dst46 = stage3_46;
   assign dst47 = stage3_47;
   assign dst48 = stage3_48;
   assign dst49 = stage3_49;
   assign dst50 = stage3_50;
   assign dst51 = stage3_51;
   assign dst52 = stage3_52;
   assign dst53 = stage3_53;
   assign dst54 = stage3_54;
   assign dst55 = stage3_55;
   assign dst56 = stage3_56;
   assign dst57 = stage3_57;
   assign dst58 = stage3_58;
   assign dst59 = stage3_59;
   assign dst60 = stage3_60;
   assign dst61 = stage3_61;
   assign dst62 = stage3_62;
   assign dst63 = stage3_63;
   assign dst64 = stage3_64;
   assign dst65 = stage3_65;
   assign dst66 = stage3_66;
   assign dst67 = stage3_67;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc615_5 gpc3 (
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage0_3[12]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[3],stage1_3[3],stage1_2[3]}
   );
   gpc615_5 gpc4 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10]},
      {stage0_5[0]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[4]}
   );
   gpc615_5 gpc5 (
      {stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15]},
      {stage0_5[1]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[5]}
   );
   gpc207_4 gpc6 (
      {stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc7 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage1_9[0],stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc1343_5 gpc8 (
      {stage0_6[12], stage0_6[13], stage0_6[14]},
      {stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage0_8[0], stage0_8[1], stage0_8[2]},
      {stage0_9[0]},
      {stage1_10[0],stage1_9[1],stage1_8[4],stage1_7[4],stage1_6[5]}
   );
   gpc1343_5 gpc9 (
      {stage0_6[15], 1'b0, 1'b0},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15]},
      {stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_9[1]},
      {stage1_10[1],stage1_9[2],stage1_8[5],stage1_7[5],stage1_6[6]}
   );
   gpc117_4 gpc10 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[2],stage1_9[3],stage1_8[6]}
   );
   gpc207_4 gpc11 (
      {stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[4]}
   );
   gpc606_5 gpc12 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[0],stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[5]}
   );
   gpc117_4 gpc13 (
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[8]},
      {stage0_12[0]},
      {stage1_13[1],stage1_12[2],stage1_11[3],stage1_10[5]}
   );
   gpc615_5 gpc14 (
      {stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage0_11[9]},
      {stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6]},
      {stage1_14[0],stage1_13[2],stage1_12[3],stage1_11[4],stage1_10[6]}
   );
   gpc135_4 gpc15 (
      {stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14]},
      {stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage0_13[0]},
      {stage1_14[1],stage1_13[3],stage1_12[4],stage1_11[5]}
   );
   gpc606_5 gpc16 (
      {stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[2],stage1_13[4],stage1_12[5]}
   );
   gpc606_5 gpc17 (
      {stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5], stage0_13[6]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[1],stage1_15[1],stage1_14[3],stage1_13[5]}
   );
   gpc606_5 gpc18 (
      {stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[2],stage1_15[2],stage1_14[4],stage1_13[6]}
   );
   gpc615_5 gpc19 (
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10]},
      {stage0_15[12]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[2],stage1_16[3],stage1_15[3],stage1_14[5]}
   );
   gpc615_5 gpc20 (
      {stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage0_15[13]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[3],stage1_16[4],stage1_15[4],stage1_14[6]}
   );
   gpc615_5 gpc21 (
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], 1'b0},
      {stage0_17[0]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[4],stage1_16[5]}
   );
   gpc606_5 gpc22 (
      {stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[5]}
   );
   gpc615_5 gpc23 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10]},
      {stage0_19[6]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[1],stage1_20[2],stage1_19[2],stage1_18[4]}
   );
   gpc615_5 gpc24 (
      {stage0_18[11], stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15]},
      {stage0_19[7]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[2],stage1_20[3],stage1_19[3],stage1_18[5]}
   );
   gpc1343_5 gpc25 (
      {stage0_21[0], stage0_21[1], stage0_21[2]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3]},
      {stage0_23[0], stage0_23[1], stage0_23[2]},
      {stage0_24[0]},
      {stage1_25[0],stage1_24[0],stage1_23[0],stage1_22[2],stage1_21[3]}
   );
   gpc117_4 gpc26 (
      {stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9]},
      {stage0_22[4]},
      {stage0_23[3]},
      {stage1_24[1],stage1_23[1],stage1_22[3],stage1_21[4]}
   );
   gpc606_5 gpc27 (
      {stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[4], stage0_23[5], stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9]},
      {stage1_25[1],stage1_24[2],stage1_23[2],stage1_22[4],stage1_21[5]}
   );
   gpc606_5 gpc28 (
      {stage0_22[5], stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10]},
      {stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6]},
      {stage1_26[0],stage1_25[2],stage1_24[3],stage1_23[3],stage1_22[5]}
   );
   gpc615_5 gpc29 (
      {stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15]},
      {stage0_23[10]},
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage1_26[1],stage1_25[3],stage1_24[4],stage1_23[4],stage1_22[6]}
   );
   gpc615_5 gpc30 (
      {stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage0_24[13]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[2],stage1_25[4],stage1_24[5],stage1_23[5]}
   );
   gpc15_3 gpc31 (
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10]},
      {stage0_26[0]},
      {stage1_27[1],stage1_26[3],stage1_25[5]}
   );
   gpc615_5 gpc32 (
      {stage0_25[11], stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15]},
      {stage0_26[1]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[0],stage1_27[2],stage1_26[4],stage1_25[6]}
   );
   gpc606_5 gpc33 (
      {stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5], stage0_26[6], stage0_26[7]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[1],stage1_28[1],stage1_27[3],stage1_26[5]}
   );
   gpc606_5 gpc34 (
      {stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11], stage0_26[12], stage0_26[13]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[2],stage1_28[2],stage1_27[4],stage1_26[6]}
   );
   gpc615_5 gpc35 (
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10]},
      {stage0_28[12]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[2],stage1_29[3],stage1_28[3],stage1_27[5]}
   );
   gpc615_5 gpc36 (
      {stage0_27[11], stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15]},
      {stage0_28[13]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[3],stage1_29[4],stage1_28[4],stage1_27[6]}
   );
   gpc615_5 gpc37 (
      {stage0_28[14], stage0_28[15], 1'b0, 1'b0, 1'b0},
      {stage0_29[12]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[4],stage1_29[5],stage1_28[5]}
   );
   gpc1163_5 gpc38 (
      {stage0_29[13], stage0_29[14], stage0_29[15]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage0_31[0]},
      {stage0_32[0]},
      {stage1_33[0],stage1_32[1],stage1_31[3],stage1_30[5],stage1_29[6]}
   );
   gpc117_4 gpc39 (
      {stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage0_32[1]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[1],stage1_32[2],stage1_31[4]}
   );
   gpc606_5 gpc40 (
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[1],stage1_33[2],stage1_32[3],stage1_31[5]}
   );
   gpc1406_5 gpc41 (
      {stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5], stage0_32[6], stage0_32[7]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3]},
      {stage0_35[0]},
      {stage1_36[0],stage1_35[1],stage1_34[2],stage1_33[3],stage1_32[4]}
   );
   gpc615_5 gpc42 (
      {stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11], stage0_32[12]},
      {stage0_33[7]},
      {stage0_34[4], stage0_34[5], stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9]},
      {stage1_36[1],stage1_35[2],stage1_34[3],stage1_33[4],stage1_32[5]}
   );
   gpc615_5 gpc43 (
      {stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage0_34[10]},
      {stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5], stage0_35[6]},
      {stage1_37[0],stage1_36[2],stage1_35[3],stage1_34[4],stage1_33[5]}
   );
   gpc615_5 gpc44 (
      {stage0_34[11], stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15]},
      {stage0_35[7]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[1],stage1_36[3],stage1_35[4],stage1_34[5]}
   );
   gpc606_5 gpc45 (
      {stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11], stage0_35[12], stage0_35[13]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[1],stage1_37[2],stage1_36[4],stage1_35[5]}
   );
   gpc615_5 gpc46 (
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10]},
      {stage0_37[6]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[1],stage1_38[2],stage1_37[3],stage1_36[5]}
   );
   gpc615_5 gpc47 (
      {stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15]},
      {stage0_37[7]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[2],stage1_38[3],stage1_37[4],stage1_36[6]}
   );
   gpc615_5 gpc48 (
      {stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12]},
      {stage0_38[12]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[2],stage1_39[3],stage1_38[4],stage1_37[5]}
   );
   gpc1163_5 gpc49 (
      {stage0_38[13], stage0_38[14], stage0_38[15]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage0_40[0]},
      {stage0_41[0]},
      {stage1_42[0],stage1_41[1],stage1_40[3],stage1_39[4],stage1_38[5]}
   );
   gpc135_4 gpc50 (
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], 1'b0},
      {stage0_40[1], stage0_40[2], stage0_40[3]},
      {stage0_41[1]},
      {stage1_42[1],stage1_41[2],stage1_40[4],stage1_39[5]}
   );
   gpc606_5 gpc51 (
      {stage0_40[4], stage0_40[5], stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[0],stage1_42[2],stage1_41[3],stage1_40[5]}
   );
   gpc606_5 gpc52 (
      {stage0_40[10], stage0_40[11], stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[1],stage1_42[3],stage1_41[4],stage1_40[6]}
   );
   gpc135_4 gpc53 (
      {stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5], stage0_41[6]},
      {stage0_42[12], stage0_42[13], stage0_42[14]},
      {stage0_43[0]},
      {stage1_44[2],stage1_43[2],stage1_42[4],stage1_41[5]}
   );
   gpc606_5 gpc54 (
      {stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11], stage0_41[12]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[3],stage1_43[3],stage1_42[5],stage1_41[6]}
   );
   gpc1406_5 gpc55 (
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3]},
      {stage0_46[0]},
      {stage1_47[0],stage1_46[0],stage1_45[1],stage1_44[4],stage1_43[4]}
   );
   gpc1163_5 gpc56 (
      {stage0_43[13], stage0_43[14], stage0_43[15]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage0_45[4]},
      {stage0_46[1]},
      {stage1_47[1],stage1_46[1],stage1_45[2],stage1_44[5],stage1_43[5]}
   );
   gpc615_5 gpc57 (
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10]},
      {stage0_45[5]},
      {stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5], stage0_46[6], stage0_46[7]},
      {stage1_48[0],stage1_47[2],stage1_46[2],stage1_45[3],stage1_44[6]}
   );
   gpc615_5 gpc58 (
      {stage0_44[11], stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15]},
      {stage0_45[6]},
      {stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11], stage0_46[12], stage0_46[13]},
      {stage1_48[1],stage1_47[3],stage1_46[3],stage1_45[4],stage1_44[7]}
   );
   gpc615_5 gpc59 (
      {stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage0_46[14]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[2],stage1_47[4],stage1_46[4],stage1_45[5]}
   );
   gpc615_5 gpc60 (
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], 1'b0},
      {stage0_46[15]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[3],stage1_47[5],stage1_46[5],stage1_45[6]}
   );
   gpc623_5 gpc61 (
      {stage0_47[12], stage0_47[13], stage0_47[14]},
      {stage0_48[0], stage0_48[1]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[0],stage1_49[2],stage1_48[4],stage1_47[6]}
   );
   gpc207_4 gpc62 (
      {stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5], stage0_48[6], stage0_48[7], stage0_48[8]},
      {stage0_50[0], stage0_50[1]},
      {stage1_51[1],stage1_50[1],stage1_49[3],stage1_48[5]}
   );
   gpc606_5 gpc63 (
      {stage0_48[9], stage0_48[10], stage0_48[11], stage0_48[12], stage0_48[13], stage0_48[14]},
      {stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5], stage0_50[6], stage0_50[7]},
      {stage1_52[0],stage1_51[2],stage1_50[2],stage1_49[4],stage1_48[6]}
   );
   gpc615_5 gpc64 (
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10]},
      {stage0_50[8]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[1],stage1_51[3],stage1_50[3],stage1_49[5]}
   );
   gpc615_5 gpc65 (
      {stage0_49[11], stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15]},
      {stage0_50[9]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[2],stage1_51[4],stage1_50[4],stage1_49[6]}
   );
   gpc615_5 gpc66 (
      {stage0_50[10], stage0_50[11], stage0_50[12], stage0_50[13], stage0_50[14]},
      {stage0_51[12]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[2],stage1_52[3],stage1_51[5],stage1_50[5]}
   );
   gpc615_5 gpc67 (
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10]},
      {stage0_53[0]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[0],stage1_54[1],stage1_53[3],stage1_52[4]}
   );
   gpc615_5 gpc68 (
      {stage0_52[11], stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15]},
      {stage0_53[1]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[1],stage1_54[2],stage1_53[4],stage1_52[5]}
   );
   gpc606_5 gpc69 (
      {stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5], stage0_53[6], stage0_53[7]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[2],stage1_55[2],stage1_54[3],stage1_53[5]}
   );
   gpc1343_5 gpc70 (
      {stage0_54[12], stage0_54[13], stage0_54[14]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9]},
      {stage0_56[0], stage0_56[1], stage0_56[2]},
      {stage0_57[0]},
      {stage1_58[0],stage1_57[1],stage1_56[3],stage1_55[3],stage1_54[4]}
   );
   gpc615_5 gpc71 (
      {stage0_55[10], stage0_55[11], stage0_55[12], stage0_55[13], stage0_55[14]},
      {stage0_56[3]},
      {stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6]},
      {stage1_59[0],stage1_58[1],stage1_57[2],stage1_56[4],stage1_55[4]}
   );
   gpc606_5 gpc72 (
      {stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[1],stage1_58[2],stage1_57[3],stage1_56[5]}
   );
   gpc606_5 gpc73 (
      {stage0_56[10], stage0_56[11], stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[2],stage1_58[3],stage1_57[4],stage1_56[6]}
   );
   gpc615_5 gpc74 (
      {stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage0_58[12]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[2],stage1_59[3],stage1_58[4],stage1_57[5]}
   );
   gpc1343_5 gpc75 (
      {stage0_59[6], stage0_59[7], stage0_59[8]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3]},
      {stage0_61[0], stage0_61[1], stage0_61[2]},
      {stage0_62[0]},
      {stage1_63[0],stage1_62[0],stage1_61[1],stage1_60[3],stage1_59[4]}
   );
   gpc615_5 gpc76 (
      {stage0_59[9], stage0_59[10], stage0_59[11], stage0_59[12], stage0_59[13]},
      {stage0_60[4]},
      {stage0_61[3], stage0_61[4], stage0_61[5], stage0_61[6], stage0_61[7], stage0_61[8]},
      {stage1_63[1],stage1_62[1],stage1_61[2],stage1_60[4],stage1_59[5]}
   );
   gpc606_5 gpc77 (
      {stage0_60[5], stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10]},
      {stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5], stage0_62[6]},
      {stage1_64[0],stage1_63[2],stage1_62[2],stage1_61[3],stage1_60[5]}
   );
   gpc615_5 gpc78 (
      {stage0_60[11], stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15]},
      {stage0_61[9]},
      {stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11], stage0_62[12]},
      {stage1_64[1],stage1_63[3],stage1_62[3],stage1_61[4],stage1_60[6]}
   );
   gpc117_4 gpc79 (
      {stage0_61[10], stage0_61[11], stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], 1'b0},
      {stage0_62[13]},
      {stage0_63[0]},
      {stage1_64[2],stage1_63[4],stage1_62[4],stage1_61[5]}
   );
   gpc7_3 gpc80 (
      {stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5], stage0_63[6], stage0_63[7]},
      {stage1_65[0],stage1_64[3],stage1_63[5]}
   );
   gpc1_1 gpc81 (
      {stage0_0[6]},
      {stage1_0[1]}
   );
   gpc1_1 gpc82 (
      {stage0_0[7]},
      {stage1_0[2]}
   );
   gpc1_1 gpc83 (
      {stage0_0[8]},
      {stage1_0[3]}
   );
   gpc1_1 gpc84 (
      {stage0_0[9]},
      {stage1_0[4]}
   );
   gpc1_1 gpc85 (
      {stage0_0[10]},
      {stage1_0[5]}
   );
   gpc1_1 gpc86 (
      {stage0_0[11]},
      {stage1_0[6]}
   );
   gpc1_1 gpc87 (
      {stage0_0[12]},
      {stage1_0[7]}
   );
   gpc1_1 gpc88 (
      {stage0_0[13]},
      {stage1_0[8]}
   );
   gpc1_1 gpc89 (
      {stage0_0[14]},
      {stage1_0[9]}
   );
   gpc1_1 gpc90 (
      {stage0_0[15]},
      {stage1_0[10]}
   );
   gpc1_1 gpc91 (
      {stage0_1[12]},
      {stage1_1[3]}
   );
   gpc1_1 gpc92 (
      {stage0_1[13]},
      {stage1_1[4]}
   );
   gpc1_1 gpc93 (
      {stage0_1[14]},
      {stage1_1[5]}
   );
   gpc1_1 gpc94 (
      {stage0_1[15]},
      {stage1_1[6]}
   );
   gpc1_1 gpc95 (
      {stage0_2[11]},
      {stage1_2[4]}
   );
   gpc1_1 gpc96 (
      {stage0_2[12]},
      {stage1_2[5]}
   );
   gpc1_1 gpc97 (
      {stage0_2[13]},
      {stage1_2[6]}
   );
   gpc1_1 gpc98 (
      {stage0_2[14]},
      {stage1_2[7]}
   );
   gpc1_1 gpc99 (
      {stage0_2[15]},
      {stage1_2[8]}
   );
   gpc1_1 gpc100 (
      {stage0_3[13]},
      {stage1_3[4]}
   );
   gpc1_1 gpc101 (
      {stage0_3[14]},
      {stage1_3[5]}
   );
   gpc1_1 gpc102 (
      {stage0_3[15]},
      {stage1_3[6]}
   );
   gpc1_1 gpc103 (
      {stage0_5[15]},
      {stage1_5[7]}
   );
   gpc1_1 gpc104 (
      {stage0_8[13]},
      {stage1_8[7]}
   );
   gpc1_1 gpc105 (
      {stage0_8[14]},
      {stage1_8[8]}
   );
   gpc1_1 gpc106 (
      {stage0_8[15]},
      {stage1_8[9]}
   );
   gpc1_1 gpc107 (
      {stage0_10[13]},
      {stage1_10[7]}
   );
   gpc1_1 gpc108 (
      {stage0_10[14]},
      {stage1_10[8]}
   );
   gpc1_1 gpc109 (
      {stage0_10[15]},
      {stage1_10[9]}
   );
   gpc1_1 gpc110 (
      {stage0_11[15]},
      {stage1_11[6]}
   );
   gpc1_1 gpc111 (
      {stage0_13[13]},
      {stage1_13[7]}
   );
   gpc1_1 gpc112 (
      {stage0_13[14]},
      {stage1_13[8]}
   );
   gpc1_1 gpc113 (
      {stage0_13[15]},
      {stage1_13[9]}
   );
   gpc1_1 gpc114 (
      {stage0_15[14]},
      {stage1_15[5]}
   );
   gpc1_1 gpc115 (
      {stage0_15[15]},
      {stage1_15[6]}
   );
   gpc1_1 gpc116 (
      {stage0_17[7]},
      {stage1_17[6]}
   );
   gpc1_1 gpc117 (
      {stage0_17[8]},
      {stage1_17[7]}
   );
   gpc1_1 gpc118 (
      {stage0_17[9]},
      {stage1_17[8]}
   );
   gpc1_1 gpc119 (
      {stage0_17[10]},
      {stage1_17[9]}
   );
   gpc1_1 gpc120 (
      {stage0_17[11]},
      {stage1_17[10]}
   );
   gpc1_1 gpc121 (
      {stage0_17[12]},
      {stage1_17[11]}
   );
   gpc1_1 gpc122 (
      {stage0_17[13]},
      {stage1_17[12]}
   );
   gpc1_1 gpc123 (
      {stage0_17[14]},
      {stage1_17[13]}
   );
   gpc1_1 gpc124 (
      {stage0_17[15]},
      {stage1_17[14]}
   );
   gpc1_1 gpc125 (
      {stage0_19[8]},
      {stage1_19[4]}
   );
   gpc1_1 gpc126 (
      {stage0_19[9]},
      {stage1_19[5]}
   );
   gpc1_1 gpc127 (
      {stage0_19[10]},
      {stage1_19[6]}
   );
   gpc1_1 gpc128 (
      {stage0_19[11]},
      {stage1_19[7]}
   );
   gpc1_1 gpc129 (
      {stage0_19[12]},
      {stage1_19[8]}
   );
   gpc1_1 gpc130 (
      {stage0_19[13]},
      {stage1_19[9]}
   );
   gpc1_1 gpc131 (
      {stage0_19[14]},
      {stage1_19[10]}
   );
   gpc1_1 gpc132 (
      {stage0_19[15]},
      {stage1_19[11]}
   );
   gpc1_1 gpc133 (
      {stage0_20[12]},
      {stage1_20[4]}
   );
   gpc1_1 gpc134 (
      {stage0_20[13]},
      {stage1_20[5]}
   );
   gpc1_1 gpc135 (
      {stage0_20[14]},
      {stage1_20[6]}
   );
   gpc1_1 gpc136 (
      {stage0_20[15]},
      {stage1_20[7]}
   );
   gpc1_1 gpc137 (
      {stage0_24[14]},
      {stage1_24[6]}
   );
   gpc1_1 gpc138 (
      {stage0_24[15]},
      {stage1_24[7]}
   );
   gpc1_1 gpc139 (
      {stage0_26[14]},
      {stage1_26[7]}
   );
   gpc1_1 gpc140 (
      {stage0_26[15]},
      {stage1_26[8]}
   );
   gpc1_1 gpc141 (
      {stage0_30[12]},
      {stage1_30[6]}
   );
   gpc1_1 gpc142 (
      {stage0_30[13]},
      {stage1_30[7]}
   );
   gpc1_1 gpc143 (
      {stage0_30[14]},
      {stage1_30[8]}
   );
   gpc1_1 gpc144 (
      {stage0_30[15]},
      {stage1_30[9]}
   );
   gpc1_1 gpc145 (
      {stage0_31[14]},
      {stage1_31[6]}
   );
   gpc1_1 gpc146 (
      {stage0_31[15]},
      {stage1_31[7]}
   );
   gpc1_1 gpc147 (
      {stage0_32[13]},
      {stage1_32[6]}
   );
   gpc1_1 gpc148 (
      {stage0_32[14]},
      {stage1_32[7]}
   );
   gpc1_1 gpc149 (
      {stage0_32[15]},
      {stage1_32[8]}
   );
   gpc1_1 gpc150 (
      {stage0_33[13]},
      {stage1_33[6]}
   );
   gpc1_1 gpc151 (
      {stage0_33[14]},
      {stage1_33[7]}
   );
   gpc1_1 gpc152 (
      {stage0_33[15]},
      {stage1_33[8]}
   );
   gpc1_1 gpc153 (
      {stage0_35[14]},
      {stage1_35[6]}
   );
   gpc1_1 gpc154 (
      {stage0_35[15]},
      {stage1_35[7]}
   );
   gpc1_1 gpc155 (
      {stage0_37[13]},
      {stage1_37[6]}
   );
   gpc1_1 gpc156 (
      {stage0_37[14]},
      {stage1_37[7]}
   );
   gpc1_1 gpc157 (
      {stage0_37[15]},
      {stage1_37[8]}
   );
   gpc1_1 gpc158 (
      {stage0_41[13]},
      {stage1_41[7]}
   );
   gpc1_1 gpc159 (
      {stage0_41[14]},
      {stage1_41[8]}
   );
   gpc1_1 gpc160 (
      {stage0_41[15]},
      {stage1_41[9]}
   );
   gpc1_1 gpc161 (
      {stage0_42[15]},
      {stage1_42[6]}
   );
   gpc1_1 gpc162 (
      {stage0_47[15]},
      {stage1_47[7]}
   );
   gpc1_1 gpc163 (
      {stage0_48[15]},
      {stage1_48[7]}
   );
   gpc1_1 gpc164 (
      {stage0_50[15]},
      {stage1_50[6]}
   );
   gpc1_1 gpc165 (
      {stage0_51[13]},
      {stage1_51[6]}
   );
   gpc1_1 gpc166 (
      {stage0_51[14]},
      {stage1_51[7]}
   );
   gpc1_1 gpc167 (
      {stage0_51[15]},
      {stage1_51[8]}
   );
   gpc1_1 gpc168 (
      {stage0_53[8]},
      {stage1_53[6]}
   );
   gpc1_1 gpc169 (
      {stage0_53[9]},
      {stage1_53[7]}
   );
   gpc1_1 gpc170 (
      {stage0_53[10]},
      {stage1_53[8]}
   );
   gpc1_1 gpc171 (
      {stage0_53[11]},
      {stage1_53[9]}
   );
   gpc1_1 gpc172 (
      {stage0_53[12]},
      {stage1_53[10]}
   );
   gpc1_1 gpc173 (
      {stage0_53[13]},
      {stage1_53[11]}
   );
   gpc1_1 gpc174 (
      {stage0_53[14]},
      {stage1_53[12]}
   );
   gpc1_1 gpc175 (
      {stage0_53[15]},
      {stage1_53[13]}
   );
   gpc1_1 gpc176 (
      {stage0_54[15]},
      {stage1_54[5]}
   );
   gpc1_1 gpc177 (
      {stage0_55[15]},
      {stage1_55[5]}
   );
   gpc1_1 gpc178 (
      {stage0_57[12]},
      {stage1_57[6]}
   );
   gpc1_1 gpc179 (
      {stage0_57[13]},
      {stage1_57[7]}
   );
   gpc1_1 gpc180 (
      {stage0_57[14]},
      {stage1_57[8]}
   );
   gpc1_1 gpc181 (
      {stage0_57[15]},
      {stage1_57[9]}
   );
   gpc1_1 gpc182 (
      {stage0_58[13]},
      {stage1_58[5]}
   );
   gpc1_1 gpc183 (
      {stage0_58[14]},
      {stage1_58[6]}
   );
   gpc1_1 gpc184 (
      {stage0_58[15]},
      {stage1_58[7]}
   );
   gpc1_1 gpc185 (
      {stage0_59[14]},
      {stage1_59[6]}
   );
   gpc1_1 gpc186 (
      {stage0_59[15]},
      {stage1_59[7]}
   );
   gpc1_1 gpc187 (
      {stage0_62[14]},
      {stage1_62[5]}
   );
   gpc1_1 gpc188 (
      {stage0_62[15]},
      {stage1_62[6]}
   );
   gpc1_1 gpc189 (
      {stage0_63[8]},
      {stage1_63[6]}
   );
   gpc1_1 gpc190 (
      {stage0_63[9]},
      {stage1_63[7]}
   );
   gpc1_1 gpc191 (
      {stage0_63[10]},
      {stage1_63[8]}
   );
   gpc1_1 gpc192 (
      {stage0_63[11]},
      {stage1_63[9]}
   );
   gpc1_1 gpc193 (
      {stage0_63[12]},
      {stage1_63[10]}
   );
   gpc1_1 gpc194 (
      {stage0_63[13]},
      {stage1_63[11]}
   );
   gpc1_1 gpc195 (
      {stage0_63[14]},
      {stage1_63[12]}
   );
   gpc1_1 gpc196 (
      {stage0_63[15]},
      {stage1_63[13]}
   );
   gpc606_5 gpc197 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc198 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc199 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc200 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc7_3 gpc201 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6]},
      {stage2_10[0],stage2_9[1],stage2_8[2]}
   );
   gpc606_5 gpc202 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1],stage2_9[2]}
   );
   gpc615_5 gpc203 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[2]}
   );
   gpc606_5 gpc204 (
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[2]}
   );
   gpc606_5 gpc205 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[1],stage2_14[2]}
   );
   gpc606_5 gpc206 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[0],stage2_19[0],stage2_18[1],stage2_17[2]}
   );
   gpc606_5 gpc207 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[1],stage2_19[1],stage2_18[2],stage2_17[3]}
   );
   gpc615_5 gpc208 (
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4]},
      {1'b0},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[2],stage2_19[2],stage2_18[3]}
   );
   gpc615_5 gpc209 (
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4]},
      {stage1_22[0]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[3]}
   );
   gpc1406_5 gpc210 (
      {stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5], stage1_22[6]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2]}
   );
   gpc606_5 gpc211 (
      {stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[0],stage2_27[0],stage2_26[1],stage2_25[2]}
   );
   gpc615_5 gpc212 (
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4]},
      {stage1_27[6]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[1],stage2_28[1],stage2_27[1],stage2_26[2]}
   );
   gpc7_3 gpc213 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5], stage1_29[6]},
      {stage2_31[0],stage2_30[1],stage2_29[2]}
   );
   gpc7_3 gpc214 (
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6]},
      {stage2_32[0],stage2_31[1],stage2_30[2]}
   );
   gpc623_5 gpc215 (
      {stage1_30[7], stage1_30[8], stage1_30[9]},
      {stage1_31[0], stage1_31[1]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[0],stage2_32[1],stage2_31[2],stage2_30[3]}
   );
   gpc606_5 gpc216 (
      {stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[1],stage2_33[1],stage2_32[2],stage2_31[3]}
   );
   gpc1163_5 gpc217 (
      {stage1_33[6], stage1_33[7], stage1_33[8]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage1_35[0]},
      {stage1_36[0]},
      {stage2_37[0],stage2_36[0],stage2_35[1],stage2_34[2],stage2_33[2]}
   );
   gpc606_5 gpc218 (
      {stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[0],stage2_37[1],stage2_36[1],stage2_35[2]}
   );
   gpc7_3 gpc219 (
      {stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5], stage1_36[6], 1'b0},
      {stage2_38[1],stage2_37[2],stage2_36[2]}
   );
   gpc1163_5 gpc220 (
      {stage1_38[0], stage1_38[1], stage1_38[2]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage1_40[0]},
      {stage1_41[0]},
      {stage2_42[0],stage2_41[0],stage2_40[0],stage2_39[1],stage2_38[2]}
   );
   gpc606_5 gpc221 (
      {stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5], stage1_40[6]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[1],stage2_41[1],stage2_40[1]}
   );
   gpc615_5 gpc222 (
      {stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_42[6]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[1],stage2_43[1],stage2_42[2],stage2_41[2]}
   );
   gpc15_3 gpc223 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[0]},
      {stage2_46[0],stage2_45[1],stage2_44[2]}
   );
   gpc606_5 gpc224 (
      {stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5], stage1_45[6]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[0],stage2_46[1],stage2_45[2]}
   );
   gpc1325_5 gpc225 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4]},
      {stage1_47[6], stage1_47[7]},
      {stage1_48[0], stage1_48[1], stage1_48[2]},
      {stage1_49[0]},
      {stage2_50[0],stage2_49[1],stage2_48[1],stage2_47[1],stage2_46[2]}
   );
   gpc7_3 gpc226 (
      {stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6], stage1_48[7], 1'b0, 1'b0},
      {stage2_50[1],stage2_49[2],stage2_48[2]}
   );
   gpc1163_5 gpc227 (
      {stage1_49[1], stage1_49[2], stage1_49[3]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage1_51[0]},
      {stage1_52[0]},
      {stage2_53[0],stage2_52[0],stage2_51[0],stage2_50[2],stage2_49[3]}
   );
   gpc615_5 gpc228 (
      {stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[1]},
      {stage1_53[0], stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage2_55[0],stage2_54[0],stage2_53[1],stage2_52[1],stage2_51[1]}
   );
   gpc615_5 gpc229 (
      {stage1_51[6], stage1_51[7], stage1_51[8], 1'b0, 1'b0},
      {stage1_52[2]},
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage2_55[1],stage2_54[1],stage2_53[2],stage2_52[2],stage2_51[2]}
   );
   gpc606_5 gpc230 (
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[0],stage2_56[0],stage2_55[2],stage2_54[2]}
   );
   gpc117_4 gpc231 (
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5], 1'b0},
      {stage1_56[6]},
      {stage1_57[0]},
      {stage2_58[1],stage2_57[1],stage2_56[1],stage2_55[3]}
   );
   gpc215_4 gpc232 (
      {stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage1_58[0]},
      {stage1_59[0], stage1_59[1]},
      {stage2_60[0],stage2_59[0],stage2_58[2],stage2_57[2]}
   );
   gpc606_5 gpc233 (
      {stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5], stage1_58[6]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[0],stage2_60[1],stage2_59[1],stage2_58[3]}
   );
   gpc606_5 gpc234 (
      {stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5], stage1_59[6], stage1_59[7]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[1],stage2_61[1],stage2_60[2],stage2_59[2]}
   );
   gpc207_4 gpc235 (
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5], stage1_62[6]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[0],stage2_64[0],stage2_63[1],stage2_62[2]}
   );
   gpc207_4 gpc236 (
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6]},
      {stage1_65[0], 1'b0},
      {stage2_66[0],stage2_65[1],stage2_64[1],stage2_63[2]}
   );
   gpc1_1 gpc237 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc238 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc239 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc240 (
      {stage1_0[9]},
      {stage2_0[4]}
   );
   gpc1_1 gpc241 (
      {stage1_0[10]},
      {stage2_0[5]}
   );
   gpc1_1 gpc242 (
      {stage1_1[6]},
      {stage2_1[2]}
   );
   gpc1_1 gpc243 (
      {stage1_2[6]},
      {stage2_2[2]}
   );
   gpc1_1 gpc244 (
      {stage1_2[7]},
      {stage2_2[3]}
   );
   gpc1_1 gpc245 (
      {stage1_2[8]},
      {stage2_2[4]}
   );
   gpc1_1 gpc246 (
      {stage1_3[6]},
      {stage2_3[2]}
   );
   gpc1_1 gpc247 (
      {stage1_5[6]},
      {stage2_5[3]}
   );
   gpc1_1 gpc248 (
      {stage1_5[7]},
      {stage2_5[4]}
   );
   gpc1_1 gpc249 (
      {stage1_6[6]},
      {stage2_6[2]}
   );
   gpc1_1 gpc250 (
      {stage1_8[7]},
      {stage2_8[3]}
   );
   gpc1_1 gpc251 (
      {stage1_8[8]},
      {stage2_8[4]}
   );
   gpc1_1 gpc252 (
      {stage1_8[9]},
      {stage2_8[5]}
   );
   gpc1_1 gpc253 (
      {stage1_10[5]},
      {stage2_10[3]}
   );
   gpc1_1 gpc254 (
      {stage1_10[6]},
      {stage2_10[4]}
   );
   gpc1_1 gpc255 (
      {stage1_10[7]},
      {stage2_10[5]}
   );
   gpc1_1 gpc256 (
      {stage1_10[8]},
      {stage2_10[6]}
   );
   gpc1_1 gpc257 (
      {stage1_10[9]},
      {stage2_10[7]}
   );
   gpc1_1 gpc258 (
      {stage1_13[6]},
      {stage2_13[3]}
   );
   gpc1_1 gpc259 (
      {stage1_13[7]},
      {stage2_13[4]}
   );
   gpc1_1 gpc260 (
      {stage1_13[8]},
      {stage2_13[5]}
   );
   gpc1_1 gpc261 (
      {stage1_13[9]},
      {stage2_13[6]}
   );
   gpc1_1 gpc262 (
      {stage1_14[6]},
      {stage2_14[3]}
   );
   gpc1_1 gpc263 (
      {stage1_15[6]},
      {stage2_15[2]}
   );
   gpc1_1 gpc264 (
      {stage1_17[12]},
      {stage2_17[4]}
   );
   gpc1_1 gpc265 (
      {stage1_17[13]},
      {stage2_17[5]}
   );
   gpc1_1 gpc266 (
      {stage1_17[14]},
      {stage2_17[6]}
   );
   gpc1_1 gpc267 (
      {stage1_18[5]},
      {stage2_18[4]}
   );
   gpc1_1 gpc268 (
      {stage1_20[6]},
      {stage2_20[3]}
   );
   gpc1_1 gpc269 (
      {stage1_20[7]},
      {stage2_20[4]}
   );
   gpc1_1 gpc270 (
      {stage1_21[5]},
      {stage2_21[4]}
   );
   gpc1_1 gpc271 (
      {stage1_24[4]},
      {stage2_24[2]}
   );
   gpc1_1 gpc272 (
      {stage1_24[5]},
      {stage2_24[3]}
   );
   gpc1_1 gpc273 (
      {stage1_24[6]},
      {stage2_24[4]}
   );
   gpc1_1 gpc274 (
      {stage1_24[7]},
      {stage2_24[5]}
   );
   gpc1_1 gpc275 (
      {stage1_26[5]},
      {stage2_26[3]}
   );
   gpc1_1 gpc276 (
      {stage1_26[6]},
      {stage2_26[4]}
   );
   gpc1_1 gpc277 (
      {stage1_26[7]},
      {stage2_26[5]}
   );
   gpc1_1 gpc278 (
      {stage1_26[8]},
      {stage2_26[6]}
   );
   gpc1_1 gpc279 (
      {stage1_32[6]},
      {stage2_32[3]}
   );
   gpc1_1 gpc280 (
      {stage1_32[7]},
      {stage2_32[4]}
   );
   gpc1_1 gpc281 (
      {stage1_32[8]},
      {stage2_32[5]}
   );
   gpc1_1 gpc282 (
      {stage1_35[7]},
      {stage2_35[3]}
   );
   gpc1_1 gpc283 (
      {stage1_37[6]},
      {stage2_37[3]}
   );
   gpc1_1 gpc284 (
      {stage1_37[7]},
      {stage2_37[4]}
   );
   gpc1_1 gpc285 (
      {stage1_37[8]},
      {stage2_37[5]}
   );
   gpc1_1 gpc286 (
      {stage1_38[3]},
      {stage2_38[3]}
   );
   gpc1_1 gpc287 (
      {stage1_38[4]},
      {stage2_38[4]}
   );
   gpc1_1 gpc288 (
      {stage1_38[5]},
      {stage2_38[5]}
   );
   gpc1_1 gpc289 (
      {stage1_41[6]},
      {stage2_41[3]}
   );
   gpc1_1 gpc290 (
      {stage1_41[7]},
      {stage2_41[4]}
   );
   gpc1_1 gpc291 (
      {stage1_41[8]},
      {stage2_41[5]}
   );
   gpc1_1 gpc292 (
      {stage1_41[9]},
      {stage2_41[6]}
   );
   gpc1_1 gpc293 (
      {stage1_44[5]},
      {stage2_44[3]}
   );
   gpc1_1 gpc294 (
      {stage1_44[6]},
      {stage2_44[4]}
   );
   gpc1_1 gpc295 (
      {stage1_44[7]},
      {stage2_44[5]}
   );
   gpc1_1 gpc296 (
      {stage1_46[5]},
      {stage2_46[3]}
   );
   gpc1_1 gpc297 (
      {stage1_49[4]},
      {stage2_49[4]}
   );
   gpc1_1 gpc298 (
      {stage1_49[5]},
      {stage2_49[5]}
   );
   gpc1_1 gpc299 (
      {stage1_49[6]},
      {stage2_49[6]}
   );
   gpc1_1 gpc300 (
      {stage1_50[6]},
      {stage2_50[3]}
   );
   gpc1_1 gpc301 (
      {stage1_52[3]},
      {stage2_52[3]}
   );
   gpc1_1 gpc302 (
      {stage1_52[4]},
      {stage2_52[4]}
   );
   gpc1_1 gpc303 (
      {stage1_52[5]},
      {stage2_52[5]}
   );
   gpc1_1 gpc304 (
      {stage1_53[12]},
      {stage2_53[3]}
   );
   gpc1_1 gpc305 (
      {stage1_53[13]},
      {stage2_53[4]}
   );
   gpc1_1 gpc306 (
      {stage1_57[6]},
      {stage2_57[3]}
   );
   gpc1_1 gpc307 (
      {stage1_57[7]},
      {stage2_57[4]}
   );
   gpc1_1 gpc308 (
      {stage1_57[8]},
      {stage2_57[5]}
   );
   gpc1_1 gpc309 (
      {stage1_57[9]},
      {stage2_57[6]}
   );
   gpc1_1 gpc310 (
      {stage1_58[7]},
      {stage2_58[4]}
   );
   gpc1_1 gpc311 (
      {stage1_60[6]},
      {stage2_60[3]}
   );
   gpc1_1 gpc312 (
      {stage1_63[7]},
      {stage2_63[3]}
   );
   gpc1_1 gpc313 (
      {stage1_63[8]},
      {stage2_63[4]}
   );
   gpc1_1 gpc314 (
      {stage1_63[9]},
      {stage2_63[5]}
   );
   gpc1_1 gpc315 (
      {stage1_63[10]},
      {stage2_63[6]}
   );
   gpc1_1 gpc316 (
      {stage1_63[11]},
      {stage2_63[7]}
   );
   gpc1_1 gpc317 (
      {stage1_63[12]},
      {stage2_63[8]}
   );
   gpc1_1 gpc318 (
      {stage1_63[13]},
      {stage2_63[9]}
   );
   gpc1_1 gpc319 (
      {stage1_64[2]},
      {stage2_64[2]}
   );
   gpc1_1 gpc320 (
      {stage1_64[3]},
      {stage2_64[3]}
   );
   gpc2135_5 gpc321 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc322 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], 1'b0},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], 1'b0, 1'b0, 1'b0},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc135_4 gpc323 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4]},
      {stage2_6[0], stage2_6[1], stage2_6[2]},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc606_5 gpc324 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1]}
   );
   gpc2223_5 gpc325 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[6], stage2_10[7]},
      {stage2_11[0], stage2_11[1]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[0],stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[1]}
   );
   gpc7_3 gpc326 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[0],stage3_14[0],stage3_13[1]}
   );
   gpc135_4 gpc327 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], 1'b0},
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[0]},
      {stage3_17[0],stage3_16[0],stage3_15[1],stage3_14[1]}
   );
   gpc207_4 gpc328 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage2_19[0], stage2_19[1]},
      {stage3_20[0],stage3_19[0],stage3_18[0],stage3_17[1]}
   );
   gpc615_5 gpc329 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[2]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], 1'b0},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[1],stage3_18[1]}
   );
   gpc2135_5 gpc330 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4]},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage2_24[0], stage2_24[1]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[1],stage3_21[1]}
   );
   gpc2135_5 gpc331 (
      {stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], 1'b0},
      {stage2_25[0], stage2_25[1], stage2_25[2]},
      {stage2_26[0]},
      {stage2_27[0], stage2_27[1]},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[1],stage3_24[1]}
   );
   gpc207_4 gpc332 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6], 1'b0},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1]}
   );
   gpc3_2 gpc333 (
      {stage2_29[0], stage2_29[1], stage2_29[2]},
      {stage3_30[0],stage3_29[1]}
   );
   gpc15_3 gpc334 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], 1'b0},
      {stage2_31[0]},
      {stage3_32[0],stage3_31[0],stage3_30[1]}
   );
   gpc1163_5 gpc335 (
      {stage2_31[1], stage2_31[2], stage2_31[3]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage2_33[0]},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[1]}
   );
   gpc623_5 gpc336 (
      {stage2_33[1], stage2_33[2], 1'b0},
      {stage2_34[1], stage2_34[2]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], 1'b0, 1'b0},
      {stage3_37[0],stage3_36[0],stage3_35[1],stage3_34[1],stage3_33[1]}
   );
   gpc1163_5 gpc337 (
      {stage2_36[0], stage2_36[1], stage2_36[2]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage2_38[0]},
      {stage2_39[0]},
      {stage3_40[0],stage3_39[0],stage3_38[0],stage3_37[1],stage3_36[1]}
   );
   gpc215_4 gpc338 (
      {stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage2_39[1]},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[0],stage3_40[1],stage3_39[1],stage3_38[1]}
   );
   gpc207_4 gpc339 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5], stage2_41[6]},
      {stage2_43[0], stage2_43[1]},
      {stage3_44[0],stage3_43[0],stage3_42[0],stage3_41[1]}
   );
   gpc3_2 gpc340 (
      {stage2_42[0], stage2_42[1], stage2_42[2]},
      {stage3_43[1],stage3_42[1]}
   );
   gpc207_4 gpc341 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5], 1'b0},
      {stage2_46[0], stage2_46[1]},
      {stage3_47[0],stage3_46[0],stage3_45[0],stage3_44[1]}
   );
   gpc2223_5 gpc342 (
      {stage2_45[0], stage2_45[1], stage2_45[2]},
      {stage2_46[2], stage2_46[3]},
      {stage2_47[0], stage2_47[1]},
      {stage2_48[0], stage2_48[1]},
      {stage3_49[0],stage3_48[0],stage3_47[1],stage3_46[1],stage3_45[1]}
   );
   gpc117_4 gpc343 (
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6]},
      {stage2_50[0]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[0],stage3_50[0],stage3_49[1]}
   );
   gpc623_5 gpc344 (
      {stage2_50[1], stage2_50[2], stage2_50[3]},
      {stage2_51[1], stage2_51[2]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[0],stage3_52[1],stage3_51[1],stage3_50[1]}
   );
   gpc135_4 gpc345 (
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4]},
      {stage2_54[0], stage2_54[1], stage2_54[2]},
      {stage2_55[0]},
      {stage3_56[0],stage3_55[0],stage3_54[1],stage3_53[1]}
   );
   gpc23_3 gpc346 (
      {stage2_55[1], stage2_55[2], stage2_55[3]},
      {stage2_56[0], stage2_56[1]},
      {stage3_57[0],stage3_56[1],stage3_55[1]}
   );
   gpc207_4 gpc347 (
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6]},
      {stage2_59[0], stage2_59[1]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[1]}
   );
   gpc1415_5 gpc348 (
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4]},
      {stage2_59[2]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[0],stage3_60[1],stage3_59[1],stage3_58[1]}
   );
   gpc1163_5 gpc349 (
      {stage2_62[0], stage2_62[1], stage2_62[2]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage2_64[0]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[0],stage3_64[0],stage3_63[0],stage3_62[1]}
   );
   gpc2135_5 gpc350 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], 1'b0},
      {stage2_64[1], stage2_64[2], stage2_64[3]},
      {stage2_65[1]},
      {stage2_66[0], 1'b0},
      {stage3_67[0],stage3_66[1],stage3_65[1],stage3_64[1],stage3_63[1]}
   );
   gpc1_1 gpc351 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc352 (
      {stage2_7[1]},
      {stage3_7[1]}
   );
   gpc1_1 gpc353 (
      {stage2_16[1]},
      {stage3_16[1]}
   );
   gpc1_1 gpc354 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc355 (
      {stage2_48[2]},
      {stage3_48[1]}
   );
   gpc1_1 gpc356 (
      {stage2_61[1]},
      {stage3_61[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [67:0] srcsum;
    wire [67:0] dstsum;
    wire test;
    compressor_CLA16_64 compressor_CLA16_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8fa1acf0f874f7491032087f8a723d8d173d1ef79b7ed276492a0b1050dc97e5d2f3768f7dd79e0d69dbed634928d100f69dc119051b60db22e85606c53fbd2a9c8c69ee9a1a9fbb0e3802c7db62db3d0ff41cf38caced8807ff0c15f72df233047f4b89ca850ec605abe4024f8774395cdb5c6f4b8e807f5b99e42fd40b9d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h536af076645148ee16057b35b3d7398616dca57e386e72d365e6da1bb8ed40db74009f03d4414e7a165580c2bcbe2b2da2a90aeb96c3f08cffa7653e2c7ccd2a1cd1e98d869aaca402e6d65b44ef14ddf47d2c7e6745d6da34b643e0602357a7446a5db53b9b537decedd0e26f35ce5f95330ec6592c0b18062902b95ed4e690;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h885f2313cb788cdfbcca35817558c88eb4fa40244e225840ba57f80475cd48a907d8403094973e94acd76541caf86ee91515a0c62bff806a84a42f534dc9e3fac19da97ee7d1f1df618fb5722806c83906ca98ba7ce567c19329eedb07625087823332c7d9674b8c732a7655a460dc321c8ca2a006d5161ca7061b365985a18d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46b4e16c050ef5925553a1aec9b57b0466a4e7dbc7b9556861dc33e1a5c6593c1589e9c360836f0b6fd72d28f928ea7f4a000c389021ef13303ddd6f8debf0e35124a9972217b262a93ad3ac483fda262efba73fdc3c2c5459239f8a60243993919c47d54049c7750dbab8f37a4e1bf079932ffb26f83641935d5944a0f5b377;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9817a3fdf963ca953470a1344a59e1fc8c5cb91a94253fe93f7a39c82be08a8a97c55ed56c8ee899689b4e8b2aa3babac65a48edff80ec45bdd9141aaf8736fc74fed5365dc5a91b9253e36a58ab08e03e56cf37baa3c9969050ed8987ec2a967da01d30d668638676d3688de26f2d3d5ba41ed2f21c8a064875ce2fb15642f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc29bd59b1a5cf88126b65a8cc6ac7be5575dbc1282dd3c6c9b3f215c7cad3a30706b992851cb059f7a35fcb8c5869d57c7d50186ccdcb7c7bbc5e1b07861920ca51e18b9683cd356797f1c0ad4f632ac6dcce00e61865c1f60c61b6f87eb31e10e7ccce01c33e79a337917997475722390f7daedc0a987423d9f1badd96ab68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b4f63513798a5ec715f4a00ad4f148f9c5315ee9bb4b288ab0d5a4fac0322e4d17d924dcf20d26d596fdea417c1804854f39d2a3b1a8fca0cb2aea873e2a6d064f409eeb698c8c88d427c8ef08f4ca6649e8ffcb0569834072bd9aca5b281f4fa5c2e9adb622315fb8c050cab5fc24200840218746a00265a60a9002f69f339;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58d48d0074c3b5e2cfa77538e9e4c58ff51f299ded21556dec67483ca6908c7f2873dd34198389b2f68308b00efc80cb7076e4d4a8e68d95b4e608b50a85228b255260548126183569e680d25655783bc109d5d6a8b9f09b15d62d13049f2fd1b38ab012ae727238089e7c823a40b7fb00531aec4b6d3e9c4719efe58375f65f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1806003dbd71b1a57cf816ce6f5b5ccd98a76f34c748d2eb99c45642783d8afc63f24e323aefe2b6dac4146fcdeeea79bae56100636b314c6abed18104b5363557649260b6b7af3d32f772e35cd7b8910397c3bc3ac7293fd95a6df27d75f831899ccdd720447246d36dd4239888752cfd8f09e2295de68a697497d882ea090;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3d4db20ab331403a57c7680a5a4b2476541ef2666399e995f7c74631f29b68e8112c3108c710853609002c385efac8960625cc22f9304724a4200e10953f63f387d1c6181bf1cc00ab13ab882b48a25803b5be8faced06fff5e22a4692c3f28024a1a5bc03ded721a3aa1a2da5281b9f0ee6b7ff7bc06ee558318c03e55e26c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8986cf5d081e58a4e64f507ea22cd7fd25f2d810f141c0d9ebeb854f4c7999dccd35dccd0b7a57cea0681556fa5b963137fe08511e04fd752d6d92e526268f4d82ddef9de64e34fc6f77b2b58d74b6870929c57347f0eef3ca2d75b65af38c22b58037bdba20c4ea16e0e413c051746b8bb7660a6fc85ecf277f0f2eb3f3e20;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2d64840ebf622952a515b45ef3bae37df8d960b0430a9262b6194c20601cceb3a2aa4227e34d59292331d736a2152839992e8fb2cd55eb11e59c13cbb2974df95885ff9146a1162febb2a3f1bcc63df9824494b5b78bd472c3c8c10ed66d8ffc5f892b5324df7a36e0e90a756cd351a13e1787e9e62751357b8d1b382cd5606;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc39893714c130af0b9db9ba395513b784f80e5df461cd94ae804ae81682ac1164d91c00c5fe71008a0b810eba083a9a7ed10aa89818643cdda7ba0008f5d430f5f0c808f6a4e8eef36cd58f34a6f5d764c7b03b41ef5c51623af3bb96239a453c4afca14957978a87a69c2bb766d6e991ed8f47359e98832c12ce2088e6460fa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1f08b1d0fbe1635e7c2c933a91946a48c52805493a1c0e2a60b78341608254708bb709c268f883985046e6894c387b147c509d4e3a81ad23dc36a2ced615021bcd6a74bef024ab9a01c965a9d60c3a1631e84b563e7185873ce13f072014bc3c68cf3535fab2149248adce2f517b617ef0b4017c7af9bd6d105f1002fc0e28b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7171042a0abeb69c9b585950024db29483250f7c458324fde22a5dd1333c3bd59f0afcb3eeb6b9e002b4662133db0a412ed1539138e760e71d648a999560c8a09762a666c116637f111f7c188c3fb2158fc13e3de7385e67464c30917e137d3e0c0cc9b4213cab0ba457dde903c0d52aa27e267aa3a10cbd1b2e54ec5e08e2a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24391a7549520e2b216ea568253d92da9b0e6f8891d576c9e605a93d09811e52441cc32df4b07f7177c7aa79832579e4ec704a8f2cc629adb771edf66b43aa467aea594e66881838303d7f483c6d1557b805d60c53119a29e549d6738adb1bb4f029d4789482e07de907c14e43f215fa9cb31bae685d631b84a11cae0be0292b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf098abfd9f26b450037939dafaa40d354ce488de5ee3d6e0a12a03c27bad59db703dfee6081d73e441fde42620b65566b9956a2cb9d75aa852cc1e7240cac9a28aadf51a9a3c0b1752a1f42ae01d4c297b549dc0f9f2f82f5451100d6f9374a672c7717986322e5479a46354df60556dd0a3f7c39241e5dbb66e3fc3f2b440f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a4b3858fcba595dc4735bc12872384ccca6694d8e8104e0c05abe8b9579c1e6710b73b9e18361c4e81802d8320dce01510e86c63231f84026272c8e44aa7bce6eab7b594f78754ed4291f7139ecf3fe2d8ff2838563db67f864b8a85e75bdf93c91ea9ef00fdd832e51a8122cb688af3b4fc8a3c9aa62931ead9be7a70605af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda5bfae0cc855f6c319c88380ed98a2d2bfe6533df5f2527ad567f2bb1e92f84d667f3b540c8aaba882856bc5f22b59a1ca69b26f69765b5dd313d472283582c4960690f920497218a719550b1a728c929fd557caa4a4a2b9f827b8b1f25ad4d71cc50222c3d1b341c6bf5b6741038cff4cfd658bee53676dbdb6392dd8acfeb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h770507c3139020cb14df6cc8cefe003c1245fbc80f4d7055323f813c663dcf1c4a61b10b70d192d21cda3866090d4ea4bc59f9cca9a0b70ff661e1501436bc1c1ca811993961431aa1ba9c59f383cb84e4a40142fe958a49b9de03bed5c0f008f365d81e3699381498051f8c0cb9c89f1a86343112227f18248c8af8539fa569;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1c8219ee13e8d736329bd409856acfcb5d0b422048dc9f9a196a765146112c3d44b9c2d073f24b2e42c7071e2cf06c083eb2abb4b47e8af8f8a4b383fd3c6eb11d12f101fab77c91b8dbf2d03712759129c47fe116577a000d61e726f8824367446ae170363a7249c26eeec5508b53f9e8e3fd5b70fbe3272a35e65aa28e48d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4f01be63e64464f32331370d0336a25122d57d566a310b40736a7461bd02615b14f4776543c68e9a6d87d7298fb22f682add133b3cd210ec3742b0db08019de2d95df4b453df53394a5469c95bf21232cce2374efccfb86cff7e3346a2ca8a4a059b3349725b96593fd04cb94ac1ee6acb5c501166879a9083110139cd52edb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6acafc129074de54c542683708052c1efdb4801c8e86e642ca2bd35d302dc698cb84675655ededb5be14323ca6ab921f43286ec9a0fed4b4dbf4c92c979abcb6fdf2fde24732b2a67a18d828408ba573c4c77d9dd92735c4cb61914cd91f47cf844407579fcfa658da95355cd60fd773065f59ff47b0f0ceaeff4f47101a99e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff7a13b9ed6bc58d22b6db75c472a8c63eb884eeaa8e8e434423ab71df19711a8f447114ae9312fa2844f4c91f964a4f72a1a8597199a9816bb4d86ec4aaa74ff5eb168d4db4d800b94c63340ab86e0bc6ee8b5f8d919b116d201cfbe5122434c63d5a7ad2c658e833fd3ff3ca7cae385d922c77a918c80b1d54c792ecd0a7fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc72d323e5587c21b65ccc16e18112ed1141f30dfa1df7bfdb3f76667c250e7bec395fdd69a426a143e1eb0906d785b55a035e0a75cfdf3653557ffebd256cf303338afcf1799cbd6a9dd7f7186a7157d1609701c2704c8e64c4db7f784449ab2d1bdaa7018797e9865c74daf1727e61ca1b3a69a4818775d97467073faa7089e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd51bfe2ae78a0d30e1c79a74eb15ae92cf5c06dbd0da52ecb0f66f31a4f7c31b26c7d314b4d8b1112d08153574c08de194bdaf8971a1bd633f3a8ddddba0a80e9ac0990f3d4ff0bf4c18b8bb26212fe62a9c3fd191c48550a11fd69270592e4f1d9e51dcb768fc2de7887c5f8d954a6983d3937f89cabea6a3dafb126387efc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57bbf950d4a2bc6088b7f0d859fe20cecd499e8e58509a4e3bbb44d99e4dc220c97cdee1d25d1e180854caf708cf1fb0598535039e7898d1914d53c4714832e09bb46b84d9f0f50af93c78500184383bff2bf6dda7895bbbfba3c8fe981ad55eb49458c35903ec6367c0ea8d34e98cf3af6fa477ab24c34496277f1fee06cc13;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfb78164ee3a30074e0a09016db5064b53c8d02d826ddb41a9f833077733207d13fb6b0a4ad2baae43b65073628705a9d32b78250678a0daf953fb056fb8764ec74b5a86233d94ef3a7a51d5861c1c59f1ae3d42970e9960eed1f4cf62ae801760ef1dc7949b4fff347dd9bcaf70dc22499f4ab652d0abb69cfd69e1dcebab12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a915f00a2a0ec4f71549fcd3585a91365600ae26251137ccf056dc487e771ca0a8950036b122d3fd48ae83a80ece44f56f7a60587b5a969c1eeaf3a07ad4d4e1fafeb6d8685d672c5898c32d755acb7f40ff9643c0afc42b7d066de4dce9f0549c647d6743b04f08a3a6abf98fa20e50bb8246a447588f09a82c5a92f496472;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd82e795d1b1b4b2d543c9e1b57e1c08d035a6997f279bffeb3b163c434ba05b95629ebce7798acc009739dfb1a5a606523aa11a960706f2965d0d7441efd8f34e25bb44d321863414bc23db2c4af48dc9f1492adfa1684f9743ae0ec335bb77cdb72c8f78aed836d41c6643a00eee8dd73cc963fd604f3a027ae449d3f11c08;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4aa136e3d49f27ee562fce585d4bc7f24a99774cd166fa55fdf0a602e5394613eb6b47e6d35a6e900bc323508b6777e53ff9206975c61f3ce8ff21a43d50a8b0fdb9c5a46fd627bd807bb9efc44f856a7d260bbffb291175bfddbbe2caf56d31725e103d29b3aa7eb7fff34fe88f82b8b183fd7d1cd928524b6e4ed7485a3fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab676796f0f9f435571a3129997b551b3cb20d7c230da96c99dc6950ef687cf7b6423ca1ea45de988aa501a160b4cca586267e8eedf29b262c5e4eff27ce9383ae0b8f82778e6e4484105b781fbc7f38e4598cb207379af9c7e4b975c65e45913e68489292f823eab6bd5d03bfd6541a074cd159ab997da72b8e76eba73365ef;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a85b5d2734cd1fb39a250d38b34e5e29220de086634c5576fd0919ae41e63d3964a817fe89f6db4c866d364249094fd3b6a3074b54da3ef80b58298b27ac38c706150655d553489bfe59eb0c2596f37b44e8ad19a41473119464f61dea8373d3ea18475ec0e61f7e29638af38ea24ba9f5784a84c50193271829e33b0e71121;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4352ef88f504209a7b08165dadfc6af9131a8f890b1afd9f53e95a53e45d6d73694561274c00bf41b00079e4a860a6ccac60354d1656a5c1c9e6df4997b19be75442892fae9cf3eed40f2932a3e5d868232f9dbe1ed8621837dce59b04a5cfeb20e2da22f3afb2d20fe920847efbf7c322a823c9e4062bad8db19e3d2c1fa0a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37d5c0a55e4b64c88e0945a6764019d7624f69e888f1d8c831c1c4931a3a84268c022873de87db0ddd0e938eeeb35de6bf28c6f53b609178ece496e7ce024ac8a520a0ca63d4d2b57eb6761a394e997a54537dfef197eca8c54e60c19e5e051a8e503620fde9066ab0f2c74c7b0860aed87abbf7e13ea467d74c4af6ef65979e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6241da17640e8cda857c9a33d999eb28c09358801eaf24231f83036b60f373b6eb8014d6cf3164a56e82aaa7736fb1d37ca96f2ae743c774e1ffe900e670f831025840e91302fe1d481a77493617240d2b5d9505045d6cf2a0e587721b77421b0bc99aef2770baa44446658ec44f3b83f5d7556d4a6c6b404d53fe10e30ebc2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c05900517bbab0a19a72d43aef8d60215a922ec29b90aad7e2ed6a6767343843d1639293b8e245c52205b76a51d7380b6ad3e9ecf30a4ca5b6483a71223c06a0eb3b56107294b14449f44ee56de502455ff641ffa54087afd721c06dad4473fa538655028e80e6e82c05e74564e452f93615b7b8f6b427f4f4301c021eb083b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf20c312e6037e2fa14c86883514233a0341cc9029ac29ccee949a7ac90ab743a8576155ea63b0c15f6b645949b1bcaef03462105e0c3656336e3df74684ada5016ac62b1d402b1cae1ed7c9b8e43fda73d56ee7e898789a9f78a57bbbcb7eea58273bc0eb27ca313cf9640a3fc3f24b601c88a63214bdc56012c4e8c8b43e972;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6d6ccd0cff4f1ab0adfaeb855839b04f60119d80a248f9ff770ed8b05fa52a219342fe403fda382c19cdb7b9efd740aa9804ea53387f02de9a1bf0ac03ea7167791694fdddc43c8dbe34d20894fc2889678590b07b7cafd9f67b1c4579c8e1901ff28973502eb36964d83cbe46d9687fa28136e83c3daac38181aa09a06c883;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55c4cef84ad017b1e3585577cf99affe0834781faebd70f0258dd57209c02f5782ff45165fd4fcaf69a90e189ca7470dfad911b903962378d80accf29c47cffaa0096c9cc1e2e33e4033a70553890b3887aeab6f74e08b826d0194450d8e609bfeabc25892640269beaaa52a694affffcb90a9c2ccc7bbc746bbaf77968a0c38;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3b9594562fb55e67aba149aae9cf09d919f00b35104ec93c7631b13584acb87523063e5ae89844103cddc118b653cbe92c8c9b7000c554b79e6784668e4b2487240c22a5291d05d7274361addf69e9a6f58ab9957ca63e682420dffa1bd9e7531e3d45834ac2dbf481fbf18f4a087b64e7355e921b24541d77272cf2591fc26;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1d15f8aa509974d9428644ccab6592f835ebf4204b0f5f05e8dda6ae00bf853dfe4becdf58a4e6f7c351c2db32f695d6aa7fcac4f90c37d18a4e563fe0ae49d2b3ba8742773a80787e5894b7e1c091ebf5e68841c160f89b666f147f25b0d65dea78c391b70e6fe9a29f385ccdb18c41821aff7b31632cb3c311ad58a560e2f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f9c91b83471588816d9a2fd1ba2320bd7971febbb635b18736c4a03a003a86110a52f9724059267ba7835c27d54de338c3ed6c6097c16f08b8ed47251f5dce8f46453a903af027cac7a02e0fa9b3900a8782d2a8b839ebdbeb802309a04d439d3c5c84a52374169262cdc3f2c6d4219b4b21268dfdd76c1a1b5e149f839b216;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38b97a6d090dcebbe9dc7f333abdd794d32bed6d8a51361dd934505ba3ad7c11d8e15902c77af396f3b77be69b75412caf4a2aa366d620ab80fbe5c8d06acb338f01428c1814b47cb2858ca5d3068d1279ac88f511d4a7202ebb49d0e4b7da159b9b1fb02f4bc8bbf177035799efab497c1854399d8a8271554adbcd835aa14c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haee9ea0e2857526ac0ae7ac26b33fe674ee5d13ef99daefc7490aab687da956a0144c2847ae4b088730e8dbd9cabff112bd71dbee639a58a78a310f6e7f6b38ec3763546e8bed5a181fb1f2e4ac1faa6a19bc4ebafec6ece2a2f0add6802eb0982a94498119921331e53b3d289621620416fee2c21d0f82caba2ff62a583e29b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6273dbd37bdd19b7953c5d7ca59687e748a71789dd269d17d379ddf89587696de08b58712d5c8ff32a1fe3bec7438b8bc33095200dcc4fd2651e2d0150e1bb7b69a222f7bdcef15db52a730c17f5f41c483c6eead106bceac852f1e692a8d62596e0ccb3a3cb6ddf372cfab4d6b9f12ff5226dcd0ee3d8507bd3724d2a87b46;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed64ea49eb112d3af99e0b43ba5b8894b19fb978e0bc9fee59075fec46b10a73dadcbfcf68420192507f92ac2ea3802726cac9bd0da5760a2fad62505d656fc92b2c0b6fdac7e8c46288c5e56dc1f461fe0aeb1b105295ac047e904ef2457f1119f2a859beb3423a0eadfb5fce2d958a4d5d77b1417587a88097a00a0fd8d76;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8792df1d99d1805fd742fc91eb8174642449281c81b7b68fce144b72a5126a37f5050bae1068ede0d0dcfa422b5bc3a61f534f55fdb8916ea2dd71428eacef24d800e42b1728f05a46df78505ec3b0d48cb204fbef052c4bace294e99a70c8769edda41a778633d73850b15e278f81cbdd6b8dbb57d3d355085e27dea861b636;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2043d4936618944d2fe670627a2699f0b36f2652ea9e8030824d4afebc54227054a9ecf8e003796f0c3c33290bf7e33933a76222b0deedacf9ea8eb796c7fa8d39692368e211d2474a6dea20358ac3b9681ed927323ba8ad7618ef983250f6c31f658ed509b210c58704027fec58e4bc30d674e920f9bac707bc530868c758db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba65196cb3cff9d21e5c106346a37f64e45fa1687219aa8bdd2075fd3ed72d89c0dfd5bab7212df2ba2c94cf787d018f9b46e632065b6271b271e79dbcc99ee3ab030c1863c08ef715e3c9d0deb0b26797a6ea54a34d57b28f0ce6376ecd40e5d26bedeeec30a9c71dc59743bf00868c3ef59d49a37fcfe9768772cc36e03c9e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d438a08cd960571c995d745dd5b245b0a173003c7266925230fb0a1a630324947613a5c3c7503d834d7162ff3247e9baed014c1e9bb5e1bcdce3496a9b6f11fc9367dc71b64c4d59aff5e6f034ec41328def088d9ca928637e4498e77e1b5903ad97e08b4b51fe1108135573d2ef0d18d1819234ad1915a3ebaeeea188bb23a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fd0bdd517be38e216d63b44eba5330e80ce6d328efce688e12591ca448a4920d433a8d10ad3d91cc9008babf205b26bbb519f06022456a967e58e4b625dd6420bd2f73b46fda6ff646573c377f890f7976a630dcbb37ce40acce6e8dabbf9830ad237535c0141c2930f98933ae3e17a084a95244e72fdf6c056bbfd2b52eae3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8337bbaf85aef2f12117ee5f25074d8f0c320f8e28ed7899dae73be4671af05ec2a337e4e9acae0a5b844483ea485e1962419277a3ae8a3fe1b536482d9f89e805e3c568e11b46782b68bfd03c2478cbb0f6f0f3c0f8e475ed84881929593f1d4c1fcbf72939e160ab36fb1102d7655021d9c65162f318d3f3d61368908408ce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5330f2928861e61b06af3c45670cd902d9ba656f875e94d2c801f6219abab65fc8e4a8d9fc96a2552e2bb86626c5338d7c38ac5fcf2b331a43fd85502ca610be63a645dd558b152ab53fa740f332805a5d1fb5a74cef417e99f61ba81d8f357fef141d91b30c963fb790d3911d3ed77708cabecbd44112d4783de62c801ed94;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30a97049aa0402474c14009697f2a2b68f7581a72f319595fe1a96cecb1c3916e11d336532d5472688ab6e3d513f7fabc23d8b03b73b67353d645f66d2d4cc3d27cd30a3742c36014bb3e735584ea71b5cf0c88e23b84eb103faa7fa851c6b7d6672c18fcae5938c858f28e7880596637f8c6dc7c20c97896c3925e123dd6011;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd686ba846f6483439d93c60696b03a8e9b945b248ebc61156331eab5b53522fa3d246220f5b499fc338494ef779c686225cd4ce61b42890f9ed921fc9bfa68a00bcced171d4f3362b48da1947ed47fef57da8114572af2817d508f0881492d5cdf545601ab8f46d00d452793496198e76d0ef7504444724c8c3c6bb645502ff6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha97d8bea00943ffca48e7cd57baf1fd0341015508026e6d1aa42d5c81b4e8976d33c7d802968e9d53ec752c05058c424bed030de8e36251151de22afc81e0455a54a3c800945d6380eb465a518cf7a28882d4358d9f24abdb7f9aa17d0a7e6db23de080b34de7d33393be1bd3f5e5a469f2a4ff2d192ad747d4dac26d211c21b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he22653b4fb16dfae092aaafff9dd1bdaa661fd9285eddc5f3606ace0de070c2a3491cc083b1f0bd52db1d7728a2060e9e122150a8f08817b7d20075b037bc744123396cbd6fe9677a0c37982623ea6a1942844a9f7393ef454b8df98b17052117f3657830902d7d466841f7000f7296a29dd5a42628581840f94d3a2df5761a9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c4ff0d4a73384178c33df41f133652c2dd4cf07ecc43760bfc00bc9a035c8f6880c8fcfa3de3fadf9634b1ed91a1088a8b516ebcda17d3205ce751fefa2bc2fab7aadc04ebfa34105c345c403f1d3fd109e4067c57f7d67144f04a2feba0ce9283ec5635656c616a4e2122f77e0d39f5ac35bd8e8f68bec65465cdfec666f41;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4316b45d0d63ce766c71dd72b19f737bf31be7be2a1b383004bf3ff9f80e78ce14324fcee40cf5c282f44d743d4de682df64ee1711d13dcafce10a69d018e7d83bd037738192bc15323c6d1c95befcb26b855afd3c696975a7d59ee7df7defe33e94317e96ca26a4ca7a3b7507123065ab98db982d55b929006397ec6f1b2dee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fa3068fd0a9a6fd95f80dede67d9d12df41909430c7c18fb56f0aefb0947a0c73e689bd769739a638a9aaef1546b183cbfc6c205da9dc36d96b2003604f6128ec2032fcb67baa96311fb7ade61569ffaaa8eb47da9cc68ca3ee810ffc49f26800552797cb07e444b7b549186989f59cfffb9d1eb6fa7865ac211c4449ba50dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf98e07910dfd5af97ebc3b99ed919d1faefdeebefd21a277b74f1bb2493e0d9147570c36a1ec92943b8fe4ec9ea34346720710c3b797a73956ab126b29ec93ca03080d5d2f168132007b1229ca4f50be43b6b99ba514fb2abfa11d7c6e01fc3859530a9738a0f59214e90413d7d119963df8dd4022a0da16db9c4af0e0f4d5f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he19716cd849145297f13f9e6f16cdb4ae5c3439ab3f83abc31054b0c6c636a8c399663edc7b97bdb178769eb0dcfd9cc963c88de0c8c358e0225b2012bde6c9abb7ceb9d2d9c9be994ef1d00a028f7de4cb18b3e2b139e9fa0b56582ae9c97cd6d91f9ef924c36422f015a961cc49626c79e66d035a2df5a16e9e9573ed3a69b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ff895d3557a2d72cb4df99688e3f54f487e85f84e5b1a0add9c26a9fe244740e90cfcd2a4cc9931d307fd007b98e7d758adb1532f6f7f4cb722f2d95921f7ca5943a22705a4c4e7a3a312c6b69008b81aea9d22843c1a76b24c5afc9f496bd8d914ee7c534d2f10bf1c11522314ccdb6f1cda7365fa639b26cf5906b1300c71;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c742a6ba311e36410e9b77608a99919a86f2a61c8eaebb387226fdb21e17d3134a4cc2a885decc169264d31bc0941c49406067d666f05a6f3b1c828db3097f10f709c4e6fe23f7ae89ece436ef44f7fb40633f83ea7297f22712e75e38916d2ad84c18249f1500bf9affba398735d71751eba2659459e59e8dbc981fc336684;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffcdaf8c7057ae65f163a15eacbf74c921af44323562881a63705db6458de893052f1087a6b95f282dd51033ec82d4c7cff329bf215c227238d121b2174e50dcc5f7ee1003c39e00933e009060641d8d9f005470b3b7d50e793449cb715f4bd4a6f88082a482bbe065d9f62f84d6a237ea85d74f0a06edb5d5ab9a806c71520d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8925e40f6e6e6e65ab57fc6c3f26bfb35890f685579ab6335deb113b58ac7c3decc3f9d29f2f17065023faf2699543917db402fb9b7afe7dfd82474f63c916275f1944d6c0495f4942f283657cde06ba5ec91c7cc959fa8cf30d9dcfc01f5e7738bad8e71618e93e619463af7fef351b5d0089c0dedccfde6303974f940fc828;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb415569faa5cc13576637a5cdfde363e93aca9923e927bccb6b274fea79006d9df2d8b70e59cc8a4548a86bca324d669d30daf5ce5cd7d852f49fe84b360a6cc33d8a0a4929bacef89334d120bc8eb03f6e8c0dc1e17443ba4fa91b7ffe73b3c20cd888f48832ab777763387ce384c83b922da9fc6c68700fb857361e7e754aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h675580aa067f44d2403eda93a96a5bec0eec13a57b584e69888f39e641e6d9583e93f1a815d9ad0f6b3b51010c87aca5fda43e7abce3b1e0834234e0fd130077e8b9df25bf28f0fd076891e2d6ae772edb4e1992b01caf85ca2c20ef7eed7780b260c2d669d3e4548753f594257abafc8af27d362357748c45c99a556ae0f17b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h815a8831eeb55e615ea79d85f034a4a205bce926d08dcd1166420cc85d8ed4a39accf773fc080db7862a09f8d4e523d8d29c392af67ed84c38fdbf952c3e95150b071a35a36096249405df5996521d4ce398fe93394ac69ebe0b080a23f470e16e21bccd40b7f4ad26fd082e09a692ad7adee4d11e31ae29e3d50bb693bd65a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42a0dc7d599b402f1c50bb7de6231f9a9fdcfce6de45b0c3ee8109ea2a6aa249c9eccfadf58903e8877a142186338d4577fe15c6da9826cd06292d89bbe37c8762e35467c3d6c86dc61f325ad29e4832c24a7f154c8c5b96f893f9c564bf992017e926e1fc7d9e94aa6b54c699d061150083b1fb4deee556eeaeaa45285706fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4eebc09260e2ba8efcea3a77ccfe7d6d88733ce09058bcd29b666a300c320887ef1e9e87d285cf80232c51c9ce66084fb7e099cff92c5bfd86754405e4fd2ef42a7f5ad971542735e7c81a6bde6f54b86bb252438b922fede25e5c91795f303014bee979e4037f7102ba5677f4a40037cb1f9db2b8246106573deb1bb41f7698;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dbf1305ade69941677543a4c15aff57d0174697054c5eb369e739dc7c56b7b9ed8a9752d807188cfa3f4fe1a8cc25beef59712680b79f451f4ee641d7e88bd7d8bea45fdc2bb54fa048a4b957c9264efe417ff4b09cceeaca19e31718c5b05852d5cd9b512f4d8a1e898edb74c91fa22f5049dfc6563ab2c57f33f7e28750ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h179729ed98a04fe16cfb3924f4b43caae03fe1af7580aab40144ef29d9fba6f56ef306cffecb6f38d8909dbd216b5e9ddf49eb65d43d1feb680271fe656f60f6f14096a923453e40e8a60da6183e4a73e351a095e6e2700d25c90f13d4dc659f404bbc7ee5b0aadad1de4341b2d615b8152592c13f4c21638d413f8ffd3ab6dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8f8216dbf5bbf0f8603ae45561588735d97cd549a83567aafb5e06a5aa0187c30d52306a980e7d54e6aaaec5f312d616f5ead1f0d99bc1b7da456f2500f123a18e6840844a39e3992ca9ed09671fe8ef15bc3597f64772bb7889664261766d332ec364b5a42bfa061643d266a0ac41b1185e3788d730afd5dcbd9a08a59d5dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b2510f538b12276394878d48b9a352db46ba298e2cf00def7dc1acd61a25f6320179bd4a0e2620dbf7f79fc04eb48e3dda90dce46c1111af89e3ca319c72f3d1bd2487c4dd8a0396e1f82214568b4aa4ed2fbdf4c1be2828a046dc1a3addd9f8c5d8b1cf9132d41fdd4e5a3d5092c1bc7c1ed99c096afcace6d0ed22227194;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e71ec33f50e00570d886d5ec46a87d2e140facd0342c15dff643fc04b69727704a4966c64c9dd7d650f9a64522571666acb881b1d88e4af41e16eb5ce86c1cb1d638bdc1a9ef710c21250875325b1df9bb129c517066a8029879d604ff4cf2c6980529789eee088461d7d74c46cbe1881a809b2fee86420c92bbc677d926b68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23fd3c50beb20ca290c20e19023758067ede95990478cfc36c04468bb769194bb9ae986f00f5f18f33655bca2dc561dfba465c781d901be67cf027589dd6f4b89d84e58dcde78488a0cf9a797f03215e993f740e832a6f9ada38dc72a2a48e4e38e22f8de1b8a260f65f2d6796f7b8816abe11710ca84ed8f7a877eaa64feac0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc294ea607abc695846b10b738cf49db05af326acd6badad4e80da70861876ba0ab2df302c5ad35690a36246de35b2707cdba6f813d3f03bd721aace2d81238115294fbfacc8dd72d358659acc28bc1b041e173ef01017188f25443fb61e07e57ae3e459a8086e4d2f14c634a312537e3310bf424d6981f25b127bd5b0869b8fa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66611bf54347e1dd97a543b42e25f672920c9544617b4ccf56509f99615391f2a4ac316f8121c33429c1d9676ece7e4df8fb91a66b806f13dcfc67fcf304293c691c731c2cb9eaa490442610ca9a1f691ed46dd7d27ad5d73e65922a0a71b2dc501625f865fd9a7fa587b16ed3be1cfd2e5fac41526d40dd6c9f192df6574819;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ac8813af717bd439d432ec71a416c1875461f6bff10897e9d6637a64a744adbd456ab02d74a42d4421d624893ace5b706568daecc20006fbfd236186d38c05c44638a56169e7ff748aa933ccbc145f1237a0f33649f11c938a0527f7774a57c3c268a6e97fa0fe6cf7e1b21221310c9d6380a70baecffda9d31d778c221a748;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e2a9f44c8299c96f1907aa5cd8dcba4d13fadaa13ded2921c8a8c958f2e5fb9765496b65ec9d5fbb0532805c1ca8813db23235471454ee01c6801621b3ae546b8b08dc1b05d41afc5bd17e822223518789211e6f9ba9ada898da1fce24592067f48710e4af5d76d19c45cf65bac05725d0fb9da935bbbd415c18f16116e08b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb23fb1754b9dbdc88b807ac32eeba63146553f65bb6f80f263910cd599d87a6464957f9007356efec62000d42e5e73075be74848a75ec299add49202addd165629ed197a12d291c8c942608d5adf9110aeb5631a1d65e378f37467fcb2a2295576576886c2e55ce4acb07ac1a53f9ae9c7cd379ba7447bf3c6a71d4e050fc95c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b18747aed28ddd03d7ccae91b7feec0113d9a4ab30f47da40ff4cd9fce6efdc89f1ffad86306d97d52d3607964db5772f5be102546cf1b5dbd342087f92af5d8082f137980c92a0be3507d331204a8295930bf545cd0bd63877559fafc439bf5e38db762d3b9a28c80d0b9efac5f3512e0dd57c33058901f23a2aebb8811e74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h820b0484a42771c7f74b80657d68b9f8b3f5124626b4ad55f4015510473412ad366cdfadcbbec03cd49288806d58d76abf1077b3be9e5294a28ff5ba8c31a082f193d66365d4265b7b35268c9a76c0e8253a9491db724484b1c5c6471bc9cf6b4ed1ed3423a987a0cc70916b6030c1592c42f78ff0f49c74283fbad6325faea9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49c13206c2dda0ede76a2a5fbe12956ecc8b2f4c905e8513a70f9afcf8da82a3469226365e43d81b2c904173143ae7ac0fb6e57c514c1877e7b3f8036736b420032f944f494c5d6676433fc33c31940c4b231fad6411a38068b6e8e3e37d6dfe420e1777de4deba1dbd2f6569d2b1e84d44f84696b7181969482417f162aba07;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e7677d1ef86e717e7452135909ea2be08ab3049503778b0fdac7c2e745c391e1f0c63219d1635f4ca98de4380194232a86bbf41daab6fe433a5f1ee40a3d4206104d1a086fe3616aacf8facc0e2df1d9e45250467e0e948a1b0145251dd3a2d2d42fe79a7c49b8bc42316333f6b7a9e914eaa19e59426aeec57dd082e3d8c41;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb10020b7b6d78c9570d280c8abcdfa5b3f8d37607fc810590ac6576b8930712c11e8907007598eac3cb2fcf229dacfb044ed4504da2673a83d5c7c078d84378c69e6ad4cb8a2957d1479c91690c2c111f24c22ab62f308797921f24e1576132b74861173538a2266923bcf2ad679d148c2825fb0bc7c9ffdf6ad310567f97564;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he649f4f9220467e9ac9868ccec6170f15a17eb34ddb60419d077f3c9b38e8c150e3d65c347f16b979b64d5d45e26601882cc3d5128271e089070d32e557e8ac5e9256e8b199606d49a289f626c2240c81997b94d841c2acdf222276dfe7bc4a3afb873656f58bb6eb630a1fcbe6367dbaf6dc47f462367e4f96458031aab88e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45ba13b6dcc5a8026bcf31937032ae3121e8907ab358d043802260aa34c1c0aeb0cc397e08c8d87762831a905137d0c26658e66fafe648ccd815f01915b0a8b1e1cab86602f06aa16e2a378da091d27746efc552cec739882b7909cd95002c2ec61b11522a8cb0c351c264a7cef27bf418a04462210480bacae21fdd46a5eda7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53ca1bc978fa0d39cbaadb8d4abd1824b6589aaf684f200e14430691467fd7a2403b965a8589b830ed18558da53c7bb61de231e634f84c764a743f7a8967be915e9bb0cc8db732e05b326db91c99b4349a6240419dc894548b3bb71ffa51493c921384d35c74189e74ce45743041a2bd8dfea69d90cff6374446da514eb6a4c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdde2b38f7c2d9850c153f158bb8c74914b9e05133d81a3e1003b4d4598f8cfd3beea75734e09650550a29c145ad5c09dfa4c8096db135a7f0a408ea09828679d1bdafffb4c20a82af9c44f6f0012cc23cc8dc1dc4c43960e8e3c566eb939217cffb004578670b5e76c6db778526860e82acea3de0757529adeade19ca3e36b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h980fd9bdc4b93db126c27c9bd20048c49a687ed74e40494704a6902393b14d8803e06ae2b26ee08de27eac5f5c891edfd11b3027e8a2b0d5b11ee20f55fc90030ec8d50f2ff6a16fe3513a8597a4c47fa3710ca5319eaf1f96bfc4113b0b10e99eae1272cfa8e00994652693c5066d67b87d7261c0b52e1e62b823a5c0f11819;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dcf863b0da29f8486e72062edde886feea515025a95ca040a4ba67d3379be65c82a37e0774944f8144c2e7f508af0a46f94679b4fa3d3173fa31176b2fc96c737614f1ee2d669d29705fe80b334dead3f7ca7533dca818e8e295173d4f347da282b2d2a5dd33998fc0dba24ff1bebcbac147cc44e17dba9500a557358377793;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h154a5baed7f5c8e85037dc968b5644b3bd0285e98ad299f8ee1a0b1fb277fcf85496c930429a43ef1182b8ce739183c0f88f6546e877999dd4bf814e2bae785f1b88cc79c774de7f0d06cdcff8241c9da50bd74ea9d4901681e8d1a2f7404be26b138164f7022e6d7eea473572f888d7de3bb0ed8d7d2c7416e24e966f527874;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac3e6940423004b5b545b80842eca788bf670f70e252158d68635e5ff1f94616ad190cdf037238eb93de016effe0e492b8496532d55b0f93ef56e632e005590e844480e9c9d66c54f07fe56c3c7edeaff568252f59e8e3a7d918795ff68a3587923282954e5ebc45ea811cb38cf29a18bf0ad0c7d0a1f7280f5d65d5b6c9434f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c46b2a7aee2337991d377b8a5f5d1fed4722e02b52e254d0da24a58c3c5cfbc0bb3b8ba806504e0e653cc314af5990972821aae039a9234f24b12d475eeb3d4b3b23863e597b7c99cc59ab4e85e0b6dd390ee5d7c00a68cd0161599ba5208d7d6eb8f9276903608db2d291e71d57c1b4083ba14f93f1492ae99b98021036566;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33e8fd2607ed82c5c86bda402ee9d738c862fb5cfbc5e75a7e5f0c9f06217fce762b8030ca8cdca1d302754874b59dc69ccb3081a454b8543e6347792cd10102ae32a7da12c4a644e77ce456aa809459390c9576c2ee3a51db6da6b1095dab39de886c12968a97435f188c276ec539667859394bb922cc8fc4af269ea9aeae79;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h891c29acd70e37ed18df265e7c3bb123dbecdcb76a9f88c7e3d21f383a15d25798c4a6e0be77f374ca8ac75e0e5efaa2efdda8b2a67d05bc2e55786d3393169e68a0cc362ad772ab115d052027d2c041d71fc1d36b720bab99c2d762df2021aeee56d8dbe0a10a6c80dd455e0f49ff399a58c52d329ed5e063b29f6e7b201f75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d2607942ae2b27ba11d1b94bcff04cff0bb07f4ba43f7628aaa7f99233adb0e474f737622dd292bdea1b7414865d7b98db0ef7651f5feef862f7d2b5b46a13ab0463e21839ad08c3642fffa17e6283e10f615346f4dc95c12a458697a845b2665125578298dc90e21b6a2a891a01f3e1d4df05a6b439d5eeb1bcd45011c9925;
        #1
        $finish();
    end
endmodule
