module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bfdeabed10535d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h688d22f8f3609d37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d6093a3561cd62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b66f27ed05bc063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96024cd2a5e414dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h478b24b6c2b0d4b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee3547d4356cfdc3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c15f2996e2075bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d83a72fcd635254;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf3dc8d4114314ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92662701bca733bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4492ab151bf9f8b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ea7ac30d27afba0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c41796d3ae8dd37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h969f3b2bafa67c47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbf21c5a44820725;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66233081f0b71f3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68639be47e203159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1382c34bb568a7eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde30787fd188c36a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa87136dfd361b5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfa2e66fdfa3c3c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3636a146f05becb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b6419982f0a1135;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadee40c3fd455fa5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7481281469bbc67a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c016ac06439a59b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b0cb9c3e165651f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd40e73f6a3836fbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h966dafdfba40421;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha844a8a5afa9ba9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42cef7dd9a1e2fa5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21ac1db50d6483cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fcaafea225c0dad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70406532f3184a5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd37bba35f187499;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1511cc92d93434d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h114a9491c66f01ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed00c225a1735cd2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73808fc8c5d890c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ab6b38b0e053db4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bf0b3a0ff4daa7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c586a074c83338b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe93ef9187f48204;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ae22abe49e0f1ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b2eeaf76af39104;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2577a07b0dd278d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32db809fa6bb3a47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9786a45ab44711ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h758c585ec18afba0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h650adae7a0a9c68e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h551ac1f7ccf89e07;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h887ecd5f3977df01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc86d66ff7c50fbec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h513af97a257a95aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4e54c8d8ad106;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba9c1ce3968195ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecfba394ad0ae944;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h551b12fb7ec3620e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f4a064b780c2389;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28bc05498302ba64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7894ba5585234e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc100c6f7c7043255;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacb6a139f311e096;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1a11136d44bf912;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5671b6755c46a7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h976b25f5501a9e91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fca899cebfbb3f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0407eb17ae48987;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he05a9b8ce9e36551;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc99b7e87f1bf46d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6bbd60796973aba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8084584a86f3c796;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56eb425db3aabaad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3921a0c957d707da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cf7645bcc3d39fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3351562b194570f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf29718c96dd871d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbc07fa418890c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36eb053ef280f954;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d625fc70433e699;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fa4d137fbd61ab9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf7301202a98fd7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec14dce3617e14d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4628ac673f1fa4af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0dcb9c58d04e88e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58d7ab0ba5ac38e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2e2398e1a917e8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66b7779fd2009e28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb53743f7a8b97cbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a7ffd484f6998f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb54ef5e9991782d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58deaff3f7685298;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f26bd60d337778d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8ff7b1056a24d37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fe0823bc36334f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60cbaf0424e072e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e9bf324baacfb52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57bc0891a9bd0237;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8fed433ae25388da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedd74c53be2c337;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd7cfea78bd7489d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h932288cfeecbb16d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4a77b7d8bb2170;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c7b299890542;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9756f655310b37c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fa70fd84fe435bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf1d0ee39ecd7bd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c2f24c865b19072;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca4dfbad839e64eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha71b9b2ff26cafe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea0665d408333603;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ac226e758105e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb5d391ea84e7960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9cbb005ae5c1f12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a65eba974f7c0b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f3dda4259c4644e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae79f40dee86a98e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8922dbf994c132cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cb1f8212ed31e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38542fd2cf15ca85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c81efef83088214;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc184543751b376dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha573c2979f8bef64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6879d187a839bcf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1341ea48d5d7a148;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ba94549fcbea19b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91fe679aa380fc7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36c61f3531183b5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6af6db9d62751aee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd11bdd205c43fd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e9c52bbf4a5b936;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4367c78d18106d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50c48a38ffdc0c12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5e9fea95c870d9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ca084e006ce68dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba17643f5cf16ca3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9817444fef8ddfad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd5c9bd60c410505;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee966f3217e87313;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ba7253f9ce49d8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d95e7a02d6d713c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d4e7659c1b42225;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc01203087872fb0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c39013141621b3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc200e94af8edb06d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2e6822503f8d378;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f7fd7f65b5884d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38c2e0ffe059a490;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a23b0f1345cfed2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad976cb48e88872;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98739ccde62f2f6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb782fb68a721e22f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2e4f02ce01e3aea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h313d1ce8b8481540;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33635eeb68e943d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d0df8ece3ceacb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5da9ab765633c3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he98d067082d162de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc164c2c3d9cf8649;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb509b0a13a0c718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2acc5173ec41d5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7be2f159abc5823;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1de8d16ba5a86aaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h484f86494d4eefe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7a64866470976d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d43928e659c0c47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc364bc6813828cdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0a5d4b5d79c85a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50c66706e04ebe6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc005b1ed137ccc40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2307ff034f96ae06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c1caa9acf9f1e14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44200c43d14ac9d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2117ca9b8f46641a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c1e898e5ca593cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd20c12741be9b512;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bced64cbc41ce1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6cd16e2dd81dda4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cdeec20dcdf3194;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h659af1bb405b2b14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bd153b4968d940c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52d69fbdf6e1651;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36540e3b6c56c3bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4efa8a96bb48ca63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57997d48b109fec4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde107c1c6debc5b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h763eb6fa806dcef0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h816318f67c76006f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b2a549440724929;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c77bd75e610ac74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f680bd8a8473f09;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba7b4dbe727f54d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4bbf82e3698fb2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf8c58672145f1db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h865bc1cd27f384f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he289d2ddd973f8bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7ff9efe46ebbfcf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf463a6b1d26af6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8065b0facd19254f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9419cbea27e55366;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c59855578f241ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c862c4621f68718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda4c69c1f3770f97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8326cce5dd9092cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9e0e82ead4ce25d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62958d4f4be9d3a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a1544ed91b4969d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec34ef2bc396b538;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9da68de4fa1c8903;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fe086c46a409a1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e5e148be064049e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2da780ed11f8965;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h879b4f5416858729;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9bad4f31a751800;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h527c8ab42b5d188d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff5fadad18a8b5b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a70414067b5f2d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9edf839a087ecc41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e660bee0b90c894;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90bf241935c9253f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdae0f6cc8b30a6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h619c87e5c149337f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c37cc63e121027e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81474953e73acb96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2125adf1d1151c39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8171006388067e8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7bd33431e1535c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea911a84c948dc41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he68d12a4b92f8bd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7ca1b4f1cc3f69d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc88fb0863a00f643;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81d919351e8eba33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc22d139086e17631;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha75fd01755ae82a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha961dc54b4d94b3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f2418b6c2f39b70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6960fb5b75a9ebb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2770c8ffb706d96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ffec71ddfa5cca1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f7d583db51f06f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73c1e7985e40f9c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85a2bc09427415b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha00c635757489fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35a730028be31a32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha31eeab328a9f47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f3d932314bef9c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b5dd5ee66317621;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f7f607b471b98be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c832304b2c75a9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6384dafa4105ede;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b996ebe2069d0a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10fde4ba7cc8daed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaa5755dbb6f9f73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he91ed68f0732f0bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h149308a89b7a77c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f57d1521f631c0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h233a5ee5e75178;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34c93df2a5ba9c54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafac6c45a4ed17e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31dac7cd410d0589;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90c34d89e3ba2349;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc06cf21cd6ac06b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee693ea1085435ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5a562813791f159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3333cf1f493ea72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h112551eea8c57622;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9e204645483f997;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8928ba8c7af854e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb7e4f154dcb55ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1079675fc61a3040;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76c56503ea51263c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18b1c799bc225311;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4adb457a4ffac8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe59126ee5a7d4d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha825627f92ac053f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb530e258e5c3ebd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha44fc9cca726ba63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43bcb1d9ef2973cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf183d13b67feb6f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3e9c351e81c154;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbafed8296aab700;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf195d3c28fa37a28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b3bff015fd1b072;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h366a7779fb1df624;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0e925f56273f174;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44142b7ef6c0afb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf1d60739cc5a62b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40be2ac01701240a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h219da3a698569ffe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dd46e7f157ea234;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9f4000cb764d9b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a53982d4d42909b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc09b40a8a8d3ad4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41b4977ad434a1d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h123d21280a030894;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h720dbe100fc13db1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc87dd2045cdc2a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11a03567789b6614;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe2b3d642b263604;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4afed784442583a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91fb72e5c044d966;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5828eb8dec64f2ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb737a8a368fa3e23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24109373e12d8fc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ca832242071f0ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80edfb5a72b3b1ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11f6ce80df3a623;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h651768c1bc8880f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32595b83d23b49b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0b120af701ea01c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d65a88de6a33213;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2c9a2fabbea890d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h457d94094e4c4e57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d6d3c5fbd3a548d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef946a6f00462d41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h946543fe063ca75c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62e2d00f714e4168;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b083420c2efd980;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28c71d8c1c2a9778;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe56a9fca4261451;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8cbe53db79ad09b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cdbb5dbeb85e410;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9147a0165a4c920a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79c159fedeaf5469;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d9c47486b897e17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c7be9ca346f06cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31fe7b368bc97163;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6e4a0b5c13fdcac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf039b5ac591c8081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbef017ffbd34bfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc8261650e80c4fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cae60d312af1a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52583b68008c4f4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d20d3aff51b2fef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8971ea8775ab1f48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd58c2ebdd1c2bc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e92be7b93174871;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd58a670194283ba4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc953530d52920c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf02a56a2bdeea07a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf77482e81cad0bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed28e98e5c5a13d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha07821f259992fdb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d0391b64d783210;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ec7cfd6cfdea990;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcafbd03af74e8ee0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h643a3ec2932c4444;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fcea2568c1538e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5811de27f60f5119;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5f17face6ed77a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a7c4fd7785351d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3277ec43844fbed4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hade507cf509adeb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2877524ac11ad648;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0c49105758cec4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0809702e1114ea4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd0ef0513278cfac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h183089bd5b80082e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70594dc850dd185f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67e3554493cf3ccd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9058cca23b4de8c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2cbbfd3e56406f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9260b7b72fd7e18b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h102edd468f987498;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7574af0a660cb188;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8805084cfe3657b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49df54e8bdc9ee08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h579f28ef39644804;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5eb0ebd592386437;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebd4d2e42c87281b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5905e73a3f689fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe4763b30fc4074;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h543d6aea2529fdb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2148e41596669388;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90c38444a74d20e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he604e747a4eb4dbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h212b33b8bb5782b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8c5b1a3e4d8a2b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h903d913083520f3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1284e2dc5a7dabf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b6c6afa1f28ce21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe8b9a0d1bdfb5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4031b16220d4a993;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h335d906a0477c925;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4c14f3cddc27da6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h809d280b0989a907;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a6ea4583164bd94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bf741cc80589bc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heba2604b0fad8c10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d68b3a0b5eb0fea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a181c754a079d06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4efb877a9ab57e4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h122730b03e42914d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8981a86de862e54c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha22abea06ff26e76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habc69590613d80ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ee66511629e12a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd20b0d89302512e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67164472022d9e03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a564189d18720f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d269930fd15d7c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heda3695f1283da10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3519b66931811c31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h194a35a64f9a2551;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9460538d0384795;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2e439cb73ab905f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3682a93aafc12dc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c1f2a627e19f02c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d968c7da78a7166;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he963db167a993ca1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h443b579d1f1f4429;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a89a6f4757310c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32790e2108e53066;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h579e48b41750abfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6aa9bf38fb535060;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa33c2077080bc8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c33eef58ab5cee6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76a89760fafe9074;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43ecc5edfd3196cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc93e8a28fb2f5d56;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7fdcdd42ae30172;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67bf98b850e06d14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h966b4066594cbfa5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab9fc4193ba69f64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6ee0dec02b2d84d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2667735d777fdc10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h911e0de21723a9f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h739c33ac3531b261;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73c8d4a4ff8b4665;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha900f56b87540893;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4db9a7ce0fd6720a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heab8aff52bc3497b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2969973eee744972;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38ed40f87779460c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7e253c8bc711224;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30a7ff8f0e0800a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6477c194f7d0e768;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce8410d2999b549a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h351f350c16450665;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha894ce09fda2acb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcc76a5dcfaab585;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h984ba59de45f3f86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46f0991d0fef8fb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f3d587d9b7b2e8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hece3e07e9d56b235;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cbf4f442abfe86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcacef12f8270b534;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2196aec17ab9103f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac790174c985e09c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ad97e586e1f9e9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbafa9930b9498c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha158e07f86a59b51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha41beea4fb1d4e2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h536a80a7096787b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha166ba500588966e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf68f45b4712b847c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h658967b75484f94f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60fd391cc81a22ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceadd41d90769ee4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83a18d52efce7ed3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d59fbdc7ace3b67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd3b3d53dbf8e4de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had5359a1e839eed8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9017beb006024a8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89715f30bd9c4121;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h918ae9d85bd85cf1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc85efef77656ad7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0186450b0555ea4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he78fef0b42282227;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb35edf85f2d95086;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h787c852b59878b19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32a888126613fa76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb069e9db316bb337;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c89361feda0262d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72e865e35417ca1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd3768e85fbe9f67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfa19ed43cbcf80a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fae6c0ecb47ca8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h871b566626d36e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h289268e6311bd16f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1039f2f2ce2960e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82d53390939ded65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b5c2fbc5bb39e94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53b7a8f7ad14fdb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdc83cc996ab1e2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3365eb22ea37a0a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h976efd26917adf41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d7e862285169fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd97934a6cd17ed27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a55a0cd1e0ce28a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8d206b02aa82557;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9329aaeeed5ca5af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h387d19e19e8ab7d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a0e41301f71c5a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5ebfab0ddb6b4bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde0f92b3ff1d6462;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1c0bbdaa647eaad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haeee56c45e21a68f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53e55394c58a86c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5cda3108e4c9aae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fd0695993558a8a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87768136e8456cc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h697ea7a86049878d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93ef4e0ff29dbceb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb45ecbea315ab862;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7b24bd0af48669a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha60a05c1ad3d1465;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd26f08b99b46b179;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f3ab157e4eefd8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddc49043071bc8b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3323b2da2ae1e9ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65326c5fc671b1fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed31c6d2c3f9bb90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69b0cdb1ea11bb81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55bdcf70ff9fd170;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55e1bd24bb924e59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2f96183d659bb13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2903c4d4cbc261f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62b1f53e2bb6db73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h815584cdc5a83675;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda741e223b96fb0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he80cc0614d7ca542;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8bf9200c8e5fa21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a9f6b68c73ed903;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc105d0e75c30d25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe8f8f16d2b4b47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6285043fa831cda7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h860c5dcf61dd07d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h993e781af2d111ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc35ac89680c6e513;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e3d05abf39cd2e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc791d7f12b2f50b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e8ac256e061aba8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfa970ef09f89e77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18a29b37d98a536;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd965245933a33e1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h268b530ffac2f5f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24cd6a9f8563d32e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h509ff4ee7e2a940f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a38c132a47003a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cf79991a18a845d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63d31638f259ac8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b91e482c34f9766;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa94d417323e9d91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h529e48454dfc1fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6aad940953205af0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7cd75b3049d61fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2eaf83ee8d9b5ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc58012814dc5949d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93bd7be4c9890d45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h915a74afe3eae7c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b62320ea4c2caf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1156b445a14d3751;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26a826cea87638ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25ceb87bdcb68886;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72637cf0bb9c7d76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85bee7b2714cabca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e2a545ef0b37d91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf0e55579aca3055;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7deaac45797300c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e32b46f37945cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b7788eebe08843a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha902cd592104feb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had9f8526e978c92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb56374897dcb1a98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69328ee245d86c79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h232aa52978f83a85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc0ca7058969238c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha58b3a60293733a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf7d2cd77d6caf42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5910d9a65f0bb101;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30f237b0ae7d5c5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c5a8a2dad32b326;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8b4a377aa4b710b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he458f5fb39d18747;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee6c7586a732286f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91bd26ae1cc06f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b16c8f6d167e79f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c1eda06caedd4ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b616f613a248549;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1c65a5a1cc2db09;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1a00c2dac7c9537;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfab7ae22211d45d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88b1f6e3b50a9f15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b01ab9908eab580;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf220cf0361b7ea5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8efa6f9ca129a087;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae27e7838bf07dc1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2428c3dec6e26d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha269560e9eb11040;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a8894cb968fb165;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdec810e9be83e1d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18f1341591c56e8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd69406df1674fa0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb22e6035df184b58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd690bb4302d43edf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h881e44ebb2f7e13a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e73db5c24758b6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed36bce6a251658e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1195a74a5b86d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2840558a7246e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb750626c8c11c663;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he04c554b1a9101b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89449bcde0820097;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bd6a38f833725e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c2f695802070078;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26cb69e93f366496;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c7d546dd3c41350;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6eec550c0a29c5ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h303b16a80777e14b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59e1515fc06f47b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd158946c4aad1bfe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dcf17ef19d72352;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha337fccfbba89418;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99b95cc2f2b760dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d1c24a9d7ae6f34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18b11ec916d6feb6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfac964faf90bf2a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4f7b88b45e48a36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c3b79cedbe8508a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h782ab5cca28a1a2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcda66b8ced10c149;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ebbc3e01b8ecd5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h561e165eebeeb257;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf49fc3b40219e181;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a027b1344250667;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbd3542267137233;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47f14b8b57570e9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bd1586e7634d568;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb75e63609c609c23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8309b8abc5a2a9e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he91e6816967db85a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he91a944edb4300e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe44589ba6e52b43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf455a4bf090b3b0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1506b0a16f6a4f0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18d62eb070457008;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h227325b6abbbfa90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ee362b663129cfa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c8d5542b1b325be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc3512594e939ed8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd347336461c8fab2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h997f3baa3b577d05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c705b941e995399;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54e480ee1ea97cfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20fc7584e9295594;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6b0a0290fe8a29c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9c313a52bcfae75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49aba04d03a4739;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb19a1dea10150860;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1845122cd9798260;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf871ab543a03869e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7e6debd5249ed7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5b9dac4a673c275;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd27a78d5732e03d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefb10dcf028cb60c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2dd5c190861d730;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e64bca7b085b574;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heacbfda34090e108;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6aa136f34962f7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc98bfe22324861c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1dce019290b5b324;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf297d0f50a400e20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb12e2f46afe35002;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2a49271ba6b4d44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e5b82d7d2fa4016;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h118d2700eccc45d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96015511ce1ec66c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf0c2a3c9add4499;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5120a061f32e9ba5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ce16a65dfc9d93f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e8ad32e086bd6f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf77d63266147b1ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef1fca57e3614064;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12e8bc85a9f68657;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a815087b3d353d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfba02139a7717f20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83773fc7c6d42241;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25f0b6838f86c7eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a6773d0ca84a198;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfceafeaadb0b803f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62a33fc9c6f1fe95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb855bd51919f65dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd72c645cef349195;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ae64ea8c1ffa32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafca4268d966dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35ffd89a729fff27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h441d74e9da8bd745;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba3cca8daf2ec11b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe2f0a98a90dc677;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he404a41a5b7842ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd35f73241770d320;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4eccb7431c85daf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3b5fcf33d031749;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4587c244a18535d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d211bfbc1902ebb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20198aa3c5fe8098;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5577796ef9b0edff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8b992b5b2712e47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heee797c37ad23084;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h646817d6b3c2a761;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d233162175288cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fa2163760f232c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2767049583ab5397;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf430dec5a2ff9972;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha55284e401cc0a96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2180324b1166cb6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24585255d91d8a02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h917cdc1c6e1e6173;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37c6bedfc165cab5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d741822eb91a1eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha32edf4f590d4536;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9ff578263d8c545;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7cd84feba65c353;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf32da10d02160c29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6571b178742b0e1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h651a6d0ae2d2c37a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71c225043ec1196a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h465f6b89f9be4b12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9392f1ec3a90f8af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2857e4989957ac0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6603ad089b80525c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fdce18613a6d22c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6099c7dcf46563ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98002d29f6056329;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4583935ec1646b3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e1358155dbd0b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h958212f019a159be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe3eb106f465350c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cbd7b74112f9b80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3899c2d0730a55c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb5589a631e073a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd19a2117e1dd04e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b72d9cdf7aff55c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf91af37dd676ffc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8fe7cff82b980c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35e3d9d85d790877;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa20f4a115be1530;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92c71d148207dbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha379a07fb7e186ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10c2205efb93b71b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66ba49075bc264d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78a73370e295e6fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae639da715561a7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33a065ac09294861;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacccae2cd090ec74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbb1b91e179ebadc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h217e1578f33e66b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1739006899ff8653;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37be34f94f0a107d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55f3c2f8652d804d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc87592d2602f2f8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e3bf68cd6e27049;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h435712d60bac58b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1bf3e4bde223846;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9ad2b39ec1cda1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h477ca494a5ad1a30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cbd16ba4cec3512;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeea6d5992bdf655;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h463a92c1d21ea112;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9633b76d3aae760f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bce426a32613ad2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d72e9f2e84d8de9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57e3233ee95e4f82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b2cf2440e9d061;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4f37c7076ef00a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc384ccb8f9392110;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b8ecf6d4b061c2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89b8e9d583d53e54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7701ce4015749584;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb8ddc8a38fd48db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6a233886c4ac01a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9630d406f89c1303;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85fddb57d8b67d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0ec00c7a48ad353;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d0e9e29854c522;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he116186c197a736f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5be52a34e38b7b92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6eb04a4ada25792b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8bee7c460452cb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec1f549cafb12585;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14adfee89ec21d2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2094f6c210df118a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e5b056ed79edfb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b3ec5491d540542;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49fe0a71ae47106f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67f56b424d13ae82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9724efc6b2973db5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h799541c47239ea9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf541808f8ae29b09;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b91fe3a155173fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b3087c0aa8b9cc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bb0ea4d9216f707;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ffaa0be50ffdac0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha46bdd1bd1e9d95e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcc6fbcf827b7ae9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dab390adea2e8df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd62b376e8c18ddb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6db639739e4e4f4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99a15fb24512d68e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fc68c0ef969cccb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9ddcd04110f4aa9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14c6056b014fb8ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7111579a69fc9081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73029ce475bed9b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8260a6976db6069d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he005670d24c178ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1babe5c4200d204d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a7c8faa06efb1e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h525136dbe96fa36f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddd75e41bb5ada0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b08c51864475ce3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe84df66f7a96c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h567446b6b06e7ae7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc15cfee46675411b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94aa5ae1339458d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf95f2ad26fcef61a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55a3e548f057ebc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea3c4e18cf1e86a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h122abacbe92151b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4cad1fe4670e80f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h870fbd2baf986ee5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53c506b991831ff3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ea5136f9e09d662;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h262465ad7430c7b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c489dd34fb3b3e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1555796fc82fd854;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf73d5a93b9e3d790;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h726d37f27997c5b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70660706cb5ce2c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2731e78c5b259c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d181ec2c4bf1253;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dfc4642e2aa0288;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b81dc927943074a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h168578a09938c70c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38649f6039b69e75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc5f13e0ade878ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbaf327f88d3a95ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1270b2317c8bd0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc876043cbe2556a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb29e803fa3032f59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fb75bcf471b5104;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf54ced55cb293489;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f4a961197327f75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a05a362275591c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dbf73bf15da2408;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7fa3aa24c32992b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha064be13bd6b4041;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafc848dcc6a3545d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79fe414830094643;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h557ba2ec9900a08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h872412d406fece9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b7397520c0d087d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7d5f70c5a7c7822;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d3eb1c0cbbe713c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a0a479dc61d770c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bdfef060ad10eef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he510bb4d7f93ac5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4f0455a3bce1d5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f0e4586ddaf15c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h897722dd187cb954;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e891ac1f7711f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecb6ad2aa2bc2db9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56b30c52caec74c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7974cdfa66fd7e5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48ee44d49f7f1d40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h392c36c3e9ddca46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbeb071e65d26c8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he044a752650056b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14a00e9938393d48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf77a806c561fd44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8405a0289900cd10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8297ab5b6efef322;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ee5500d86087008;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f976dd6166883a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc97e928dd1277e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a5bcc9ef8a6067a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6dd12e2adbd6d1f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e31e5c8553508d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h776219ef5bfb9085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6131b0daf7a0d0e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c7a48e85ad719b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3337d1ab0111ec4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48242a78dce3688a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd92b2ac50ecaa70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dc3f90dc3deb0bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb45dca89c7b5e6b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd8943ef483d39f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9f3475a17dc3a13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec7ca59817e40df3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95d9d020b863d240;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d92edfbe92ca475;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a29deca3ea32767;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a20c923bd0196fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9705317c8c757540;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1bdcbfed1307292;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdeeeb9eadd765546;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd1fc7f65080392f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed58e711a7048ab2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb5aad4bd2a054b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bf3c7bda6fa9fc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1bd6b8a4972e7a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab056a850c21d8e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64b2858a9b9dfe43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8697f3a322ffb4d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f7f12838fc1365c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5ac0afa9d0f3e70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a32eafcf3f792b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb77759ba2fece44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha523d952d3ab307b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc360daf6a979ee9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b023b1eba907967;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38924172703c2fe2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7e086eb23810a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7edbb90d164cdf1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb9272f834e647d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf698f39b312376ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb2d23341b7226a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7aab002684d0dcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he915a8b70dd03f98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5674cf2b10642f06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2a27582fc107a66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h569b5a986c49c361;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37c5fc6c39f9e091;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68fdf731cca438fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0b2253276b08bf1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29fb79d8c5d8c32b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90f6d9ebfb7af9a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed6892697858cd6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cf0f679119c829e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19a517d8839bfc84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfced3288a109faa8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9cad43c7a0ed3ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9284c7c49147e3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6660a6cc28ff06c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h633e2c71f85f928c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h715c71651cac92f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97a1ce030f79a2bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb07dd90823d8c603;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3c3f78bde45a915;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64a7d52e6b22f7dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d3d04d123486044;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2456690ce353b9e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dfe49123391c7c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7f77bda3fae36e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71c923065fb0b293;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h215f9e5779daedea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b8f2d9cd98ce07a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc31a231443df77e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d60ac6341a386d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8608cfac11712d3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4159f85e0b78fdc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7909fdd86ab1d726;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h329bf389d8a7a883;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6963109e346eae4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc290704a68c6d989;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22a848cd27d032c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7ca1e7830516dfa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b063a7abd2add7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcbfdbbb5106f1f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0d62b6aab533bdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fde29d3677e5458;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd97068bbcb4f5e87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6052ce3b35a9b1ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h380b9984c005ecb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7621586aabe3dbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73deb5c5134c616c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h834d747d426223f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed9046fc284c328e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c25a01f3226e4ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb59131d5ed2c65ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70d10524e6b668f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a91ee38e0a36cb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b2d3ad88babff8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92c4ca8832f99a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h378cc5e7155c0f3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64409cc28c2a02c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ab68b3fc382d937;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca098e605dd03b40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24dc1a8e5ce2444a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd363bbc748f5e259;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cfad9b72d69c07d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e46b9b6486e2838;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h725d13e65611d524;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28e96afc0a3090f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3bd2e683e950b46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cb57b38ecdd306a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9504504fbbad6114;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58b45c62374aa1e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d635868507b0905;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc83cec2fd028329;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4f8243ee5212d37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91b89cf62c1de7a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf74c80adc7d33eec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b608cff718e8196;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae58061aeda076bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dd1312996394444;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bcb67f96ea106f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6cf9874d22838e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h310c808d3f4d17c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f216f63ce44d7b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5626bd82dcf26ef8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37688458c9f6cb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90ff5418943c3959;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39b775a493ca7733;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61fa78f27b9b765d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ea9d6f97459d99d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3524a50e125a291a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc19b9ea1063578a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed8dcb4d0b22e66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he63631a0b204237b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f410679f2a58387;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecc05ac977b94dea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7390e65b3ee7754b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfb545ae0efd8e8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdffb5238ebcdd5cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85086769499b352b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h512304536d761749;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8abfd2e3f9697bc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8acdb5fa5a1a27d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e22d9e485b289ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbd46b5910445ed3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h429354cc159a9728;
        #1
        $finish();
    end
endmodule
