module testbench();
    reg [25:0] src0;
    reg [25:0] src1;
    reg [25:0] src2;
    reg [25:0] src3;
    reg [25:0] src4;
    reg [25:0] src5;
    reg [25:0] src6;
    reg [25:0] src7;
    reg [25:0] src8;
    reg [25:0] src9;
    reg [25:0] src10;
    reg [25:0] src11;
    reg [25:0] src12;
    reg [25:0] src13;
    reg [25:0] src14;
    reg [25:0] src15;
    reg [25:0] src16;
    reg [25:0] src17;
    reg [25:0] src18;
    reg [25:0] src19;
    reg [25:0] src20;
    reg [25:0] src21;
    reg [25:0] src22;
    reg [25:0] src23;
    reg [25:0] src24;
    reg [25:0] src25;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [30:0] srcsum;
    wire [30:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3438b8d65c0b9f85bb5eb00990822868dca267adecb862d4ff3e5ca5703105322283f3b2d693aa0c76759562460e20282336291d907d749a6fff13b96956c6b4d52caa07fffa23c9be64e4844e0ec8c027a1e371;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h988d97d98ce013337eed76bb4776b30bbd2313b8072a5ac032ac0176ae1ed0ddca35846efbec5da178d2318c512123244039108b413a3cb7fc909feb71a89cd84ee252e6806ccf87b7620c3930fb13f6c39b041e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60cc7abd59e110f6b0bb198cbefeb9587d219c82c1f90de6eb433ac2c4eec439123b7540f430e04b3a67ae11e84761b2d7cd76a7b281525a29b355ba56f024cd0dd25246e71a6fc222dc1b5130f9aba8c00721587;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h892b1a35ed2b908668b7ba26c56b46ae247159515b427791d93b01d33b5fdd16a29bb19deb768c49b2ed4c4d3c26eb77f5f7707eadba36c72f5f92504f662f8b6a5e9f30cd5870e4fa55e42e76e59260d3a2dee70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h769ee584231b702840c69a66d93d9ac2cc59079a6fdeefd4e228f5527afdbbcb28c9095bd6e70644c375c0dac7cdd4219078479bfc75cb1fc3b5473ef5ac24938054ff48172f634afdc8e2ef97de7740a97390de2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72e297ca3f4db844b3e632d71dee2750f5c507e7094c3421f9d4569d60ecbccde5c78c7cc79628f9ce95c765d9f32a1ca2bddac090fadbb861bb240cd0750a1845ee230d66a29d0f0e6b9809b8b605825c0128631;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha78c7b98bc08a8d33f38526737376766675bd89d5d7625bdeff377f41f0a9bf4aeaa11294066c093ae8fa126f508d7c076127dec037204f0b34481fe2f094a102171d1cc0aa16a33caf1e3337bdae9b9105220aa8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa4c3dd2171eed9f7892281bf02f91de7db321d1d556471646bebfedc337ad71932c02dd0bde0adcf0894c20e87373a7d7e8941b8c5b2606106b836992f85eff7379c941501219152713f5659b670d2a88bbd5fc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b7ebbba6e1f6a0ab27b251e6689e5ad5cfe9e5b706389a0e950e40439751a1167ecba07f05f61f0259237f1857ce38edc1ada006090320c92277446d63ca63ebfb99647d6af30ddb1ed012f06b27c05e022f3108;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h963797558b9c47d272cd6847cd36ce7e69e832774be539326c207baf14dae6ce389e6719568772d554e9ccd490980c724e970f2fcc094cb7b747049ffdd2ff8495dfe9e0fe0ad81bfc23da2211e4deb68cc2363e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h990e549a265254776f68772701b3b36edb8e82c3b7b31c4d5e0780f57669e2cc68c4805e528393fec0671608d253af296edc702dee24cc5e8616e5c0465b538d2befd432b15b52cb21b744ab8e764bd1dc6f72074;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h298f164f59bd8a7cfffa2de6faae147b3db992d93ee9ab0911625042e4d14b85285038faa18ac3df24438b2ee3fabe12c827826e99ca678fd7a6c10cd2f195303b7ca51aec573e4e2a702f3cd1c08f02a83ab0891;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbd84ae9e97bf57d6833f468ba1926d5a2d281acf7e07825c1b2686d69803062b7e515f3ea018409b23293c765b28bb79d765063c5c477c1adc0c7ce2a24afd619a0534a3bd13fd1eb5a98c447d4de9774e8be95d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h533f23fc9a95906a859c3bf5ed27e7a43ba5840edf62008655ad83a0c3546140a52f156d0464de81cd8dfae0b8598d0c75895667ecee7682fe7f628f64b50cbc22addef2205b9ae868dcd9218c726bd669e2280ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64e7fb32236ae56638c5f3c405fd8e85011b90ff685573726d7ce4da5a0acba446ba472ceb457078dd7ca7352bae199d73320934801ebfd5084a4ae30e30644a3e4f38798c7f9dd383f791f06b3d4d97450a6f2e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b12e5ea9499240d6bd01b6aec44f6f08980f1632ec53741d6701a7d4cd210a9a795d13138d4c3f8a37d75f0fd72d968f1d72f59208f36d8dcf1095abdcba08c1adbdad0388b427df64e08bb2ed1850cb70830a01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffb0e1e5128309a5c9f85573016449273f1bf8b86c020dc4f22b10126b3713ee39843ff174418f6898bc50aa2d926683bb9e2463696a0813836242a6fbf419d34f56a40d8742e974e6e4695ba06bb62bd675dab87;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fbe5ca655ac1cfd45afe45ddf8e0a2e0feec7f92843a492a907f814c0e1d7da2adfeff5382b6084ed5d918e9fee0dfe0405de3814a1e6633b35ff629e7587b13748b5f9ac987eac42c3ba0945803f254447b01b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76bd06ac53dc78be0faedd07df725216169d7aea5a2963a2331588402c8cba7a7f2e280141c13987580c9e9087fc3f80a0e42f0974c017859d9bd0b92312c21f715465f376e81779c6f05cdcf70cc5bd27c5b4e6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c1da09106831f6cc7903f3b76d1b8ba4076337a0387d7f635da97c2834053a135355147f25f337c786f5defee83dc09d381f23115e942185a54170982c9e74af8a0166df67aa090501c5557a2301c0866ef7697c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a49d7f9789bd3f0ffecc589d592db28adca5219fb49fa19a3d313c0fd10a57546e0c58181bb66d112204b7e0187ccf19e38ca87c2722e6b2c90a941d6765bb5f59371385fd0e655063ec979dbf2642c8a2fca21f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b47b88ff7f2f438b9de3c4355ba2818e500f7eecbec340b373804c9aec06e627cb967aae53a6b611ebe97f565b16b9480b34e07c8557e27faa4dab5185891f0b10b762ae6d821d35e95b512ed5fa4fe48f725a6b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69ee51c3220e3f655f5971dae9778a24d08885c362716d545c604b9f85f0a2642311b9532078ccc8d730d4febb437bafbecdcd833b1bd752e4913f975212988f1421aaf84eddc36ed14f0a5da4b8cb7a83b72f099;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h518b0f499ae2f39d5e41ffbfc5bf67fc08c9b06aa072dbd3fb0489c6708d8150662ce885c2a1df38db65e8ed33e78b4aab4b1429989980509adfb690ee8a9c4ff88c11a9ace6988ce0902b97722397255ecc5e13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedcbf3b0a7122ecb39b07b5a0dbbd0af4750992e37e410f939be97c02cba53a6c691d10a87a93a981f4938ccd243cef79c450c541c5701dd73819f8496d6ee95aae8c8670f8f83121f9fb5b7437df206c2192ba17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2d128b4c5b239a85efe241428b30326576b8b9bb3ff5dbf939556ae676fb14a9b2dfb35b2327f7d17843cb42b5e6cc34d1bae9ad678f859a2eac42913f67c0b5363cb3d6575152dbd76810ef3dc28834c0fc143a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75acd3c79d8f21cc09e52ff3c72511668c3f4bea2b043c7fc32467dd362ad9f63603d62fd814a49dbafcc8c20d9b6efe58880daefa9806e2d832de2700f3ac084a4c27182b505dba66f33b721d3e5fd1761f31b63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1510d9f75dbc4d05cba1d2bd9e4d549c35584d01e7b64fad4b4c3a009b6e8b9896a4f69a1f5bb160c1ab55e40f0c2935d6898ec5f4d23c35e62de802aa287c187ff376837352bc3847c652c1242a583b149c428f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10bb566665e9f009e018b1b3d0a7db5da19ab287721b6c0555af98acbd20fd5402809261ebe7e105794249fab20d5b417b2ca8cadddf1268f3d53ddd673687492cbfaeed90c0fa1611c18381131da732deefb03e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h274281110386aebfc62dd3931227380769db2bed3a717a49c53b04573835617dbf9236bc6b71c16832b11b5c1a9fcc1edd132293a124def8a0824a53ecf95aed2f6eff1e3bde4f7e12e2c743d9405c896c7e6ab1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe4ed552ade8e83504a2c693ee8d42361cc7e859706a8c75d4839da8f0460913eb606778fb8ac2fd13815054033f6290270ea02ea4fa1a03b7283143b9525a5ddf8e2ebc10039dcd5bfe33eb74fcb19b3ea2e7772;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c2339942833a27a200e6076532487ab6e28b02f8ba2ee1d0b4d3edbb32714fdc3f04fb7de4d5726dd0c56694ded1acfc1d9f094f3fff48b473306c35a0ab04862e2d62bd8222af1e9bc3209a137d700128f89be7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h245a65a538595fa82eda48396c5323389ce92450022cff8882f61c8def0c3ad00d96a80b89fe532a59d17f83cdacfcffdb4c19ec2d798730c71b088a5a12916d87f0a267fcbf0f9fe5cf1bb94b28b4c95cc6e257d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd6c1e80624fb465b378e30218c1a898f55f704d14e0c713844ad6b7eca50a0e33c08ae4a77562df5f6a147b3132a1726faaac870b9edf32519409b010223ce8d2ade2a7ad9dc4d5bf61768cb7f2e88c139d8da8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48e48ce90b463c241f88d70c402f494d47565196506840dcd5248730b7ee8ec7ea54e0468b28470bb5ef52a18a76499c6f42f7281efe2d63f9e8e6cc28d101d448ac595bb238cdc08174adea64bced7e971ffc4df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dbdbd83fb4b99d61e0ff99195f53a4e58588d9183e5fe4745b2b8d61aa17c3a4e77bd9ef585db569af25135b57e27a61ee5cb865c87d38ed70938efb9919d790941c66fc7534afad704175974ed33cdf2303df9a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha84fe840d5509c01f895f59ce3755b9cca49dd18f0b595a4c2de1bfee6b2f33569129a46e63224a1945111801cd50e026ea5c9d4bb30109e4b84e01dff41e4f5e1005b8513a59b05eef5e8ed42682058cc8387a43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha74475aef650e29eb52e3a3a78d242a49a18bf189a40898a28014a683fdbb261c7d49d0fee2a935a631997b76260e4b6efb0ec15bf8413679b375cc59d28f3f9de0b714ac3a2c72e0118206b1c364e47e049bcf56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b4c14e6fb61ab523d7ba88c1b5bbc3c310a9fbe8fbc8521d416408dcd441358b4304d72bf18ca91aee9beff272d18f76907a56bb9d36e285b4bff8a36d121c38cc373bdb3839b09a0cc120bed8d84edf0902922d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc054efe793fd0e1d0665fbf7824a10ae03c46bd7b03201de678a48349a3d4806b17fdb781339d1845388a4758cc8424e6f5b533b2821543d3ca27457c66f9675dbf69040aae5d7fdac2065556d5524817812fe2c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b201861e8923416d33cfcccf0a1dd152dc0ac9cd12087e06401854bbe1c0ec891a46437f966fe458f51e580d7caaa131e761b4ff280b6f5635d122dd47cecb5912b408f2193bab279b822d6885e8a6fd2ced49ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2be3b7744cbf2a88aec2ec201369388d6b0b06cd7d525f13edaa217e6d769a97d985e1464ac002868a5a1713835008cd3b5b57cb8785ee4ac59d68a52a29a0b181252746cd43f08d07b236004084ae56773b6b07a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc25f880c277bddb8c2738e1b217517940415015b72ac4d8a209022614302fea064bb8449388840cebfdbe48168e05ecc9a236ba85a9c3ea11fec2ef11506968b3912936642cc6b0020085bfc4cd170e9ee7f2dd56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc694d5b81bde50bb7aa1a3315e559b0daa0c902320988243e6e2d4d178565807b8d4ad5cc31deffd64b3077ab8f4c0b7b5237f7b96cd8e5b3237a6e0b02e08550c91dd38200410fd7ddea8703a068a0732c11ee4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h184c3dba65398a8421ebcd02c5ff947a5ec016be776ad138e8bfe749af67074aa00d750dbbe44298739cbe1685f8fcf4966bcf0ff78b13522107274c30bfd3477436a1e04c7408252e71e5c5ba43ee764a38480bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e333f5bab2337d0ee16831d5d084ff8dbd9403d18989d6cee0650c1efe06f9822d7893292fefffd410b51cf361de4da63155a3b270df775a39de9395a11d59d5e0902e37f300f8cd3b967e1ebd7e67aadfa91c28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1629be6a71781ba4bb7059e988597ff8b571812510c70be8b9c0214f2690dfe3be1b53f4ba15c8bbc9b1c4d7a184b1946b4baf42152b14e74bd045b076fe2b5865277a3e38d0934f0be903ab1cc770927271aeb61;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1332342382b3a26b331962c9be3eaf13eb733be89ecd6ae43d4efb9f041f2e7e1833bced9cd0ca3133b9a64afdbccb14e058a76a026230ac5b9cda0e27525071761308c60a642705f9cac49ce3eaf6e287bd75e1e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8905873b3fd6ef8c9b92bdd48fbdc93b500cd4c6289bce2c9167a3a53181ebb87613579e0123978989a718a0ab94925da5dc1d42aa9ffd1c48cf86c7eec2e9ac9dd6279cf403eb630717ff297a2cfe7c124e4489;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6474e766be8153b822d33889084f8126b30851f186f567b336a2589ef9336d6af9698f654cd8126fb74303924b9ef4791dd9f7345bdfe83a32404ff143c6a58472e58c6ecf5c67b82f3f28a8cdaaa4f946b06622;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dce0cfb760e390a2399f2d7142d77c40a1c91e8cadae826af1283e3b1044557fe7bec0270992ba21bd704455dac6b6c96fb32ad66bc2242ba8bf1fc0643f1f295d050c641a71f69f93121124e0d0c0d4e4dc901f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4314a4b8cc0e460253145d0557760a4f31ec93fca9e662e89f611acd0a26408d5ff8fea318bce40245680475f90f6c52816fe08566f3a733dc2b546c0d7b2550c7478db25c4f9f1c2f47f71af193ccc624e10c2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h108caaf36a81b6544067ad2049f9de03df8afe85e34fe2356a34eb58328ee493de2160cbcb7711b9d241c66f6cf3d721e7e0dc1a36fc465dcd4a7720ff516a68886a4cf1a5bac0b8df40b32c43879f699ceaa511f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef0ff2657b4a9eb4d52dd4a371e56bd8c8b2db05948883bebb151614cae09492f57eddc9007150a1a5843fd931cfda755898043c94ac6e2d3e70de43ef9c6fa8eb68f071b376b06d7cdee418152df76a8086b5912;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44fc387df54f57d3471b3f51a465458c716e340c4198cbc8bbf7c82943d16e4a18bd7c27da567fdab3b92b791839dde5cf1f2925df9fca69c6f8a087eae95ffc70db7e0bfa5255b0e34c6f3d7b714d253f473ac6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc927595b8099896dc553ecb1cc2b927d9ba57262812e175b09d0ed17135743490bb67bbadf927a688608a545a1c5d214a34c3bc6a395c0458dc5b3cc8c2dd0ee439e451a4e9f64f0df73e9ef0e7ca032b7468d9da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19041b630e3b36287b4ef870ee6a1ed769561827d3541f1eead5fee14bd2a256a96d647264150e51ae8bf5147f656fc0048227c7da2fafd0bf9c18869caf5596513ef5979308bfc87688866be82d0cc7c67b0a1d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5262d1f73308fa6510fd0adc1d96e5196cbe83b746c052f9844b210a12f5c3651e277ac378cbb14a106a471dc2f7b9339bb22beda6e62841210f386804f3a3ccd17faa5d3fdb3a333093ef29073b3bfc9a981787b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5b3fd99ca90daf5895505ee034a4b6115bbb5b1cdc51bddd01dcf22a4a544a43ad96024e38d077f99f139a4bbbf762036bad11279bede449cc13b3f159848afd228929f20b475174d0710de71a44e9338cda1213;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h329fc4ae875be53c607e68c25dbde1f8b4261feca5686c584354f032afc566cdaa536ffff1a91a6a1c849a993aca727520247d384aa6a60b5c23b4b9b0d7a7651f2965e8437c64bad35b7b5e27e324d42680e4ddd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h838b7f45ef8df5d7aeca8a75ec4c06d6fe7405eb63ef0978f7e7528242db82885bc211d856e192feac25e565b1ec1508e1899a6857ac08cf42c434378f45ab1de514b9828237ef55cb34094ddbf0f0f269ff71539;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he18b1931ba0c3bfc9950d8288ef36c25c7c56f201cd94aa78ab4a559e457705b8be900858fdac7c4f5eca8207b8cd7780495705f2552bc1b67162e9c4f2999bfa2520995e68e63aa52b3f3a4dd297cbbe16694c5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62d2bad7fbcd23cf52f697539c49b0adf71acddba02626813b4bf867caba4f68c6433dd9f847c4ea543ae8792fba2fa95c414eb7c9d39a0c9b2a5f4cc2c08cb713db4726207a7481961b9bbe5b49ad2e2af0f6de3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7456f7e02a19c94f000b227abcd46e5767ecacb605506427e3cd39c848f64e6ff14ade3bbbb16a8b0805d76509156547b763f612a6d64ad1903c37d1dbce36d332c5ba0cd2c47a0566c50e1809a619fe5a6701207;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h621e400c7b5797d1f4daf9b3959b0cb04435b98742bc225791a9e87e5944da26eca7c4435d5ff599b1cb7c698b9d57edb76be3754c92cb3408cb86361ec3bf471e03cf39196faa00c5808916a1de086837084b289;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb51b25898b43ee74a511e99d7a3cfa5d99d6769c10295e3e2e29ed07c3b57b081bf9b892b8e471686a3804627617722ca9e01c29332eb33e9f2f2e001a0e18d0a205841220237ee82d210a41d5d8fd48f184cb7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62ca86f5753fa4e3e5466a15b2fefab3cc61006c621e41d2b7cc41232fa0b5236d9e88cd826ab198eb1ccad62788ff459871c21d7f989f3ed1802195d8c821679f9068db13702cbeb56ed9b8a4078cb3c016d4155;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h427fd7fa8d8a2be3ae928303b816a2d425cc0ba07f19db8217fe4da900e8e11fef03db363c018dc68aca784fbfa2e3c28fe011b2740d928b1516e59f2672917f82c45b71fea85a66d7b22725ba75681a527612356;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6eac42c62f5eeb99e7039ac214ce7b946ea925e3a0cbfa30a7a4a47ac7acc2abdc0ebcda06d8da2bd899d083b1ce1864b1b9e0ba5c4b362fd624c4e870c238c244cea73b2fdbbd7bf66b34d4747442747c54da68b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48d2af2d7e62733e99e5859955ff74196569e079553b0c202744de33fdaf05edaf7581a6fe3377470ec52bb81d63fce3c3603ad5192518bb048206f41fbe22c768eb26e8c07162260be6127cabd8f1cb1847004f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa1b200411a9e99299d346f1c264fd6a4588e5693956be9edbb01f09e9fa893be50ee79a004d1a98a4a434648c5c27dcd12033e1f0b4e860db00271e3e8b3796d991ae3c03acb48879e58b5d9eabd31618a9d7292;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f6f3ccb08f8c8ebf82bb6225f465cd4e4d4320f19392907de919573bcfd96d204b93592814ff8811018191a8ce4478032f385a819bc100053a827369d85a15b4ac8a32f846ebf39021413cc91e299e1c5d20ee3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cd9db816b42232915bd24194eb32e5417e519a8696f524ad523501783aa1a766ca0125c08f6805ea1aeacccec8f2436f78f3d8b449377a40fcbd747268b723ed59d807a6dfd582e0c7cc3166834efe3707fc5efd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he42b0e590a3c6d8878ea7458fc8e37a4b65c2ff173c8af01345c6af5e25348783628bf6d0a1c90b428554c90e4947ad991d68b1bc59432fcf6244e2ca50e2246fdba446ee03315ed62b7c7846bb724a156edad68c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3104e2de7474cf288680776667e4e6505207fa0f4bd7ca9d25619d3412d1e21a6b7215562b51e40eab1b6c1c4d88912e6e2ca8f047c58576c4f072853508577d9becfb8021f2c308c3d502038812513e5296f1dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0256e6f4e5d68d879818dac4cb2cc308dab7d0e1ae234c7914efeb84980287106590e995e4129df04c3f5229919105e1f18696298ad6253c4ed2f592af448dd4fd731b88be13a86205b0b55be6d651c089ef2df3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4eb2049cb55f29c2cfab4fe1752c7aa50079f09aaad530c9b146b150db3fb93ce04d9baccc8922bd367496d106e81a9b1e6d100be0a4187f8019063ab42b32f2f3fcf52e2a5d2d065bbc91a72321b3ba0d7696a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8c5d526d1b3a8a57ef7d00f87d0ced5bca99f2b60be8b956ed0776b5395dcdb5a80995a7ab58379c4647038624fb9ebbee20244344d6eef4ab7bba03bc499ac04f73f9b1d333a6c64e2ec8584b0e11d95f1e9da5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45425457ad82e7bd141b5c8dbc6355ed15bc67aafbee3602c1ff0b529df30f0cbb89125d560e690ad4209455b0cc70cc68c711ff6ac5509a337c21fa7a88fac47f398766544af9aa1082684332753c828b74685ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h283d81e0ebe9a62bf321e89225b48129565c30368e307e5d7e1a0b41cc360d61308bf2b8d069be60c9962c0d6e6217e39321d3752b35379f4b6dfd068e6006160530c323cf3c4adf9ee8e091fe8c19d07b59509a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc087711c0461eda34910aab44d22dd6370e4bb6147f785052a49d76cccbdee50ee067fa64a29cb1f2b891812e11d0dba8df6a6c481cc0a608f075b917d2327c219ff94374ab3b04969237b6daa3ab650efc0c9c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha87a226d07c9ed58d905c4a5428c61f414925f26eebfa7d000670f76a98ad4b654bf97a56459643a274376ad52f4df8589abc0d2756884f83d09c966eed927521ad0780d8cf382f18442ab54cf09c5c6f4ccb06ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h214d3c9356e095d5b0113591eca1e5856f1393596bfa6b56ef54e04b72b7c56eee8785599bcc1643b002deffd78f404205efa57c79998e56e179d9954bd7be244c722996faac8907a720c4938acfec18f5781f386;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55d1ac930bc56bd91ab3c9cbd7b8ebfa1645452e98462103b116e9197c50cb377da84ab2d104edaf02d1b0ae75f7ee0834079212d4923e498266169ffcc5f93b93b6b83d3ec29fa4699868cd6f485a40bf8c80e5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d9701633649deb401e4e2e5c7e6e5203ca49c01dde4351b2bcbdf661b94dcb85ab95452662cda0c63e3abea766a6494687ec41817cd71c48220c848919b50f0b921bd96d2a94359348605befd1cb6499c0ecfef5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h316b1aeb2e50bc34a15821a7327b95eec868f0fb895abf74834be3071c1d7711c6ea3c813768ca275c81495ac499dc8ca310f19c257690841e7fdfa103892a48c40594a1002fb3a7700562d15cf30cbcb8b89e56d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h550f79d988dd76eaef3127774ebf901900f73bc81886267fa120887ed30738d8c7b71f600e0983b30688eccf4277bb4d04bd85ad30c7ed0746458466b4ed8e58cc7bf7d23735ef79c112dec22275739f89a4d433c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f20a9301f581f966c69d60ba07ff0148141ba22b01871d687d4836888d7841a49ebdb4d6b823f99dbfd9ada6552317994ded818ee92644b5277f699026f5db309df180b3919e35055c54c9dcec052a428a469a25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f6b04c8c45ca8c264355c5caccc4702c34a0e4122ce8884b2769dc55e831c1f0831277bbacc3d0021bb2e933ad5a6647eda5ce74fab7c80e53b3161198cfbfdd9dc3e7b7102b2cbd9fee1987bc61bda68a07839c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dcab4b8d3e0d239b4f23f598cccc2ed16acd15977409f714282e26d606ab85c7a1c58f7ecd9ed7b344e5e78aff3e9a58948830c4191e407172d76842783db0f9da3e24ffe06010a2ad344b78ba02bc56c16d443a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4a2cb6d1daa1dd135526a4b1e3b87e9140dc1ebbc75122ed75e8cfc4eeaa0dcd1e7c296d9f5dd1f0111ccd803d9ec3d06a60e1dc400ebc68c4833c89b8b176dbd9add91fc02b1f9649b7fe2d03bdb3c855f42927;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h516ecf3f518fbe4648fc2daabbde7b0a2df2c692564cf8d80b86e9fa269e35b9ed4902ea7cdd03fe29021eba96408930d322329dced965b2771e661848145d67821dc80be5e7292247c531d8fac94ab276500d57f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4373c03361ae48582b0d12a903c9713dec0746646c0f1a7d9db4a81f372d526b1c02cee4c1cb8e7add49dd28c967cb9eac9c89cd41bd2b5893e8e8581f2d1acd98c86d3c02a110591c4b5314fee70b3dba50462ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9a76da6ed117fc2b798b9d1d9b32f46f0747a675c691a0465b6925d6d33a5af5e65adefd489e1d090001ff76ab29cd5a996addcaffb59dddd2e2461c8e684db1ebbf4a87ed925bfa8bebe09e3e3b26162aa1b0e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd7a2e436ddf22e086e279e30067ccfb6992b0006e398795658ccb02b7bb58320940aa85aaf43454a9288eb5460b7ff04324f372c1e22a6768388a2b4aaba114e4cfd928efca7633ad0736195e2ce1ae961a14984;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27719fc3294444a172a6b338f25fa3228a1ded1435feb24075cecd38ae4dd80f8fdaabb16477e4214226c92a1f580bbe6d8f6fde08c1d4285c163f0b9b09c886a3c38fbfa92102582d663708f68f33cf777f38c9e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd77643c35e7de61e4e4584a332b8239521e16fea91a07e978158890a6bf7192cdc2f5eb1dd16b429a734977e2e2686394fc7caeab4b6b26d060d3b5db0ce6964d0134dd7f0c18c2b94e07f3ad668096160d331a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebd1a7d1215524ca55ab5f7a7e98a702bd4f12e973b78c8228e182b7c6978256c6cd304b91893425b2eb0839eb944e78783460ba843047228d9583ef07ad1b7bf4356fbaca42b681722b81474b1eef7973a10e930;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha597053521d915e19ad644beccb45e08dd893920933925ae0d5afc9a91a6f24355149459e4f02e676eb89e73f2d45413efffe74223fceef16ffc9772ec47a241e4691a1a538ba4993a4e108ba9cd4c4bbe074d218;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35959a099b2d76ec3c18715249a03c262f26bea55f4450c01f26f54a667d2062e48b301534ac0ce5bec45d6abf34aa83642c864e98c343b442298d3c3a74cf7f3d80e374b9cbc74f72a81b0c71cc8f181250a0b88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha58a9e5d1923939372af3e5dc7f2c56f5f440f0bed29c6fd0d9cc7614c705b99951a2ecd3874f7ff8875d5d4eecc222a32a26c20d0f9c84a1e0ef46729d527b18a0efc3623600c1e105cb0b6c14b25cc7d9492d93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd0f95f607656e6fd02d5f34db13e11964eea06b9c82c8d39fc55392c252e421ec3d0cde5c52e1331a803b104c1e896142110273adeb0fc804b8bef4df0be9ef30562367d32aa278ece907f3eaabc8ca98491daba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26fc207aa103901c89071e7bdb969c3f677a19d0c4d6aac67479effea23dd5aba6c989e69dc4cea26f08ac46604be5e014662fc7e15997fdbabeb5c5f788b702b136d3b02526ff27cdb77eeb366c0913edf07caa9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ac2fd95089ea45fea04eec17043f6d5aef481cfd3bf7b1534b9403a2ee17ac24286ed75c61c187a08a363875724816595dee6608a100529e4ddf1c0d4f381c565a47cdbcb8c0f9c672b5165fbb77899142f88dfa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43abf84c59bb833977529e6e4f1ae246d4e17f186769a57eb7caa52ffa666f056c8bec11b539076752708a42130f5a7e75040ca54e5a90b73167423e4a46256b07ebbea851dd2dc50791c64acd62bbeab7c831958;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5064fd6c4ffad9c19852273b36a1d3a96a8762a40f638b96a64e4f6ebeab15fdb90ef7791c2b167b9c0bdf9c1a38afcc97a6018343374bf1cc5f3a0ad6d736135a633dd5bf1191c9999bb9a19e068c218e22280d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dc9316d738fefab1191138233783d0bb56e6bea9ea33bc21f13489201125e7a58fb3cbb4af57d9ba18c9a8f15e3634716beb1cc9fe9cdd4d9d2ec737da9cac7e05c5c699a0753623f2b9a151ccc6dd5caa422e6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h271dd3444b4b635f5ff7a0db464278fe4d11c32780cf539d528dd4107df75dd7a2de632497fe053a02eb7d35c38ac820af57345cba7f63dd5dc8f67cd1b036971d8ed9b91f10aba79fa91b1c0781643c5d484487c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7b45e8686c9b1bd32e37fbfe304bb8d4f376385508cbc4a23e5f37c53c2cee1d47c3b0b8fdb95bfb4e7af78f02282c99ab340b866d0a38adbe3a2d4720d21759d38b331a5b2c0bf8f5e10199bde91cb8cad70d0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf714b48ba3dc6a37bf648f36fa750c5aae4f3256c47acff0176582a8716c20eb0048ac8a59e354095349b970174e0a0981d2dda86850d6243216e7426c23108e645e6e96a941f5ffcf69b33cbe5806d3e61ffacac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed75de9eb63bb6c55fb9144e6f79a53de3527bf04ad1fe104b9832ed8f1cd5da1155bc17135c207f0c18b794f412650893b7fc58e35503e0ed8b954649bbe1a7ed314fafe6ffb1b551d1f5c0b46e2c6acca005392;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88d452aafa1003eb720c6d173d102078233b8d3f9ba8e4937dddd461e01b93eeb3d9d70d5919de28a52d6b6c463d8f23b5f56c217345e54787563d0dc0be93ce752d789c966dc117b42ddd254cc9db7d9578a9a8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fdc510324fc2221eb61cd7165120f00096cfbd1c2ea1741555bb6a75b81de12e0f43a405d045c77eddb5f0bd6e6837c42167f43fe08be814d4bf1e7138d5833b731313c909b19fb692710e2767e0c5d959fc7cec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68a82131d3d4597854a66a41d510613a690a2eb76fc5c733235b36fc28cfd94524337436af0a896ae60cedf3af6850623943db7f6b22bd475dca518bb8c8860e201917213a82490d51cdc24cffea4f706f1913f55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h423181d1fbc114528a08fd31ca2dfdf8b94e2c9f627911ac367f79a837b100b8d512d38c1122989540159282e7ab25bb26db1002aaafc10122ac05a32402163d0b4ea3a69031e62252c3dffafa1c2053e3f32b806;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c3328dd93bd6bb6df6fc95f3087b9113d496ca4dd46da4a0a4b178ac2c4a1dab1c435ac120c8c4d140f10e8ba7f152e61b10d5d58fd5b33ba13ab493df826085f25ad3d212d2fcb7f712968cf65c41226956f51c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ff0d082786db45bb305fc0106d71186f6d00608f073183525255dc6db89dc8e2ad6cfd67ddcdfb00584c076e34325f0abeea7013d1ccef2bb5809430f3212d925f5c53e20dc76c78079ab14efd4d9a1330310886;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87f57f6b1c2624ce87fbd05deb4d858e48e537bab4c83ef0465fde018e6a94b4ea8ca3f53ef4dc3b56fb8a1bcb82c859a961dac6fb895c9051179b1d676cfee5ef29049bd1cdbee0f0a4861e6f5fdb77812d09f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbaf6d2fcaeaf372a4d404a443134b6a85ef0fa0ffc5be1de4cfddc382533ab12417d6d53b7e3eeb41ef57397d6ee60ba916f642c78bf24ccd345400ede24ac9fd23aca0ce46e2fba5fd15a73115795fa76c2de45c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53f9aa72cff73e547b2017e141d78571e374360de0f1150d69a6cf04ebd6876d4ba329101f618c01b091379c0bab00d43c01bf71682706d214a0b9fac34ab612998e381351591edba1b8f41735a8dd11a0644aa22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1df9b7f48aef93572238518225a801da7547d58e7223ae036d4f104cb586bc15ceca6c5feb5aac4ef2fc961400d8cf2fb9e9a52970628dea1432335a245fe1755da530373b40a2b703d701133872b4cbefad3babe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadccb5d8923a0dfc0f9668615552bce1d43ed70c7c06a52ca02f3ea327d51ffb63d3d24b9a780517bbf1bf468dc0a20afa7d0cf24f4265083065de9bafaa2e3de4c9f186cf630da00b37486bf869536c37f3d1be7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha827e83da36652befacc310cf05f2f4d219c7b7ee23f03dbae45203ccda2759eee8e47a9f0bd6cb4078a905d7304402cf96d8bf59b99d310dc4cdf0321e1b98c657363d6f0c94bad990875ccf2d9dd64b848477d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he02d7d6d214747c946fada63ac77e1fda94259173d2c1f9ef6bb1cf97b0eb559f00ac1a390c0a04272dfd5673f4745335fc738779edfa06d9060e7b299c008290c5da03fed56c8362baa6462502f7e15a65a5d402;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1585a57a2bcb36a6da71a162b1c4cc5913b53ac3090e92a7d8bcbfe086d7db54a7df615bdb82a1be17b811c2432a887a84c17fff655b38de5b3d2aa355238c7d420288d60ce2c9891496b16123541a09c4ef2afaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56bff306802429de94b60da1a83e027cb93a563dbad3cc3af2bda20f52380da6643bc2b62cfd046cbe021c3b904af3f42ef27879e9f61e1e2d187fde2ce51f287c020d23c8e2ad3ac2d2f74e0c5f635628c02e51;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h681509214ea04c15a0aef3bfb092e050899bb8e9b4f3c4c0f7548dc3a57bc50147a6225e28b396c504375e32421bec8a7f2d4c21a2f69ab25b87631029a6a05e3e35e496b4d4b14bf89371a5c4d64732044a55cbb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea749d15e8255ebb731ea3d1b23a904cb58fa97238a1edea6b9d40380d3f3715a38b32b77e7b6d63c4d9d2240f45ba0b4d9529eb91c658127363dfcd83ed19e4c4cf552845a23a01abef67fcd2774e0d5e9905e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd54f37e228aa33a3eecac85ef57266b98315501ced85597a77ce7528b35384d587572fb3f831f997a8fd26508059eefc46e60fb2bfeae42a9206cf4b52e56dd90351641bbc103281eba8e6469ded16c1fa122f37e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70d28a8c68c0fde9c03f76e939e96d02b79efcd5176822df84b96a70c30b44920a46412fda68630550414c62cc4db1fa76d0b94ea9f71f307eb073fa56b492f8351154524fc1b2814dc42dd025a6e8d19179002a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5072a7eeeba3e6492de66fa971146ad8d17f5c4f37c6d600968cb60b828dccca7099ac7ae7291f80a096d294b21fb4393e19814127216c4f13f88200e649fc8358cc8b9a3f0ed063daad2ef9ed75ef4ca5081c728;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h465e02f518b1d8a6a91cab0627323cf75cd59ae73018ce87a3f87bed6b3dec559deb8d843f813376792f2665a6a2ad4dc6c89805f783139b5a5c610deaba8d689b1b6a5aa17c674c8645cddf348aaf74e073db36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h965dfe5dc4b6ae0f41b5299ed3d976820d2e9cff648796ff8823f0aa987f9eaf43fdcd09a4952832a6924f6af203708bb3c7ca7bc610f80141dfbc7a5aa3deb5a841a99ae42d45354c00c87e04be66312ddb19f4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h286b1467c1d0be30e3df23955fce3e6f4595481ac163cc312eafa988755f8fdb0ef3ed5d2cab312eb97d16efe2f0882ee27b95ffb0f5f1210f7fabd5c1aef18aeccc57417180ef433a3480c7b64f3f57a8c30c5a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdcf531b05ca4f6f92017091781a97c69678e398ca41fe45f63034f1646414e31aedbad2c2be110c82d3a4bbe97faca15c737b63b089696a3d680c96374f3881a9653ad2df81f521adef543e2863b9185c909dc71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ed5c37d40cd87a45d9af1a0e95a6ed405abc3cfdcc5fd7a13e1b75056470284ec2110143e9add78957bce7b4229ef21a002cc0254a5439818cb4d6b3fbd61e0cfb88cb9dddfe11a2908d2595d9ff9a88843782f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1849d045e12f7a1001c2c6bbe5e34a1cbb66cd450a7434d372f04375802991d6f52ea656efcb81fbec1cee6286447eff802c4d78d6355679ba399bf3fd7917dd4d2cb36ca1eebb7d197a3942868efb494510176a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h876cf59b765eb6ad4e66e18812b5e37785eea42fb3f52c424735f495c47787f9cc540874475c57bb273ffd3dc5d04fa1b2085b37e5e2f5ff92aff2faeaa4d4befd42784a2219222c4d10acfe17ac23f7fc1859017;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61fca331e7316f2eb80efea4e10c8659ef66810d3c29f06907a00b1a5ad59c002e811c8fa4b106342b992c13b375e3ee501afff8b9d37cd2cc08c47248dd05764a71b6de2458c7a92aa3988c3ad4c0b1b6b29002c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h216fc85249b1a0490fbdcbc670db429e86333acffa56bf434a4187073a1221a8b9125317d10b09bc98e220a6fcb7a36870601b9cc7e578319dafc49de582aab4fdb83037572d98057284eae6aa1322ba7a09708ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7ea5d600d721791ad3648c671ba8d430ac8a2bd4f9cdf5d9659a1c2a19bfa30c315806e33a9c91c4b01e24743072b033c1e916f459ccf80d4c2f7fb6804941ff997f1d161c05c117f49eb3a0ed78afb4bd294016;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4014bf6c624f4558da3559c42d0a430c4aa0a895a4d70a05ccb16f54215cedef83cc28bba484efb3c41d31ff15574d51d0d84dc451e60a8328ea494b71f7d86ca50a87779a5e6e4f09954095145775c4eee2a1ef1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb68f485389a421971d4f11bac211613f26de9f2ba42a77aa27932f5b3f3ae851e7140387e20ebcd9a2a69cf604fea48d352786ef40eaaa51a702626ec968cb439e5004dcd581d381128bd4f8ba0baccbdc8da80e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae72d6ee012eb724d11835a1a2fbf2037a238be104e26f3bd7bca9a433eaab1643d5773b59d869a05628f1fc017130bba1854a9f2eaea506f23ac9af7da90a1671faadb7054fa1ff601abd60198fae12ca6f189cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72d118f7f27aa1784e2ff957ac92fc10d60ee387a551630003a721eb3897026c85c9333c3f18c7826ee1bae50ee66d8dfa7eb8d895f9c60bb97004be2f872928c6c601a2c657fd8ef12c4fc86382ca6b848a3bc72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24df1ace2b6a8b4a90a896f27a936d7e5b1d89d00af5186ca08f37668da18383a6410d8ac74528289ded1af530184c16c700d370887d1ed5285fc3e99782924a67369693fbe79c0d8f476bffbf2d30ea2a9b8358b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda2ba15584dfc023a3109e1379924f1cd32fb82d43071d2f8db331705d7c07e315bdd15a8589d62f73e5aaee2588bc8b0d67e74a9f36780c19425d24c992aa1e9684896c128c532720f2c24e7b7ff86bdbbc05b7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72582d51b030cf278b42aa392d861b2e3bbf966a915acc0bd8434926756d97fbc280b5f2b9cce8dd8c56cd23b88e8c8b9203661caa0e4171d5785cb7d3fb5e5bc79b81a9e22acb10f810468d0c5f88b4a247f88f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc4ee4d0805b30d45644c755b5dab44070017957415bbeb64ab344422d1b628f889ac1a7a7d10b2eabef63347e0fe9a8674a9e06c2d6aaf970819a99246efbed6f9664bca716b18affc55d93c2b503b74ea6804e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fafe17a2e40273eb6557f020b953ecab22ef3ed28538a22a0887a3772d17e26bb5852f3ae5b2dc9c3502df568dbe41d190cc824b081fd0596094edbf8bfd8cfba089f072ed1f0aef9bd32a736a4c07988b7f0527;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aced1e8b88df773e537e12633bef1a8086be7e414ef9d2ecc2920e8378c573a3be38f96f9c746390f883e66008a03793a8171f52d7ac20fff3341486a9e857697f1e77fa16524c1fb98a7b7f4774d66c64ac6be1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95d6526004f477ef6e5dcf3cdd7bb9d142d73033a39d1d73b2785db156c2ce93b619af2e65eae75dd4b82fbbb396e8ab3cbd2ddaad9f1745cfb3af50cda044659409c28727ed3b2e2e9509d17f0b5c5c1ef5c8eda;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2273885415f5ab0604f6311b5f6e731aef97f723dd47aeecd6f521b300bfc099ec3956505fae09cffedb5a4a7e4eb8ef01412816c216695be330e791635937d035dd7ff5c48741e0bf8ac0acc2bb1428c61820c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f22e46a86de1a9224246c5f68e57d32ff259db943a53337269b2246d5306694bf5d1cfc9bd532201b092bda6428453121e818742021a20b97d1c449e0e8cc465b51f202032f28f4bcd18fae22e4686fdb650cc88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha53aad8e0f70ea30883c7d1fb75227d679ee8f5db408c0d498dda97f0a8e96749f9193f508aa32d6139ced1f54d23139d7e35146bcd93deac1555103c1acea4ca7f78c4e6423c76052fd043afde115250b3b40e2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf5e4de04a7416b5dd9a68d96a19b49169ceb15bfa15330107d773db5d7baa658db36ca9e50e77007818bc74a67189e4fb82e1284197deaa1c04915403cc893f138836ad9960861a4832c68e21e19cf79dfd69dac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha90de76944776be8bd25175fe905204b1c8bbca809787372199b60e262c2bae7f713bc95e55f035746b99e4ca4990df6c350882ce64b778f5647957c098a9d62c25ae3df046a9f55782990811a63082ded4071453;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf116be615dcc9ad8ac4b39a51f8cc12c628aad6064ea8969192f44c2e212127b587f04997d08762a82f8247a0bd68458ff779e40c35a08b42f60d4753f7a5035398ee15c5578d0df92ed6aa77e83ca66459bd3df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4160f64eca853a9d451a2e5992941b7e489b5e66ce5bb74bf96008aa47e56b00049d96f5c1e9062a6ea7262768b30893370c401d395fff49cf18258d2000815f375d18cd61a6fdf78ecaa375f29bdda3b8aae8e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96c2b1b81f2982f032540b063049e2c02259f4294dbf26ba00a48e7bbcd92db0f212878308bc501513f8705b714887c9ad1c4137331e1150f9413a1bf12cc1afdc02371bfe7687759f90114215141b9d9d67731e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8520786d33c1252cef3c10577cb857c03f2d7ef41e317137a5c36314c97f268524ef3a9c99565f72f954f8408a3dbbcc538a449c0cf1282081d74072a626223da919f1ba12dd4b8fbcbc2ecc4016fc70b285bc141;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c7c2e575c49b21ff984e0fdfbfab404f1b76dcaa2bb7b80d00b8e07d019bde3f8ca9e2e8096f91b98d9115aac36d287bbccf3c88b64adafb3c028fc1bab5c4b162592e497449074bbda90af31f3dfa873b8b0cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32ccf04d2ffdafd647d6b05b1798823813c9c67ec341262f5ad20a60f9d4f247933b95c94d50c09336d207dfd4a1ab1206fca7f01773de0c0e87bdee0aa5478cabe9784e1292978bdd65a3c55e6ea9e6d89ee779c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bf53bd73c2cc2b081aa9844a6745d3fab59a0db4eab0904fa1ff5d1f253856ac67813ea7647fa94dc590a41a9d4020efe0947dd64b9192d7c70291a7607f33e482e41cd23c0e94e4716568f3c01ebedb82759a6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc10b33588359d45fa12c6bd548b2c93991c6371fc06cdf46caf3a53f23b9941889a76d6b1d2b0c26a04de2ae18b2f1970c843f5dbbd8a6214673c669f46d857758859e2f356eb6181e1a4748764ab2ba19ef9df66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea2269751722d27cdd89e21ddf8a620045d5a20ed1746bb53a90f08a4dea6a04ff9ac9cab3f8dc24882a35cd5d82f8aa9f2976d5cc2af78ec7e1523696fc8db61b4d39cba1d247d1bd485fb7a11051770229a7582;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf186449605bfeb9adaaf8543e1acb493e8b2c02280a737dc2a0a9b429d3f30238c8d27234fd82aa708119c322f4eb9de8e3fdcadb17a3459221e92c073b6df17388dfb0ccd3a177c1b5eb0276837fada8dc48c6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19e4f15825d091d6574ab61c4224d7bfc4f41a0543a144af6493f802705629558fc14cffbe45f15c1742457e4d420e20ed31773d8873c319c3c8258f7c6ab141ca04ff85118070deb59a3702a09fc1e93ed99f56a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc63eef531a7ffe26250d8ccee66d6c4cf3ef0002046b252e015af9e80bd8c09e0f1326ae59b7a7764b1a97f85a33bd4149f5fb806cb7a3d6355d89889050cf2a9a8124c1091ae6475f67d9da8627e2d58bc9914f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc22a0f3878d293ce1d37536c46003d5997d8c91f1a614dcf41065277ec5da4b705ea54dc7622482e533201589649849530f3d8b2dd35840d006616472ea279b365ac3ef5917f542397e44250b371cdc124bba1b5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5eee4128161331d74ecbe550fe9692249d18b8c2904ec7db9f11aae961733f69361b0ec3fe18a9bfb281f2057b4719c239b03085c8f1b2275df21f7485192d727b981ff4768596679b5a818efc317a75eb9f78c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17e0619a6f67a13efa65739f954068bc5abb06aac7781722e9ad2e97a18ef40842e6ac79254f96bd158e9683543f993464615a05f472fc35ac7bf00c057cdccbff45e54f80b32cfbb638a8ce108c719f18ac16da8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0923f514eb03a874ea77242f75bf18ca2c1fe7275ee0591a016349741b063dcec33ef902e0ab11d3a4c264382ca4ccdc79648d136570e6c1f2954a959edcbdca0c14a3b45a39fc708b015a7863c4b233ad672abc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeb97c541ec9533f30c3d1f9c79bd099a272b85ef1d31d71a43a63da4cd3dd5dc1eb00dcae6b1a0713baa7d183ab54feeb88890169184b5bbf315eb793890e5fcbdcb1185d4b5b3597b7428079e15986656fa4036;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75fe2c654b67e38acd09b33f4b87fe27621ac7fc023c81aa8b3731cd149eac2603da6fb364bcd6561666d17845a4c4483cbcc8569cb2d9890b4a4be2fb06a2638044c40b6f597ab753a5479619e62be2b0086376d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9db62ea796433e0376ba145f5a2b2f2cec2e855dbf07ff6712da82554545019c05536812048629594f781c8d045d4e76c9f535ef5099c085d8c43a96cad14d508a03b4352e384a92bbddc8c8c8451a7e0f6525d54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80344ad840d34231f70e6f63a63026199d18fc3d9e0b97c1b20938be1985968d5a3dfb7694aa5517b1f02bb3c99bbe8244817fb1f6b224faedab30e855ee1cc36c69941b2f4dcf0587bae1fde6956ceef457273c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dec3d52777e78fa3d20309680e4cea83fead3d73f894117522cdb2c1071ca2ed64d37ab72a7a87c26dd0a2ea4d505306778683ddbb790ccfdd65d7f4dd401381f4bc6971c4bfb0bb2857687cd0251aab42bf011d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2ad441c09414478ffef06e1931efce90f2edccb0aca5d1e1cfc4447278fd8722c0bfbb6e44a037f1147c44d0fbedbfcccdac73ffe1d69b5cba61fa7a4677d7f883ef5578139724b4390d524ed2b5cef0e71c7f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf7643971b9a9d64325e93b997107fc6af41c55f1bb0d750549a3b145ae96f8404b7ae823c4e1144f1b9e51b8d89018183a22d8eb30e4c7c265421826f751ad444e3c9dfbbb28061e60f709a1a4e3441ae7b2579;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfc4dd4fd8067005dcc61cfc8e4574f5b77191d0ecca4beb4f208a35b227a2594f03b7383d18be67947d77cdf0cf873281158b233621bda9d46514c2747a3ffc5b053353ccb3e1e230da08efae777ac00d1f38a91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21b225dc212293601f039c752299241bd0e2ecbc8c1076d5fb57e5766d503d016bd2f6cdb68cd5659cc788c476b8bcb001752d19b1237dbbdf705dc029a3514541de8b14edf688d46a1c2da3cb77f70e368e50fc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebaa9fa8676a6ae66c5d79e329f4d6ad0d8a7a6f34191e41d0ea2170fa5de46dc16826cb49b9464399154d3fd142363b8b558c0482f5383249bf4cf7dc7edbb08a405fb76e4f0482125e6f7cd4cca4c917ba96c5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e8e564a992345c868443527633088381d2169c42a2bab29e127218d0761a729d7a846d395cbed430fd1dab7288c3d365de1d24ad2675ab3bf90d9ed049339d9c4da676da476bca8b23882c822289d60dc01b27dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74abd4a8791f4fa49f5aab38629b39d3df5f4bc279d5530bb6b6fd4721c4fac75ebb1b6d8f101d2b0cc9b008bb36f56f9b42393467fec3674c54e2863a689afb6c294c762588b15c90839b091382087cd782e2766;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1558f0af4b1d0164ef3a6d00474b86d62557438a5a50a5137e6acb2ee394ff21c57be2305815229da4f116111e5d77dec7d1c08ebf9825eea7963cdeb0884e91f20778377b01d20ae56dc0c0e7a9d78098fda83ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c012ef68e54077ca149012fa6d42279b120e38fe94ec4eccd4df6a4dece0d4044ac6e5dab2e64607de9a4dcc0cc34aea3a4c17975bddcd893e9b28d9d8a5209e6c08e6d4b3fa9a27a0197f9c89b98f8f907b0f2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h989722d6d09fd748c8a49410c94f2b84d7bb14cb8c8aff0dd217c508faf4d2135f838e19e4bed05d3e956049c4962622f630995d0d3a949587fd84d4967e25058bc88f8cbbab4fbf5deea88dbd9ffbbeecadb203d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65aa3b189073f0194a9009cf5a7dcc40b82c0ce1b61769449c4ee2b832619257d0c608b7e2222bb2ded0e89c15e647957027ccef8fd83b2086e5536cd23b023fd86315a7998201ee5bddadcf0a7162f86f8836296;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ca4dd8b9751d07d7ce97a4b3c63032e24763b805d6bc2e4d301a3db90539df29e6c07bcae09fb440ac863dd31f1e26e0c80cf1a91d3c7ab37a92902710a4a82e21547d1ca73921c7daab9c6aa164c3a521314dde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a54cf1e9f62b31142817c93aa403de4b2473daa5bb7758b36f35ca58d8ce22f4aa97fc7b30ffd486eaf92bd143558c2644ee8949390e0cd45eafbf8486df454f1dc75e878196524b992d14484e1dd6489fa7af1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4442583879eb347568529e467982ad0f75c956941f6596b924831bd57c5e458c1681439bfe34f1628af31fc87d87e4c6a1917d746f8b646552bb3e5468b01524f1920a1ce345c240d9e341cab2a422419cdc6df99;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76a9d8b22f956b47eee9066e8316d075b7ff7ea57588433595683dcfedd86f2a44a6b229faf53a8553f710da7d0d32a9ae366d231e1da95b02068ecf240da718e8785b52e0b9b9d569853a638724b16fbf753ca43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc68d0bc4d90f8c4c8ca86cc48b07db6a6ca37ac8753a417e135c343e8ca9200eb81baa847923147a9e77d3c4a4981863ddf1aaa186208bf99ce25b4b756acc83c9819f2b98ba1b5299d53b27926edbb6356b0b3c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1101a8e97a28096261329080d35fc89d17f0f0d716eabead9e7a88176b13ea030ebe9ad12e1d480597557dc4be6358f933f87c282ee8b3e21d99230611286f67c75e246cae4855ca8b2bf4916b04288c31ce51558;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3078187c2d55306d776a35e94b3657c84720dd75f3d2d3eb8bf2bca134a7137e2bb81c0fe9c17ba9b3c7eebe5bf276ed0b0b82272649dcd68757cd871ffb78cf9da3078778336a8facc5d4f975948daa23d7ec27a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f8cf069aef908497a64ab4be7bc7876e4fedbb57548beebac34aeb1a07cdf97112ef499bc7127eff714d8d6266ffb6c22f5b06766f8dc60e6ff2ec6dbd47d1d8531cf31665864cee4d99f83aa50820fd60affb64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8955e765744436abc9ba6b95a1c6591d23a5884c7a7e8f1a25e10b3569bdb00023129ac898d0e837075eabb113e6dcdfff3fa4538a9965ea31d9f1670fb0a73df0ab1154659b5adb7bac09ec8f58e9e84b53dfae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ee89005f66e3df92fbdbbde1d378cab081d0737bc8e7ff0c84c194d7639980eaa98cbe9e2d9738f5d69ebdf96bd6cd9b9fe8efcb30f4de9328c428c52dc10fbdf9509599d482eafded56bfe577dc5a449f111b58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47d016bf11c8754527e949be668a95b8d719206880d3e15013f18872cfddb887f2a2e3208910fe9b1f423b1b2d2c80361fa84f7f53f2b8973fd467d595705c7f807ed660d456429be13bd6e0d2e95d77da20a154a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bd42acf13a9707dc2361e2c3c215fa024370654c3ca241d40014adc6344a4e114a18bf349167d790a66da2647ede765a61729c17055a983b1d3d496bf01c75f3a555f43c0404e25bf93dcd71f5ec54b332580579;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaafbdeacc7b21598fcab48d369986ff027055ad9e6ceb9f29ae3d1abd178318fc0d5dd52baedce749267eb1ded130a641beb8efe8275c08c7c78fa36f302bbb598101dc384d8307ee942a903d13884af5799f38c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0200120960b71c904988c904e91ffdad6377ee21df19ac322d04660f844366c4c945aa8235109d577893aba312b30d310900aefda686893bc30ad65490aebffe8ebae85627dee207e02d432821c7cc6e7f20a7e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7336e2f2456f90aa1f60876d955a0252dba23f111c00626950ca17cd8c64cfb7a5b5b09b0b304a02150a148d6df02de6d616fc016d5e632714852b6a40da65a98c78fedc64af10cfe7412500d76c40cc3a23e685c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3442718c63b16214206439e9b07e64c94b2f66f701ee47fba1282cf827cd662a4f99c0f402096718b01dcbfe0563f33fd47222950330deb68d23b5bab4c6329c4ab57e5761de64b632ef536d17f15dc1f858cd2e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h965b891bd91a4f99c6a592e999b703825e9823e664c86aa2005b5a8e69bc8fa3a1c4bfe121c5066cfdc218ec21cd41eed1354326d1a912b57f598e52b8f826946abf2965e9b8816de2b0da7e2d9c37d5155346ec5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c6da242f1f6d3b32dfd68fd844f1d74ef9f93c239a1cb3be65a63eb2d3d789542730b48637064106b3eaa32a349808ccae5f7b2010efa39ac6d270505333c4d533597ca35254105664ed9c8e32940cdc5d410820;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f7104d65f7b4291d58d9b13624813f2268db0045b9dc320168fb7179dc0933526bd50fdd7cd619fbf45f7d95182ae96b6ac41b448fbb414398d32d5029732cef3835c140e8f5363ca1566f4c674d1bad64a43248;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h217f726173efbc1d4d906c65d3594e90667f37f866ca19fcfe696f0663d365dec3fbefe290b9828ade1f08c478973728969a7d6251aec58c67cfc8da0a75c5422ba8e67e557c67ceab02f2afd7b19f2f656cbcfc2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45124a55f45b7bdff1acddf45f6681122607d2f3dc04e762f5043d1195a9d451cc47804c1b0076434d483d9e687f9926b92bea63df15ccdf424bf63f37c10059eca08a567677cbf23d0667444f3dbceb90114bf75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b35a848b9afaf8c4f8e801478755fd1a7b68fdf0aa64895d270c7f6be6f837d23bb1d9ae8d22f5132153740496a9c34606a90883b5fa914ec83482c2107ab3a09ce246e4de603e294b0f49512ec7a4b8392049ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ec93017c44a219cec83a6091a2852705083e1ad382573d4b38072f72ec276d6a907a8e355f31ca2f1684534cb6f460333af3a9852ec19c65ecec9180cd7afb5c049f58ad009e52e2e4e0506cffde53e6253cbb31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc36626d4a1be4b57c65307db38899bcafbc194d8bcaa345e64553e1013704d51dcacc0b24d0b26addde2601b0964bfa4e38c773a409109aa942f50a5409958e391dd437f6090148e193e18b19d19d6d2821dbb511;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd3c4a414595364f421945ffbc89e294124cb3d2818e0b458ab715db63d56104dc39527a61366a237af33c03af8a3600c66ab3acf500e10a7422a32222dfe4f8b17f9423912a8558fddb6e8c914b23a1b6938e416;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cc938d72ad9692a57805a6c232bcf427007b3558a5af4de9e4b195f735a1d076b680167dde8b609242be952ad6378c713eca8b1d9b9c46aafe534cf30485cec18ed5041dafdd37d2f678f763c808ea6c70830a22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h195b43e90aa2e07c75d9e500e8d1ac65d0cfa472f29e2a22cf3722f903e2f8cf4c49b4bbacec823575c20cca447ae18383e935fca69566c6c1df81f4e48fe4a04973047b2abb27f84bb717e402528a6220e885b8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h399fb699cbdfbde5951e31fc01df6e8b1a3286f7fabf5b7425ac14244d1167a1904544428800d9d323ba9185ec7b712048ebb9e1ab90253bab10fe20b0a4761c9fab6290d43b29dc24196e464c6f163a5958a32e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73fa6988661611af7f8cafb0d1336a726bc0a8050a56f2fdab54a3274432bb529c05fec894a99cc14a9784404fb0786d1e9de6c3bf992bacfe89910f6e44250c6bf1a135d401095816e41cb259b2f82389c30e0b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33fe416a46c4558728530569b10031113f2bbbd2adab110493006fe570de2cf3a680f60e96a42274d3c0e793e249f29c43e39be96c1b07486afbcce2cd94ea7eca858219aeb16694e940602e5717fd17efe08dea0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h569218ef6ce5af3322d89121e3594b6126d7f180fce8171bcd4b4e5adf8e41eaa39c61611f61a220159a381b1086cb2ea8d2ab92e2dac1c3dd523b3c4f4824d715e682f260b03defbc8fb0e143d798d0692f003fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdb9da53b71f4a153d52b892dda0ddc8472fdadf7843777484dfed0cdc2e6de511ae48442e0677fb7c3778c4ee0572b527c02976801a40f25f9bdd0f4c789bf6641f315eeee9528b1e5c5bea3822abc3d5de4cf3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1aa2207e77a3b283abeb67c684d68a96260a346eb7d97699c4c6313ac3b511a64843aa1dcd2128766538f22529b6cd1c6ed7d3c971eff30352eae4714d740478e03efea55f561a3711c92be929818499ec7490970;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29800a2f384d62181cd0fc81442f4083a5d94c716fa294aa987746241ee3d889903d30a98e211a475faa23e29533cafc843029b62bae318349c3add19d2c07b3b4c6889a75900dff5b14403c9faba08e89e2aeb21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc4d8186997c9c57e26c6bd36938c953df3f955dedc2d369338d1af86b8444bbcb73095be735d05e91eb53a58b2b81e24897b2798ea331d7f75ec7b3a16ad7bb1b6e6d0a388fc9a0e640b2551b4b8f888cd7eee6d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62ba378775a88f515955c581adc7202592bbe9fb787842551708c78cbc5a2bbb605fcc878750e7563d3e43c6bb14d7426768d405800ee4062ed8d0fe624f483a8a6bbccc7fe88dd212455dc8bfa3cabdcfdef05fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf781c2a37e9d4d5f82d49821694487eb81064f7d6d6b94ba298f4439450fd54ae66d00893eff9602a194d1d82093eb3e6ba5f5525277885f49c5401b97da83088357972a9ac4d2e89fba2d5e29e9f860917a5a640;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had4687e8ea38c586002ff678846550da7bc8cd349f159dc33a7ded3fe88a9379f5b5ce9d36895d0f6cba37391b57add500496868d0f0813ae8e4e8235c304e4a5fce2978cec971abc6ff35740dc22a1b6375ef492;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f3393055dbda16caa48ff46694a61c0a1316b32f0be3b689901414aa2e166ddc4d8bb8ecec2beaaf24bdc3aa2896bb38b899217d26b624c03a44054dc131ab5d6087347559d8f4c996a8616957ffdbe65d8124cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb197014c6cb10332ce53dcaab53e60ae86830a673772f945a20c6b012e43f0bfe7cdc02b503604dc0aca2e2fe69651551b24041dd0f1468def0e2188cbba9e461fc275938a1e18bd127a7644b50042289b73666e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcee4e37a26ee4711f3c57493366746b95ba6164d73cce910ae05f463b4cfe38b79d9b48c5e3d989f5409bb3d8e22b2cde74584dab1a6d6f61ecd4b0b84a20d492188668cfed395c16e247534bbf9c22d4bbbdbd40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55d76b0ab44f74fc403c1e9fc6a33724e58456e0c8495e94d5d17d91261f61cbca48036270305c9af51e8cbbe7a5e7a943ce323da570e096019e952cce5e9f11d71aec31a58954bec9656f546d4ba3ff97fefba0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb28c22bf0d6db72e431452ffdedeb6042d78e54b590c14cd8d86e21a25164a8536f69f63be7ace7b15d8e84abe2e00a1edbce8ee58e7181865c767c8a7173dcc7df597e6a794fc20061bbcc42b4ccbd741a5fb321;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec6816cd2ae6655970892f4816818e041841c5ed95763abe9d8604cecb9f8b17dc19278db18b156c3117ba7b5671da5acb56e7ffdaa692e69d7bb65fca878be58afe566659ab7ce62bd77fc3b87ffdcd8ebf653f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3979f7ccdea8cc418524cfb71e84953933304a00f388dee1f2d748d3fd33327d1637668fd1bf705cabf12cdac1ff951eaf8f4c2de2e9248995a294bc2589b56c7390d66e074f1a7d9340c1274db0fc1df953728;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd7b167257b7bdd68439141cbc33c196c155a9438dc8ab8f2896ba00a016ba7fe3ef274b3290cf5e68ceeb1b8904f60fa88ebe9fbf6e94fcf6e77c87e2e6b359728766373e0dbe1842c1b125e22babfa53bbe1e90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64490a091a23acfd921037314ede6420ee9d1d6437a6cc75bc923d85da3cb85bbfaf71ee55e839f07bb76850f7ff9c34d51d18f95a5f332f8a64d7cfaca281f66378aaac7ae6cbd00f2d71bf1c660b41e5e9fe326;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78afc9383aff4c03ee32f6086cdb2ef32328be00771d931ea30303014b10a6dbd8018ec10c5ad5c1eb5c7f16115f987f20c5b602f20fe0964c957ce2247394da4b890e10a9150e52e296e31ceae7b7b738dec12b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dadde8a89b2ef8194f541b66f3707f77bb36cd3baa783523b53d37328586ce01afc003c86ac468e49a0fc9aa13d58796ce410b4ee78582f0ed2c9ef722d50b3049d008b4425d4bf018b918960f5b4987007d2314;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ec972d6221275f2eec9e5e62a6fd38d9183438b7ce0047a05d953a79519ec0abd574d1bd46eb7797efee1216005818ad083441962ba131a03be062d816c5067aadb0783818f278f20b01f5044f2deda5caa8cb03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb22b42fefccd08fdbe3507c1aae15cf8028a9eecd738198d6c05543d3cc99555a330b290a4b99e5b8e8bd3f0ed1fe3f3b135af1c30f63ab9ef3a7cd8c3dd58989d2c34c59ce8fb5a72661bd4e39030c4da9d1e8d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h303dd4ccb8f69b1e0a591087e9facf209c221a6ed025fe99f52d5a51af6b5a9b2162dee41db5355c15568ad61ff538ac4dc26cede974f4d172191f9c020aab0d5a26acd31cccbeb407fc8ac01e64ed92305e901e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h826db1b4a96bbe43fcfeb09ebad2d80ff83b91bbcc206c2d7248488509446095282a3730eecd80c4aa6fb0560b68660b0a0130b67dbf126cdfc91d23c3bb315fa8afba11b8d60f318e940049b2c4835d2e7594ce7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde104cc40cbf35fc95f892209e423171df8f781d19f5162256829016ba5b3ab250f27eb42d79f5d3b91501747ddd7369899b287f2b2beb814adf00e57eb701e63374ade90c995b473f8de60f041284f138d5cc7b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22192a032309520fb982f0b6bf75e86aabb84fb282875983decbf85e2cb21a452e45d1268afa3b644823ea9381c3782d7556041d6d04175254d7e3085762e010660ba12d91d78d57e6b01152c5837a0d4b1b8cd0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d0560aa1b416a8327d8e19d076baec3d837625c108d6c08c309b82cdaed187ad1fcd6a1309df0c00f1445c0f435b1cffb86f51e1ddd09fb2147ead7eab78d8ad8003d237c11c00c5ad0dddd8de54b7b56d68add6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf2a244e9d58e213e16b6dcc682b24fc3ed2bdc5290ec85761779da95d4f9bc9c19baac3b2d08ce87fb828818310b37ffd6a328eb103c95637683fb8b31aaeaef3cabdfdef7b58caec56e0562623053e522c2cc29;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6392aedbb66a6107b26868382b4a3e619ae75b6acaa9cf3c12c231b0a88d3d84ad026e8132bf855fe44559efd94e6f03fcb17c888b92a08f74ff7af5597c300ec97141d2b2d220c15caaa866f9ebc65c38e1a2f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46d65587705d9d324408cc1f5354352f903d7393ba0a8ba7f01d72ae8f327d601068595e1fd87d6b9b1b6365a9621cfcdcf82364f0c473a7e49d3d1e21c3b99827d67990eb153c70e0567d649274201c97dd2522a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h933c03e7f1ff1fecde42b6a8e66c7a289578143c62c9c1eaa380a33daf785d5145b0beb965ed24325e9e2ec007307202ea94aa20eadbffe36c429778ec0c81100774fc30d9e4229ba46e55c7685b7fd43f9cdbe54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13712af9595ec1aede3c65901945bfc07efa511f355840fd3c93ce4f9e73f089ba748a5f5a2bcc2c5b6a27bc9ec026ed765a09a4b1baffa9c00a10301af94c3d56d96d9e33d000a9beb42a24110611aedca3d145e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32c1f801ce6bcabc1fa5d0363960e993449483c88a6d8bafd8cd6f0c55d1c8f2f66389223ec4a9d0e2427e685e5fd3c95455c92ead4a0e119be7e7f65bf06edede47eec31df1cc105e9705c9ecab5f88b201f69fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b448b3e8f2a3d53c45e73c0ead86320798357663f3473643e930eaf406f8c8258ee9f632f6e29ca80460ec693d7b000f88fa5ca61f7bdc6c5cda13ec0a177e232d661cbc8b9258affbf8d13ec0a8e19cf5c90f48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc79c573cd172f228bf26b4b9041a4df7cfb26ad4a77b0dd9de9d36f382e97f85a41c8b505af7f32a1794736857733ee48f5787abd0decb6714fe0bfd205d19c078e18a8645c9f3e774f8dd135492a250ef511554;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56f2242fad1b06c8d830274fa9afc352af538f46c9994ec9682dd0f4e0dd7003d2d2f575b4fdd592c9410f47a96782eef2bb5a529e88d531c1bc8c1a4bd8b35336dfecba69bf0d8781ea3aca71b0459f34a77261a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9affa8b86a540a52b56c9ba8496707e83dbed56017f79f28f994158b1e7ed60916e72c395756ef38a07af2f5d4ca536d8304baccde0184670bab7859bfabaf779911ffaed7574aca9ae723925dfb6bd5679188e76;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h833502af3a97ee8626662cfad0756c56d8dce0d9c0fd459ea36e1e35e0ac802ecf6195e5394a6b1a423fc97420ad3f4c59b88cc62973bb80b3ee566cbdd7e2c356aba1e87ad9e34bcc840765219f5ddb20b496938;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c0531732f6117e3f13154d13b869554661762e4fc6f39d9b1a77182ac04bce06157b9c06b33847b1cf17d91829a44b5291a9d88cb66cccc64a13d09aed4751eacbbf1ebc8d97ac6077801f668493cf90593c13ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdc8bf0ee50af5dfaaa0fcfb99116cda29cbaccc3c09c4352e81df86273542a14fa1582b1d8a51204d680879ff54e912c1eae9cfaefdab334eb47fc91eb89c0469a325d638a5e7c7cb92afe0f48b53126178f545b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda2eb22b3fdf8001bcc6a8b3dbbd3509a923710497f0a68c32ed9c4bba01d1da3328fa0a81af5d375b3c004a0a487e6ea3bb529e9d1e089e2dd8c9d92025a5a0e95edad1a1773f74b14beb53c6ecc01eac8070df8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec96dae860c2bc1b524582d918fc93cf2f4bc610491507bbbc5532b4101a3fc1001d596ddcf5e79282f8655adf921f7460362d92a36a8fc60b724a1057b3920a515daad758003ca7a86255f7fed69b43c8b63fc0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he99d2dc6be4d8aa33da831a359e9eceebd6e525efb0ae1ce97692f863692b70cd0a324e3f9cae5a43f1081b0b15c5b187cbc3da762b0ce9c7c18055751512ae0080c74fe3abeca46f5684ed1dc87af07e911e6a23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f6fa2f33d20e2a00719a9066a603cd7efb7d965562ab6dd4f190d06e57c16f3ba4f3df11b7ffabc570c404bc179e6ca2441ee5a4c8be1e9c4f3465d79bc312a88a80feac0c550551238177ab0ebe42c6ffb3f2a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de852230e3d7a2aeedd264c1dd54f2dd9032afd4ff747f5588d95d1fb8a7899357a803f62fbb0c7d0691cacf3f6a5c04540d22b9fd86453b693c069fde0266177b5d81cfeb7f2ca59191fb66a25df327dd24d359;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff9a8a92405cd0a986959af8796a9059c8bb1df46946c378e8cd4e008a2c9ec75d31a625645a3b2c6a647a461330819cd4ec490b05d381086f428c6bf38917b15ff18261b4f341073d208e7ea94d27a0ccb1681cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79c5f494ca9f65a1bf999b56fd272330582e70313fcdbd6e9fc4626c47d9936667331094f890806991b5926215d87a18de890a2bc389c5553ad27ee995dc128ec8b38938a8448cf2ea52bda30803a3b0e221aabf7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e7d1ad9990c883daa365d269ea9351004375b6b82774efba2cc2f0aab3cf230b1d54acc55a8f45aea328cc998af814eb7da191c6a93ad767834e8ecb9f2baceceec9153c1a5068ce2f9468dd71a732dc7485074a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87d973c8fa287f29fee720b6520d5c796f0c472e14553e6bad6686144124ae760e72dde77d0b6b97b47feb0029de44f4553119dd9840b79fca2cb7563b8aaa27fac218214e64a518074281bf53111b3ab1b529bec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c53a4e3d30d50d591e3a9002c25adc44c7866412c0f63a3cd9993b6bb19cae407ed1d89a91f79a5bb7557dcf5f34daae6b4c2ac54b607d6edf8e0245569f3850c546660bc72271594308c788d9d1beb34e9c153a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fd285e4d12ac82d4133916d6155dcce556ac674379a37fee089010cdb07ed7ba32c4d91206a06c48c7c9395dbba030773294429d4228addcfd3c1064e90dc3b7a25e1fc48a80b1d0788077603c7c088a51fc3937;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb2040dbc4f809ac7924a9b53504886797aec9c8710e5ccb9f89a355571cd2b5bb2f8010fca2785db655e25856841d365befafa61b44b3136e038d63dd01868a935bff27f6d81e8c39d95f59c772d7fdbee3ac8a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h733d2dd6550e6b9fa86531c867d8a5aa7d937beae1c48b0542b925665c1cab803e1ec670ffdb4a09d848578ced537da5e873a2b77e17933a056781d4f644f63257ec3548e2a6005091befaf6243640b96ad832e50;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha366684eca9b49d44ea2f816d8934bc1735e470a9ee647cd573e9a9e71442471403b034689ebf76caed8ab7ebdff8210fea54c8405671505b8834fb2a784a116c83ad923cdd6b004c9b686cbf27bb2236f96cbad3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb5a2415a6f0ba47a2bb8deb92e20f60c293ac4a0cffa1eb7bb1a122f26c82d6e2b320f2631892120cff6a4b1627451ad3efd72bc5de8730e666a79e6fc2db270ec4cbfc688637c8b06907553c60ccc3933c69945;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h715b8140dc96f591af7beb6d921837f58fdfc5c02321accfa3accfdcbb8681810bead169987ba6299d5edb202fc5446b08a30cf42b1d3a388f356c13aeefeed75180fa9d950387f66aba90d82b4cc3be6e6f60803;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34d556484d346fde4ad8047dcf1874eedc5db6ac568f8fa94c7dd397d03f373ebfc6db9e8fdf92708296c7597b5fa591441ff18842d2db8097e9666327889f3856dc050485b747af55bf1f85d054feb73452bb712;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d5bb16a079c0d5241dede5e3c8810804d247c59ba8e9d86538ce7b76686641bdadfff5ea0fb7a71af215bc90ff2524f231a18bc9d3e75b0acdd2c885cf27d95956d53efd2816d109cc5bcca680d4ad2ce292e4d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h319d9ab6bdf22045c78d0b65a64398085ab3377d150cb7f2e8a554ffef3b30cba33f841d74c6fbd3acfffd7253216aa7651a0ba1013f14a585fc5bfea8cf727ce2fe19413265ef4328b574c60bd4c1a61995c9cb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf59b1d682067f212ba33540c26ed53dc4246369c05a9c44e9775f06541f70063f87c45b445373113590bd7bb3ff0966f359255bbc988268a6873933abd5e5674c9522fb4aa6f3c683e68afcbc651712fbdfa9f13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c0d3f356508ffd299cd0c9139844de0b58914d7c75b1a231e5e58602b42ec236fca15c42349385e8a91b469fa06f8274c193088f0abef1febaef5bc76714349af54463c639bc542cc7bbe9c7e5279c15e1727a57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h417df56f4fa0adf369b83436de513224a37086ae9577857308a972f129967445145a62f6bd095e387afa3682c6859dfe47da8b1efabb69587395b592ff23bb80eda26770544fbeb0bfe4195e8fd7d2a17a9a2ea58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f6b318d7489d7d3347649885b4adefc9e32304e62d01be86a03ac97c0c3dee2022c3338b852b9674e6054ee274d5042c6412a17c6c7b921cc8041ae83791a3cc5f4bd28e381d552fd4cc36dff4b0f9ec5fe84c27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f294f56eb723e3cf67c35442fd5710f9e6357f10298dea3c7a04bb352ea9f6a47a2c94861f00a49d475823cd7a5be15ba6cfb726f30d7e3d6544d4f8f879d9eef12ba0877a23e7a43ce61e78870d2182b849237d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h902f697af675d4d6ecac6a73b4b046175ccc07419a2aab769527ab735ad83c4fce445640411e715a9470bda95c62f967a914d19dbabaa759ed1878430646a71253a8fb15caeff864b923187a8ff158b4680d62c08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81ec5d876eeba0fcbbe4a9eb774d7d55ac3b86555a0d4d3e270ac4cb0a04eed1c23f2fff805168953b6ebc3ce5c105c691ccb0283e97492bd759023704953e926f71f81e5c7c1c3976246db63105c0657c6320f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47569b661c90d66646ec45cff7f0c4dfeffe30ae150c7a1e28a5015579ac8264890bf6c1a3eae2a324c110f49cd43ba34d9bcc5c382c6a2b15c916e8f6ca89b69303773b020c35c3edbf003827bd06e24efb1f314;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h269cf81d77ca255e6eedc7be78d65352b05319226b23f6cda80e95179025425a886626135014eb0f4a3d66dbf4dde2e7b8554548f4bb643d6b7f1681c31ea0d3e14205cb66f1fde7a48a2dce39b4f5c28996dbea0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd21598039d9210595737c5280eb5feb5cda1620ae44e30185833114b38738fb907eb55580831221ee1534d3bdbb6aa3dd30165a94572fcf1024a3c96a5dec76c6e74b6d91cae0c83a0adc00682b2ccff21c4bb968;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cdd9a8e51eba6e7dc3514a5a169c396465c987fb44a174b2566d3d262215995f1956be682422b0da9b524694b77937cc50b88eb4dd0d2f6ecd309c51728c48542aace462ecbc2f4c2d573fa38c086791904f9b95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c1cabd03c330401b9fa561ac37c7f03bfaef694a585d3791e01ce7a3230347dd710211eba960d3de824f4ff181a2a7a1cb5a68bc5486289994513d9bb68be1bb510ad1fdecc2270b3cf3b1af2bfe0fc6f5072ce3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ccfef0ee6c69808202316c717c9deb141169ef180d59bfc540f30be0588961823435c279ad53900b530f2ad077a487778dd0404316d67950698fa3c5ae286ee15be0883132001f84e5a4608e6c79d32c15ba7c3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h380469feed01d48aa2a10ce06137a7334489e36d8e3552bbd2427ce83a0e4aa50fa955e92cd0515798268f9697abedbca81464d0851fc699909cfcaf6bc5e4f8268169080b5543a2813066f6879abff593f24343e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77f70372802271addd062c2e7925f32f2c41bb07529506fe2084128caf8c4d0d9ba590ce7f0146002191910caaf37bf6387247a12c4ebca6d2f2bb43651af6c79e02ff409635e0072d388d6f635a7472e54a58c4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f5f3716469074de196c33d470882a407884ccc758cf9d66c036449123df4b9f0d0b1201bd43ee0b71186229ddb713aa0243d0d870216b89e6aaa3d7d4567d61aa02f1d60d150f8807e583526552a0cb60a201db5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb965c7e658be5f6cdc8c4528001a8e3eacf90cd4c3818240cac525140e4bd60c834588b70c30403195217ce3aef14a5e26b64418c898ec45cef322527979f3a5033c3076d33300c52e6fde4867522692259002c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81b64c4a7c06b384db19880cd1775e3c5f7ac04536825b5645f1e72228b5f4c8c749796b5678b142c1f5bb4a95759bd0fd09d70b0967e305076600379e2d9322641764356624187ebd240d9ed8d3a46103f8cab87;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb15cc47080b8245f1b27d1563a98ea987300770390a6837a98881272cc7fd50e366ee2f636978d4fca694538f6e52ef00faa87f0e1c429b8544f81bfde34c858b4ab25e8910e52d777ae27bb654089eb9cd929a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he62542592509f579470910aa9de6ed2663100d8418db19012974467c3bce9a671a21892aec3a37203ba0f2f7ee1b277369474a5c253f45ed9e5bcc30e3178feea9b2a4fcb13d9d84c626f8f6d0173cafb7b58b108;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c81ce5dfc119f3270d1dbeb5304831485fc2cc39f452c57c728c68dcf93eb7d4f6446174308665d88206f05805cc4f724de1d9cd5e7a5ce3af978054b591160336782930da0a0abf7f8c66d5d0bf1dca4355013;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a67c8752cbe6d189564f33fe27af05aabefa40037e24c7d4f909664ece28ec81c875d5cf9901171fc293750538cbcc58884bef22707df2828b40f8afdf861785a0cec68a7524e309dc120e795b42a508e6de3f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c5f4c87eb9d566aec7c92e5ceb85fb9b6bdd3ff7a3a3f6439246d2f5100d83747622c7f07618e6b7479265e8aae1d421e5e01a349899f555af952e240f0987f10de851913e8b7f53eb840fc8b56db854279ef5d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaea9f0a10bdd7d105f12297d228fbc198ff22e4415c17347d060c4dc4d9b744784416b4dbb33b00ccac03a601d1b7e60dea2c6f7d53e7b7c76914b8a101c11becd22bc553af7df96218e90d2264c2b0e12fae797;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82fdc3c9268d3ae37e6c3fa9a8202be89b11475528e5f5c302eeee109ced6db86afefb4f40e14e4f02e94fdbdcb2cc081b1fda5bf95b1fac03beacf09763f270ff8ff5f8dc2781b72e111f330753a14dc6ed4ebbc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fb428d34321a942cea0078c0b213fe54e5d6dd18fc7da3b896624a1a107b9bd483e0f0bd2e1efd1aee8ffa373f6f4e6c47a5e54974a8e2066fc0af690e5ace941d38d5ce80e0c912b9f03d58db53e1c6e203d5fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a558ccbe13665bbd75d0eea531ee3f345ef8104afd85447c3d53378d1a3c662dbfaa27bec94f984734d79b68c5ad6b41f90a86009c30dffe487209cbad2345f8ba9d103ced292d7ff9ff45f9e40c11a2b26901ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfde64753d805cd8a16941630c6f0229c27d81cd1e30adb4e42aeac72f19f3d23907c76f87ef158647bea489788209af1b1b1374b9261cc5ea4d67b8f856e961dedfc9fcd6ba94f5dcae85a6a667407e7e4a00d4f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdba6926a2e2b0904686140921257b86651f5662729b597297d06c9fa5ae25686300521746c5b054bbb3b3da3ee501e078a747cd20c091aec9dd90b52e64d0c7ca8dc5d5c68b985476f4a1dd31b92419169a42223d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83965a90c8583e9fdd87167bb777fb1d9de0a1d3f2d41ea756b3c3a55cd685dabee65c1cdfbc84e635331f38295233a1cfe184252bf9d92e34fc67af2b9b1ec624762795ff71f7d3723743acb001b19215a4c9bcd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d1655d77eea9ca5ea23b4ab04e7c7cc007f61ce7884f35d5d810c64440db9124cd2306ef8edd5f5217455774c0fbca0ec95cfcb85574ee1a53b55d654ab36210712479f86d6bf11fb5a082ec3e0d57a8e593f6b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he60ca2e34737fb543c4716c6fca8f00816a078087d0312bc5017976c23e60037fe3ee224a3cee78e55ce8673b8a6787a8534c5b5d6c8e7d65ca85170e927147ceee6d99a6791f8e2da9ca5c3768c630a68008d19b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43080db0204bf141b05bd791ed0ed246135321e1698f0ada220f47ea165fe5ddd72ffc352651116d7169ed797026bcbae4390aa72a9cd1c6455744a1f223af7f5f24311aa2c7f337c29bf6e5dc8384e7642b11063;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84be421c4916cf7b850eace85b3572e2e1a2a64a3a2c7ea742d0f5be7f37bcda317954921081aeba7690ac366ed9c21504d883a56e7fcc38ea5b0815cdde5582dbfacf55043c207b174c812a86e009cbaa6a8c230;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d0b8f53c9f89657250eea3d6ed14bdee7c2fc2719b892d920724b87126e49e8c5e64153efcf9dee2de167d51debf8eb4d813ef80fb98b29ea2537af3777b0852e7d71a9f31905a3fb7c31fafe1ae7d33a1a662a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ccfa656f88b881cc4d1b62528a1bd5a0f88dcd86799132ae515afc34204bbf1a370ded8e91d0271f6459ebca397ebc317a8f4c0a123232801a204acf0e19c0209c82cfe3a0a5accd3df0ff2c7dfe31cc2aeed7bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda7a818483a354f5b921f6dd62cf33cfb5f41f891f954a607fb27485d74125a7fd1a8bb632e3c7e170b8f93a86968551631192557d5dae8a9259413e4e7380a4401f98cbeb52cf54d8b66363f5c16cf1e12ccf373;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92d77a0b9917ce886ef5ca65b6e5a036b306ba723bd1d55c60a25ff7fde0e654a25a76bf480d8ab0c2ec9394d1ced0573b3d5310361f215624fef10afd6a59a51c11a444139db30631a082a0af15918c7457f3f9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7babbbcfbebf84e1b7eaa27cf46e681d4cfa6da74a78030af93e309f20b68872feb76513de3ecd3fe6c1beaaa849a8e5c3a44f9350074e54a26d29851828f3e890323a5517ebd54c01d53ab33c14b24c1b76c9499;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h316eafeb50518380f76bc044795995d06af28fb59b83f3c66bc3db94e6eebb3e15e023b7c0f82a9ba8b4e9a79df2c2d04629e5b8266018d439a9cd15fa8da944e26f13c6c1b521a3ec453107b43facd42e66a6d84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82272e4343f811e5bd1f65b45217f9f45336acd5a977fc7088583fba323a6144301b637f4b269e5f6f71ccd1247863a979da6e68f56af68ffaec24048344e0ac83da7e1e575bfbdf71d639001c2335f5c046c66c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b263f8b30cd1e9c596de3ecf1ea62da70ee5eae1eb2e2502e39e93b4c69bb2909dac43b4d73c4222a41dd00f8034579659a2f4f6978a340f0334e5039bb31f1c1ccbc27606a0a15715b22b2abef43443cedeb30b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3c7b8ec01f2f494055f5bb90100482fa70dbaa4c9a57cadb0b4453b848dce2c55206be518cdea0e8cde2f54154c119830b53e223f941ccdc0db31d38a68b35694a18f84736f22f53a389b3e95ba61d09e8376b57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41b18529dfa3433e45b1096cc0f7630b913cd54bb61eb8dde487885935d173439ec81e94d07491beaf5364121b72c8edcaf6e83183bbab589549570eb7728ba464ecd04debe020c99b01abb24c5c8af107f5aaacf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb27482a46bad7a1a5101c3b3c8ac1a9400a364a0ece2453ba34e6d9af41a54c05bb16ccaa9b7afa71dd8e480702c9e70517af0ec7dab3bff94aba52518f9fe7fc049aca2b72947972d4334e5634f6c699c78b7254;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9f3a37dc8cbefb0cc7b1c9fc70472fee226ac0bd41f7d3106995bbfa8af6ebc8135bcb35a04d71966efeda7830ae869a0f8d56bb895e3e54d1ef4e7dec0d37eeccc5cd2e8aa3dce0192dff5ad4ba13019afac076;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaec685481acf8ac1a781036a64ae6d5910d7d9516462ddbe02ff6312f6b752d74c19aba282f0d02cfd74f6ee1eba245058a73b1de883d4d1adb97908a19339dbd24f759b1b3ed5685999165ac55fbada3aa9161e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7b8e768fc99503bb8dd109878c1922a30e2270e1b4debe6ee434f0c64d04d18aefb520f92b4f4d303aba20791f6c14985390af42c8daeab55114150445c68095ae3da3f8d7ee00a67818af8f1b2ec2d8628cedcf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacab2bf6cb22edfcc74572b074db3bf8e9edd3c88e848c09564432f23a65059ba6592fab184e6ce4a3cd4ddafd9e7ee198300c618693d47954278f7e8883e2ea3cd4ca64817657d6cc2d3df80d2d75660fcaecf84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12e16a3202da91a3fa92e116521ef0ded03814b95273a5fd64723d851c94078a3f8f51f3b2180cb27eb84150654610cebaeb90f876a7b9cd990b705901a72b9943546ef79313447ec8b74bd5a55a051cc013a8d6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82ab3f143b3d383ee594d58ad922c5baab58d7a4d1e929a300ae4993531f10cde1f823df8ace66dc4ea0360de2b2e8d061131831e46d1637926782de4fdfd349ed62fb9dbd200cee22aa161b0a4c2a6fd40ae8c24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb43415e8f4df3df55c99a1d3f8ee18bcff3d019caf2925c23dfa046b902b3c2b1b239ba58200eec5e36b22a4c94b9a141c77f7febf8efcc3d5af174d7f1312d9b1c3544ffe1f3e800739b0c7d12361b711cfdfc2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h146b9d25fa47c2f4d3aaf9eb2312ef8b746b354883f53efb4a6c9aa03ac108992757bfe9e1127c5f569b3868ae2c0cf37134b0bd62452b7251956c741813f5fa25843dabc2fec1994bae4e021efe5ae8962ef5a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f384055ddcde65d59e7c65a8c6ba50211b3543197c093a948e01afde3dba8b94de8bee00b4f9183e85175f2aa1a328e7b27e7dfb9061ee75a379dd1b040800b62484f202dcdcd95ff9163caff568e3df8e74a683;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h350fe0f92e1f687d0907e3444d235f18f064d33e6acc5203e265d8de56dd93650b334a93458f01f6b38a9c7eb590669c875f7f1621eedd89ed8732b39d4572e2bc49d12f5d06cbedfa8729faa3d16e25c0a871107;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d67469aa8456ff7fff76eb6897fe1333be87571a1d78ad9df2346475b7fe99df5b4dff71247fa35fb93986ce6650063b3598bd7a1602b4adc3040513add9de15dbe10d2a8ec491fa973399c3ab8a28fab7bf9f7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0a3ae7060f3013ae0f2056367a63095d05d764e7e9ee46d81f3ab281067ae6789b5d35e633e9042dc3f8369107e9a8446d8ae4e4e0d1b3de85152dd8edc0d9d6386c2e929284e3dc446ddf0575c9d244926b7de5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb459a1af152118ff21412c1b7fa02c7b8348d812c8ba34faf2b51fd6793cec1bc392dbfd8c6cc9a0c01587d81b2cbe392a58206de55cc806b9763cb55aed4cf02e5e3fe7c9b178d54550663ab241b54ce6b4048b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he33918a0089a4d5d7f033193751ef7cc77fb7111bac945de35f463d912b3827c684017b3b04b4f2b687fc2c7dc6258c5741577259d43a32339c307a11f26a05a0a4ad6f092fa414abaa23946755c9e2f06c300c75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd67e312d5e86d63f192bdf571c1234dca61bd3cdfb37231ea13a3af1a95a2aa72add98b5041de2ef8fdf5a80fe757719e3354ee421163a28ab93ef99343946aa577bd295286248d04032ee8fb53c87a59cfeb216;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18e7e0a882e29a5f68e9626107bb5d9e54f742a0553e62db682b4b80ad172ec0cbdbf53e10c22dc65af3b72bbe0a6ff57e7bdb9d80c7e63a559693b2d58f90bc92510210008aede6c8c46fd468dd1d25b09354302;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h100eacbd7b836c15ede521805f92312ef5a727e578e8b66448a902116cd80fc16a9766f9240da881b098ef003e2a941c760275fce3d1ce9b8a75162ada270e6d21bcfcd9b1e192bce733254641c4844103b94b449;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h501df74c9508382eaf9a693a6ac05e0938154fe2a620ac49e774abfa8385f91287853dfa476e8eae6b83e34d93ab96aeab4764b6ddffcbd0d43a73a3ccf791bf57732cd6237071c794d32d801189106e6949339b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24a5414bb21debcefc2a984502fe849ec8099070dba6c92884b4b0dda4caab22c5f613a0a5c9750a9399f727e9dcb453462e706a9ce966657da1db35901ffc15fe7c4aaf58ea02655064b910407da7d8937e33f95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2b0a363d0f4f21b6dc41f516ccbc38c8eb6d16a4cf4f84edbda1354580e1b8abfc8cf33ae29ea05f3438031076b7a566643ed7b30c15423808443c7bf270f2d5f5664e3e56235d25ecd1d80b283fc2f96d36b791;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9798a277e95dab61a1dd60c0a70d48577275b1a2cfc172e707dd3d94ba5cf1f04c557d556b6e83cfa8943c26a20abd63e2f8632fbe655ada00ef5753cdf065970b4ed985acecd55ea972dde717546aedfe65e315b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7362739e28bc2e017eb321e14e580c4d14fab38121cfa0b36f521a3c23363be451e227e95491f3d45431ee52519c02e4087b6af0db7b2a56e1f441f56e5484c3776d0c35034c857dd995283be440c04e26b09a5dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e8e37cc2b73823f5b4550fe0ad7bc7b9b254482f16a76f4e8e5558114a34ccd099ae7fdd2072ef852fe6f93bd4169450f2174ebe4f918236cc0a2924a58269489394a01467d9b2f972f200002ea7557fb5bb7ff1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1aeb505cd8fc5c3fd7421931fa88b78552375b6adc734039fa8f7c977ba991f55b5423bc97f1245e3258c535b5b49159b7a076f9e1c07598a1542d2afa78a81ca2d159395bd3152cc772fd97f45a9861e4289d56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1272072b6717ef5e4735c7de4ebe5358c2a232cb786ae622238d35eec575272afb34eea3f4bb58453d89b337c555d64d3a46b190fa65fe49d0c8f07d93427d1d937b86c6c02f254e52640622b8e7931d885aee626;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d94e7fbd92acd8e204b10ebf859d5c2dbd508234253b2dd44ba3062289cf4f2746ff1bdfa0f18e26dd1dd869a2298d1c23d1d01f9544f34466534100c457d77910619022dd45510f7582b6bb7e384cb56d29eecd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ec920d9cf8328765e4f13fcba9ca817be985e98ba162a06f8f31175476ed6b7c9ad9b4c0141de82e1e1b09156135a2d75956642142ed7034450df99fa948aefb335426458ca2be8bc93fd19935749178413a28d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57160bd459963168c8c0c95ee4e3df308aa749db4fadbac3b4e6322fec7c25630e9db60101af56f7bf291099bb5b057b143cfd28eff79c22460c4ede2283871eee813000e19786ee383a2506a53e6eea660c6db68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f28669e4ec67cdea6a6ab35c57067905797ef5f842b4495fa62d65366546f9bd82cc02b6294bbd06f797b24227ba3c7ed25232c61e9e153f28f5386dcf8dfc6873a06b1cf199e340b13d2d55f3db3e2fd10b546e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31094ffdb48e3fdbcff6dbd3e233de622e5c7b40cc3bf5bf491bd3923607604f27df9678220d8cf31144067e0b38375866fb6acaa10a21fdd348741a2657d6e91ed2f17801b22ec5e60f957212309f16e619c221;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fe2cee6b56778f17135e6729e40b53d094aa806ed93df37c386e0e40ecc07b7e667a51ac61fd7b8b3524a391f1f0a11edbb28895b73bd19aa63d62304144ce601ba2d40d3336d130f5d1c1774c0a39d4bc16b5d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9454c9c4e42dfef29b5188e8af695f845d08858dd4cbd5f6c29acd5680ca555ff8ff0ad95adf2b716a12336d925e6731983ecca5e59d48fe2bcba73c9c71e483106e5c429b95ffe70b2887f9f7a748070c3cce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf983f66c37d8b5e713d41d064feb9d80a772887eaeddabcd24e1a04b0231f236a87534fc68148ebe969ac7c0904efd874ffb099494e42818c9586b710b4e929d6cdfd212e04a2d86ed94246183a4cf96b909b0af6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ae2fbf0ead3c40d764c527148d183731ebd8b01fcf881dffb4c6cc72ea3981fb2e0b5edc4bece4c35dabb9bfe72c65d767d7f3d01e8a192e5a0475f599d4e90d7b5dc9d0025d458fe03bc2c1500591ab273aefcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4011b04f636b8db90a07c2af376359d7e3a56a9b009de4b94035bcfd7b4a3a21d29731c840950f1a6d8dfa2185deed65d2a66c090a39ae9c357c90afc2764d2b643f970d6884b7573d577634d360b65a38fe9d094;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8d3a4b10e2a30687d3c99ee842469530ae88344d21da9f066f9c06b3edbef915bd81d4b73d516285882ab6508c4e0410b1f5f606b84e62ec58bc1844d3b17af14fb5a2ba76c6273c676d9cba95e49ee0ea028649;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddd36cab72a30a8e7a25619cec53ec67227572d0153e4e7ed976f1f25c88d6dac98ba6b1b474eec423218d47b3ee6b04fe2d9b00c7ca6f3622ddb2638b474816a967237aa029f8ad50468f55cb59b604d80122cf8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5e5f8524400bd1dc217667d8fb2e17713015b6e8bf87596af9d7e25f3edb4b02bb3bbabde0f4aa35f25c70b2832882ee7bce2a05ecf1861611003035072be72ab0de5cf2038c621fc6fad2590d1b91364788c21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafaa9fa35c59d65cbfcc857de3dd7f7608ae08769b27637cbdf1a4d84bd858d7bf6e76d9c165e3691cf59a5965bfebd12e4130eb51950d999fe7d9aba5ae655b214e00612304713c82f851b76dbc73294179f9853;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h527eac52f524db6f8ceded06ff4558b2c7d9623248524373e12f792ac6c68ff74105a9a8943ad380f5ec079cf24d192ac6080eda75126f2cbf36102697d4569c1359f420be44f4cc4ddd0c38e4dcddda670518e9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54ba754c8f8f31dc432e62895a8419519cce87197a3be35efc9794492a54ca0204d32f8a861e588eb6b5d348870716cf977f56e47962f5f2b532f481dc69e00d93ab475f9b47b6dc41a7277ec575c81264ba54645;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8994a969e7fef26a21c63e433bb5c1ed9fb0ab6ef88726ba5b22a232e35d6edd2dba373f6edf395387ee682c5fb756815b3aed32df1e3218e40a1425311c7f50ada588e81924975fc8f228aefd2dae8f78b9ad8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cc05d4fdf52984b66eb3fa27f9eb01ec0fef10d0b5835f01fdb74b4254fcc3d168a059da2d25c49ab54a346563424c78d07ff4809384cb5c31e159497567fbac7ddb13a9ffb865de6d66999aaeec0847eaeefdb2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a47e0429a80147bbca7f6f78c0bb9d8798599c7176b3926bd4dba417c6752ba679b33d9c0157d60332a3084d7300b656d6c7f90876034efa52ab4649d18b100ba74dd4dc857a4729288fe3dc06511fba1dd658d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d7c8430a2675f4220862250ebb63a2d8e8ce5f8ee306f8834583ceeb36cdd913952444b265145c594c72e2e60147d8f0f16bf365a64ba8c2f3bbc388120afcd7529137a7ece2d9c34ae461912cde9f169a1fdc3f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa99ca28bdaf3adfa03a9f740805b584ec3051ac3ecca6cdb7d14aef676a28e35d62493d7b4e195df473dd27673b6bfed1dfbd3051d12de349cf63d4a1a66d344c4c340dc5a1d20f3d1187bf5588150147fade89f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea7c12fc917b68f523d7e8e64b8bcd08195dd958b941f61c1c1e6cf025d7860c2d2d6298787ebc6d2634ca2b0b3c23fa7497fcf64656a26dd9e51503651ff80ddc6675deabe138679d7c9d6d87f5bc352d7c52a40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb82b68fec604493dd18dcb9f46d5e499de648a450b7c5612abedcb557483855302f5d5a7d1a84772b8dcd7196090033be8351e83ee842b725a765c4beb783f1dc2b5f3ec36287d85e7ce94834286615501f4e2d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd1e1c6ac58b2a7ef43894eefbc856f5621dd7842970b5e71042b6a967a421f12e1594f512a4880538e11197a7f81a4f0be4cddfd29f224b5a077aca9d428342c57eb79da438a34718a345b71621cbef4d71b7580;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21bb3673593a67d372cce05d27779709fc064a1f637389e5c16e0fd4f168304ffc64e6cfeff10a16a0383b677a13eed39fc2d2d6ffbcd21a5a89f7d0bde7453aad0e20863cdef3d09e58b72d1582f71a645c9856b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90c9d3a6f8345f2d05f1937f0529e7a79414cde0f97c8a16bdfd7288f5f07853a9962bdad630d1ea36c74887e3495bd5f93a827f3a8952a064e6b60fa0b677ff1dd97db45e17181111ee225afb347a6ff2c0233f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc966159a7e4593373c7de599ec5e855294676d9cc534fe209ea222ffe417bab1f6ff79895afdb3ff4f74a054780bae32245e8ae858e07f8aa15acee65825fe3736324c9c818525530ba699123ec3260703a9e3c5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e929005b799c08d02221acaea80f38e3620d2ac7b1880392d07c6dac4cb983252ea6d12cf781d0693cd10db61d59f20f7228b5729977893abec9d850b90a48795aefca67cab7c5fdd12e655a6fd0567079120f37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf141764bd24caa256c46542d08344a4a6dd7cc9c689b646fb2c701e6f5906800085bbdf65679ea171c86b9edf1216584ba912a9506bab600fcb9ea55cbc7d7d098130369b19819aae798c95658d8b0bc29df159e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ce5ea6c15e725b9550c507052b0cbe06fcd794c0e9db90ba2b1478edaf40eeea688d27629332b077e256434485553a1347268e7c960a9f0425b7681a89178fb5273123237666b720529f023d1cf4a9ad4475ba03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9424af40d5c5cf5238048e6793b2197787f869a73ccdd70d39da27d32dd64710a2ac013b61abd907d0ec7fa1a1c212a6ff8bbf53dfdccbc996186f2424b9ffae80f968f662a91e876151a905fddc592dcb93243dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75555941e11f4b6f555c036a25f237bd6c141f929340017a91e12d65e44108409c84c18dd80d6e15f540bcf7a24290301d1ad60bec9e1997593a36bba41d1717e7f75263e3de55c6c0e475aac47cd120d498d7ef9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4074d7aa30fd3f06c2f24fb6db86ddae0de45b39dfaf63751626289f696be7f644d30820471518947772980f5aed43cf2e8d68405374181a6860318d30140692b3e9596ddb813bf90cde09315f90b3773013d465;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a87645a6e238256fa555b5a048fd3defb614c9c8c3499d334b6b140c8de3eea0fbca2b9044d7dc169449741baa6632dbb1b85f6e41fbe01042ab7206dc56dfb419a3ffb4bd97d9578edd2c01c170714f66b3110e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69e382768dbb48eb132cdb035d96c22cdcc5e5adc094de3bdbd2bd9deae59633809674d225cfd74d47e21a36bf1f9439b3f0d746adddc2a3c3605bf8234d9c607c5c22642103e2615b896c32c137b746abb21714f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91bab7d71706d2f69356a50a12b1ae82773ebc5ea7d1c204d084e2653f1288b533eef6b34c65b6fa17ea99b08cc1842eb50b20f4de65fe2c7b4d4734b65988d0b3e8299e8a8f4633308238c5bbb90a363479a1197;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3003db2b873b946fc3919223b22b5173c66cf8f9f909003b04e01699ddbeec234a76a8a4ecd47fe21b0d5d1a06298e35f5aa924f99903b72d4ca7f3ae8566c76c5f61af3d50a0c2957d12dbbb526131d1ca729586;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb9c5348a76c373e8e1ce380f6d08a7f5142641e18167b52a00011136a3ee6036bec217c0caa72f42503a333505fde714ddcfe0030dbef5a107003db79bb8040b3281a15442f8d6d430f584d3463372a6a0371716;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18eb8d12ce711e8c2ff59d1607a4fd39dfbf2875d3a1538ac3c6dbea674955d2200ce70b25148b7b6cb937324405dee8c119e25dc5a5213f6f80ab6458c66be1986b79614ea068792fd36e757fbefe99c1233ec34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3fe2398ff02bbd2d00270c48b5a7d16833186fb3b5abce0f4cbc1d5bff3c21f4c90bf6eaf3576d6dd8a9b3f0ce9d78f9e825c3d8afadf84d6b7ea9293373a89241c97facfe5452fd1fc50f3436ca18455cb1e823;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7cd067195e8236ac980d3bb36545a6e38f89d48fe002a11ee2ea06b4dce103c26c62ade6bb9a812e38a5ebb5e881789cc498fa1aacd71376f7279ca468a1de0c71104a08fee14e3a88c8c700bd764b49824595e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41372cf193895e22fab48dd69405662f182db7c4ccfa373c29c4f0adc5bef9f4772ffe6cf1037df13a6f48fa4b3b9342795fcabd4ac8864cb6caf2ce0a648f8a183415a18213844b3e7fd87b1a2a79d55818cf473;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e12a514bde7c636dec6e0b985c544efe684ccc0bce3240da1d302bbf18dbb08f9ee54b6a762a8822370c207e579a27357e08b017b33ce5969f28a4888073d34024d49d7514c6c66f430bd2a03ac456e99d6ce8b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c112c6da6a4c5db7a104829a00eef1451ed273cebe65569c8f791a6b70d25396c4641f9e34f189d20852f0fc87c89a5cee748d689234411f94c93574d1f6699088a46395e9e3f865698ca334d1c40a6b7c5c2a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86d8b6f367351f3c8364305726bd531fa15c0b8bf99958e59c45ba84d9d75516bdf9c8253f5bbfd04ed2babc7dd7721831dfb3e1675a6fadb0b97a7f79dbfdb7ae1076a6b25df14e57520aa6b6df4f0b23d4add18;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e51dd4a2f6783846dcf79181ccac508cb077ab11cf4899862d4e21a707f612018d42e4adb4b3c2187ab10e5c7bac1e4378f05bc626f464b8e9f4a84e2c17d97d6fd5d2dfcb1c74d6ed36f7db2bf6940d8750f86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64b01568680d8f34d997bc4f42b6b5f86772b20fde8f5c9429b7c668edb5459a8915dfa97c2b52f37d6f890c517c721ef3af319dd389928c85815811495541460030154637ccea3709677f15bc0bd4afcdd2570fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h341025ce7a035101424253c8ed4d0d7bb52554420b749de2c58fba236466fb5fe6e44257afeeacc694a4f5ab96bdc9d86fde2e01317f653c1029c77c43a5001a03229ab7821b6779be95f8325d50694aefb21b78;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea10bc665090760a696b38c78e3c106b5585dc276742b9242da1754f0b1c583bb03aeaf26ce6635899415f3d666eacd1cabdce7f59910d2e4a52ebc4385420750a602951e32d671e5c6a8dd62cadf85692e2d56f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf536577fe8fd9985350fc5bb0578b784a057274f9a96b57fae9b33450811577aa678730354a4896e3c0351d23dc7f3b85f0622f4f7d0cd56ab88e6383d55decc3e81e8619cacbe2b498d4dd3915a15de7cef5d69f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha02f08b93e5b9267257a1cf606d3014b20a9b7cf745e2c70728eb60f8f006b0903896cc9a1aa4fe460c670caca70c6d25e0b7bc572ebbca41b6da01fb9bf2d181b03ed7a4d32ae2ef82ef3f8fd16a6d0b861ae39f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11448d5248e8ac70fb6ec699532bce4d5d7ae107943732c77761be192a69e2bcc7bbbd00c474ee501200b85bc5268a16e1540487c17cf276946397bd4f7edd7619c8abf0f0f8413b74ddfb87d954cc5ab31af0882;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf480b2dcbdf3d78f4ad5f545d2432d02fa5e63eb8ee2b9ab7d64ccce4932568129b6a4e4d6f7fd8a6414577e9829e4215082eda78eeccf5e097ed43d14ec1d245a9d9fb2155bc352222f290ee19ea545ed032c985;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c296015262cac282093bcc2368d2b6177d47abba52d8c2c18270227580b00463bc2e6fdaa9ab2f5c3b50e67d2a78aeec70780b746d0ac658ba89eb6baea3711b633ca2b222efb3714e00e9bf6ceb7151f62ef1cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98f05afd69c3c97df8169e296bf829a17c664c059454fa1b01318a57c354cbc2033853c0f4c16b8bd6ae6095d856158b247c0245c7e16dcbd92ebe1dd4593b5267ff2f97e1c364bc7f399adc9a15e45cca4f1d01e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8587553a8fde4dfa420f137bd81ec62c7e8cb3c6ecfe5fcd4e5971fe510f676abf0df603c99fbfaf39a3e8099e8021b04e7ab7dcc23853b7090fdccf1a827e2d5ab743420de322838e7b0d9e98d436e82e4c0ebc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c1eb1ab4063c1d2b39cdfd004ca77ce02cc0bc30510cde13a0f532cd13ad446d8dedc5ffe391531be2f2c718fd093340739f36781422f62dabd79d22236bffe6b4800ee4fd4b2af3bd8108eee0affde71bd554e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf6f2a601b5302b825780a1e72902c3eb91cf4b3e35111599a21aeb593518e330b37ccbeaf6ccfdbd5c40af2ed0686b69e875bbb86bd5516aa85f26ea5d0e60cc2ccb7fa48e274813f4f80996bb6d194d22a366bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff6788aee6277f732f77f1bf5bac1213d63e012fcdc4a06bb85081588ddb017e161adee8837680c3a957065e3836dd5b680286174de9f7b2e98a64945951319cf9c4b4b8ca6219fbc078841204440dfcd45387668;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0b9aa670ce5f9b8ae819e930a8c3e5091992ea873facbf106de94048618c0e86d18435e9bb1b8ccd8e94ebb21d58470cbaf52c06c3f8936c9dd4e9fb0c14fe335c14bde0d76cbc30552b0a7bc5c4b28569798fc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h845931af0a07cc3563289da85b86420198262f80685c6945823e1109cabe25fe79f2e0091e4585789f73c24c831ed0b1e4827d20c2ea723a24c3c0fba01b192247807ab51b10b5d2a876d9d7b93a4b85352551eed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde32f36a3662ac7c4a30c71ce21edafda589898617369e18943afba06bc6a44c035b7ec200011d86471982ff9c1010d6274891b45089ed66696351d62098967555498d9ef487311b93f82d7f631ca02dc81149a19;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81437c5d5ac5ee46b7e48273ac00471962c15fb8f0b16465bd0f280840cbea643b7bea02f89f708119b5e473e4a00ef234db3686427cae3c9aab302edb3e87dc23c1f26509f62aa01782f1822b462d281ec3fd465;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4432a610bd94fdb4fe6e012fb444887513bd91343499c6032d87f023edffe4183ecb139792d33dd4b5a25c6bbe00ad74967da5280d7834067802d03a5298ef64234af35a8cbe2487e3ba1d9f5ab42f0a15975921f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdddbdcfa9bd809d2876783cf511b1137f8db51d3d8bf56aacf1085cc6fb00e689907a86184601017209fb0634b1e2cd3cf5e9553b4e574929633974e40f2b2bd4dc3024bf82fd4d6da9b5c921c785adf7e706a563;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3116e9d5eb9b5f3e6f110e979d72cff144315cc0f69246a5b705b464b954b1943a3294b1a091fb291d1cff3b786456d7a2bf0e8da6853f56768d6c27b678c9d972d2e010961aaaf53001c40403ea01ca74780332;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha26bfc95a27a0bf8c851a610740b994a1acdce7a91a35a1f36c452a22be558f1bff073930b369e975dbfbb9a93d7a1df5b15b8a6301a6ea12bf67f0c22a8f9dde56392f5a7f408e7bd5b802c2dc62472090f92168;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1540c03bf28593653dc08fad34278347f5008e4e5feb027ff5c1bcd7869a5a127436a36ee89b42ac2018f3ae9fdd4cf118a02991aec391f595e1c2d0b2a8d463e258725d637f4b9e790a0317b45f56bce6c4abf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc39282d02192b8fa95be3d1ae4305036a74754e6e11d5b81ce603a600955e769265b8a87c8d5fe0ee2230da731277bb2791aaad4b78156a842cba65296212f0de76dfbce8930ccdbfb3cd399c988f32a0b6c0fbdd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3afe947f1caeda8fd950aebafcf74450692bd2fb4b69363a9498e56c8df8743471a9e4cf385153c1c5655674e6a47bb1f3e0aaf55d020936b5def13af13e5d82cd9f824d7ccbbb849489214aee693f8a05d6ed12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12ff86eae788028bd826191819207c4c850b24a3e46794a67128993cfb42cb5139a88528c5b42d984425a4c3c969f88f719c9ad886cd7fac9f70e590e3bc5f493d22dbbed78cbe2548f3d90df01f0de2649dcbc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4755e420e040899b24328d9d5350241c87ffba84ba00816aca8509356a5913ba4bad91d7ee6a0b48875a0590be2b9994cc17db2889974d0dba474f4469f26d8b4f74b93575064fe4f3e81e35c83f5e3d8d0ad27bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cacace6cacb07baa679320074741458f4907b2f4bcc2ef993b602f2238e7dd4d35f7396f901f866b90969cea9d131a1070c9fd0780fe2259fee4b286732a3e166cd906370c46c648189c0bd67bd427dd8365a84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d70c52bcb30cc92c30fd9bb360e2b51bc3550a513fa48bc3062d6646b44bda14ed3c12e878c546c43fd93e6da864b347378f716834673fadd6a0366ed9af73641eee4e218574166e52b4b693c6fb7903d0f35582;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f3887cf5f8c9f5abe6086ac29b8730fe1d796d017834fe6d92ed659f4559fb2141cb0f2cce7db478466d0193e3bc3345c18595a2966d6989a68743761d8864a0793dd59c206ff7ca355ab6f318caefc9e89be5a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9027e4bd040076624a4e9570a2e7bdc5df7a767b3a60c1e5a04c95e2e8e94fdcd7a2127c7541c451e385d1e34c2abaf41048e39735367d668e86d62754590df927f372e788387b6549aa32cae7312514401d5408;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habed5f61092e2e154206302107221c500df1208d4e3492de3ea2d12f0af6aea23b59b669020c27319c4444949918af7d64b22212324dbf95dff799aef552a5269af8f7b782faac76d003d4a64608eca72f07bb9f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h401ffc49a5a88c6e5ca99a47ea92f250b0a5ab3eb2acc6bd279c400b26e3250fa9b06fcbfbb08ac882b5b079e81f5ff34408e4d7ec516c2622afcf48a4b4e2c0ea3d3365749814eb9dd723cbe8b350f7c9516c5a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ce47ba0d64ad3f771d618131af9b536c422134a467d12e70a216d1ec24f5cb2a02f3ad6281cbfdcc6910ac785e07a455e37efd15ed34a6b37a53cb88b773375ecf809f2ad172e512005ac8246923977f3a33c1eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he64069f3ac72ccdd96f75063db113a308444060fbd098c395a51c284aeb0df8a51faa6248dbe9680e6f88b4dcdead61c9968e8fa42f02f1ef1410872c832bd2ccbd62972b0b7ff115571057589a340451b88b7dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40b6901671276c2dfd0d79268bf997c87a077fb7d843ab24d09d0ad012288fb32ac8a21a51d498897243b1a1cd1e5045f09f4718845bad74d872b0fad6b879c18f93260c135f05f0584627ae851f8606490a2b731;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88471f20d24f872cea76dd0261ece4a841f00e033d0bca74b3dc2d2c58cae5c65dd2a7cec63b49c01687f700f24ed2978b0d83446766a0f7d9d8c28d8109cf9423d3eeaeaf06c402fa67e5917bb7d485ef54c9839;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdd19863ebbe17e06fadac7acc353f2e520c22fe1c7d09b6dd7ec56e35bdc843c509140d145e7df0cbe7ff7491d346ea4eb6b3b7fc4842dfbd378114d7a6b9bdb15489c6d330af97878c5d0645f2473cd098b503e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1efb7d7d4ba8cbea06fd803ec446eb4c832884ba4b1bcbda4f49db894931b17c14d375a9c0738bb51f0e81a11b475b28515ed0755542d231c4ec4ef718848802052af7e119dc35d40079eeedbe3752c6e4595ee1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d0efab8210dee754b7ac79f77a34c227ae7e66811a9074b31641997082e0c1fb57b391eb891caac89fbd153d1b259647332bf002f11e965c73228427fc74ba2c6e8e11707b17856a1bf7a490c59e969f88497b8d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b23ee8708359d129fe5bbd2dff7e21cfe66e26b438948abb4dbffc612bc630fc786372bc80f24e2c494e2bc078b0bc59d90a8faa1dd7bc4f25a5e80f55e8df258196afce17dbc149d04ee39291e92d803f314ad0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff8f401cf1951aafec82a4319b788c5cc27bcdc541f62ae99c9af80a9b1acf05a581ea2dffdf8fccc3ae178e8cea61cc12edd76627aa8a72bcad83ecd0c9058beb8c2cb3229b03a831d00eabb4692a88d654932bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52d9c756ddb808992e094a445d167870dfbf06a83ebf3a7dae8a1964bf7155e79f4d7c15f5094cb9ed42e48c6b57cdd792c9d2169e41a33c48d1438e94a1d254e322cfc904ac0d737140d451d67cfd0162c19d709;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf63122d002d3467eefb8c7dcc59dd480b5c71e9e73aac324beb2543bdcb588075e85aff94a9f963f1c729b3ef405c601913e635f14e627689a798d568925a24244fbe96c1b595c46cfa46efa5ecdd2f551b450982;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc55bb77e445188943ee1f183f8137cb3f5a45d410833ebbdfe4a765951a43e1c894bed8c0b011576caead58707c0d2479c2b0fe68db3c3a326cade203d38dae836fa1acb44899e63168927ece1b245db35eda582f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h520b75499e421ae0ce98d8b22f36cc4aa5cbc0ba4b396f175fcde61a9a85b7b8681fe4d7c6bce1a6d7d556e7da60c74eaea270bd85d65ca2c9e28fac8c9203c5a552e9c7a25597ac9889f293a25df3912fc0b38c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5071a5008bcd08845654ef6047dc14634a09a0593bf94820d8ece5df573c069b225e9f7e94aedf6a62089fcf8eeba8aa2d183e4950fe96cdd9286112ba128f46ae96819feffabd924555fbe54670ec2dbdb7a1f23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb1807ba566403b01651768a1324983255f4698ad2af11455c0047d421abf93f3c6047c61c9fa6f77a8b40beda914cfaf4bd26d574c0fbba495a94614ec6cceb78fd38778995b363171c78b4372b0f5dbcbb55e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8efdbec45f93ea43c1f510bc23bd3b0dced523e5725b13ef04c24f988040a65594e39330099484ec1854a9fcbcc855542cbe004f1c70681abd31d3d54684be142b7f45f34a660a4ef5645a6fc71ac834f5a95149;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c64b385fe724b018bcadc89b7b882dcf4172c0b3568c34934521b1a3a0af4af1ec3f3c4ff8b0809081bcfa7cf1d1f50454cc67182f14dbea5898049ad7719bf86becf6117a7f81afaac3a80e876c596c73bb86f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha044bb5424a76b4efd8fe63d475c0415a6d5e4baa689ab4a9f3f1ec01685ac55dd8bcedec1ca9b290cc34c3214ac890a00cd6d9be396aba311660cc065de999cd995f76a7d4eb1c01ba6162b058606bd9fef43fd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcacaeb6845b5fe4156f823b8a5b9a0ffc915917ba499b6e72876fc466cfb7791e4e96796cb2993aa705dedd06b98277e17829a6155458b666cd9831ad934f7a55bd5aee30d41dfd94717b77b180560a53fd2fc0b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf154c1d09616d1a9e13709604f4c23b25d86bf5776aaa25a4c1cd47e4ecf1143816ca5f4eb163d04c6f32b01cb03cafb5ef3e146c10369945123c246d23edc75c1eb7591f655b7a14e80de80f66e1f245544a25c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h148b8d63314e7081405248a99ffa7ea61c68ed138c9efd2b122b1ae63389c1d0a64a2ffd0e17190388fdf3a97e12da009cce1fe1edde16265ec8857a3d8da7cf5dc02515f902f4fc1be1db874eb8ff50a62278fe1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h449657cff16af9460ebce9ed944d08a86a4d1741e3261ed7d89e22ea0dc19727462d88d59ac16dd6dff3cfc85aef8fc6248c25bded3363ee038aa9df7ea6e11d063f6cec6e5b390ad9a95bd99fd570918f6cfc363;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6f02b028d549f1d0f012fdbdb01aa53d735358b613a51a541bcf2ecdbfa9f7a7294aa7a78e1268704868e014a8de0e07ce0633675ac0becfcbc4f9933f869a94621e5f7a96f75d765f190e02aa263bb5b2fd4af4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf781b5698bd4b9690dc89e9da93b1fbbc0fecbb29d91b1afe3ef5f0627883edb7142876a2c91c43d1f28b287954b970cffcd15344ffb4dc78fbe8526f0524897766085f47b8704c5eff70de0149d04b1fb249a1d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ca6a10d306d8f0ea74c8dbfefc0faffe84328b330be2aacc39d74a737a2c374b3560ff42215e91938b84344f9dce9d4f5ff11b6e55c42a82b33ce5c931ad9d4d6c26194abe4aae2c011ef3e8afc1fe7f61474e1e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bfb645aa5c4ea2360e5bf4cdf5ef412b65d480ba4b02cf67070fc710624cd2ec5af39856a6e579be55f0ac02922e5543a0488a2f273ae4c84d50442596cff2ba3f1b5ae6a82362a2e6d5e9300c7d3f7e489cac4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf37851a73ac7a9f850dfb726ee4d8d9bc4ca9cd3aafd9bfef83069afa978a529b1ba92f0bc8ab7dd23a220ca5dd90a3a76836d0a45cd808e9743fbaac0599d8299ceef41bc73ffc470d1e57e9f53558044515669;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78c13149371cb7be37e93d9310e1e2de04f2fd063a09937aadf18f39c8b59d0d6f31d17f5b50b75d7210dab0053ab506ab104be782d1c961b5fe5106ff51f47f17698fb53f2342a439e5e40213ee80c9cc283f61a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1192012cdbde801873f0861f9a045ffc2c4da43f2241e3040a4c2c7fc433530c762cf5b06ee3f54aac5b960e33ec9f6b8ab589a988c966244677f3be056c73f9bb510d1cd18e28a874a2af548a67440feefcf06d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8553cfff31d17d75ab85f8c1423d1da9d5bd450d567f30798fcba9103f1fee5cbd9d378352a886548835273f27ebac841fd66acfd87ae3068ea5ba1ebdf607cfc1707e5c5f73abccf31520cf76f08212aee03fcd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63618080486ec195ab37f39a9f8a7c79858210c225e866ac80082c274fd4791c27742ddb96a44d17c99d1d1406918ba61f780a2d2a460e0ec597379d1977c9673b01bc1e21d0581662f01c0f081591d0648a7df0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea94816a0cf201408fe42a8a3303aaed7d017d45e55115dded944a0f589dcc4cbdd8c7d148e69980a7ebf2181e10b1f7a489734ca71e646055733d6a3c25e33a3f792a9b262cfd7ebeea48f0ca851ac8769ae32fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha86a0f1abc751d52493b48b561ca48026cc329e26b03bbeb8ab2f99e7530fa234c07c03cd0c4339367653f8d7d38e5b9f4e6cc3a71396d9fa641133c733f9263945e595648c3da9580206317df84fb0494dcc9c0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d09c24a0c9308c9f3565e54c932207a024b946fdaa1e5511dd41e913f8e72073353258c2b211375beca476f81f37060385a264fc4f4951cc0b59469cbfc80e9750301b7845c69472edf533e01cb81177ff488b34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5d2b74a88a9c971dfd7b2048e1778e9acbcaed6a9818bfc256383058bdeb865e57030328733006d250bbe5483f9c4916022760146d9dbca1cc575544adb004f6b674aeb7158fe810d230c12e131228885523c760;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8edbc43b2120a448d939538d19bdda337a688157e58895394af532376857f32a26acfb52059a1f1af3b2df2aee45f0d932ed42b5afa46ffad8fae5bca0616a4b514435090c3b04fcfaa7bf4d7432cd7ec14f2c20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43fb950ef7b09b61bb512e6131aaa6d4534a9324628ad36a8afab75b4b9893cd3215419aa0a46512c114478aec131de920165c042bf588da458eb2a6f4a2e35b0fc83d0814d3666a90fbe8a79ea5d4a50dbbe79ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98712ecd5c91c15802b2621495fee40693635c7be6c11c5b02aee1dcde18276da5e2a05eef859c476e5ae8b5bdfdd870a65936ae973adb86decd969612e09236325f9a90d555526d49cfcad6fe7dc0c75a058528d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha08efa8b546fae5db8693fbbd8306400d0a87bb9f030c4cb865cde7164de2cd06813c49dfa1fa7586bc1fc626357d32f12b675eb3e1d8eaa87240b3448b6821d6989184942901e907dc01c0365052af3f8e90d193;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82e606dbb67994a681821625d1fdf7fc4dfcc74d425c975f5c6c931c170e41b9303f2eb52baef4a03e5c69c1ecd9afc0209a6f015422e64a1a3260403487ce3c96c56570af7e86503ed77cc4558f06a7844c01343;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd17c706990936abaaebd0cde04b36233e15ed63ef0b677df6186b14cb67f8d074806e3f7d06be561423c847c0204caed69e8dc304947739d65834a1896477d664ca720dcf3d629b6a5e1b66a99bc5deadd2a23e31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56cb7fb5e15889692f0a244c3294a76a6b74632f125bfc4c5a14146186c8943c607b290a5e32770607802caea790f4309f08a801dac3e81c8e42e067e0d4e4157c02eee64ab30b49f3f60d75ae7a9e04d020c52d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42463bf704df47ad1420ac0bb24b27dfb6f90c3b80fb6d17954afb050caedc909941dd6f6f7e3ad51615c633e283305138a1437125ef3fa30fb8844c9f6395bcc64c0cc183f73b963d3cc864e055f233ad3b322eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3d5790527c6824595e7dcde18dd35eb4521167f7ce7c8fda6da15b50d0475fbce5e19587559e1856dfc5cec0d152818984ee22c57c8237d7a80c736301f5ae92a90d73e8d4b38a75ee3c67b92342029a65f98859;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94565faae85c96d723043be476c4308de2c3b125daab03ab8cedb61264510de827dbb57d1396c4a40577d529e4797a164d22d31d5725a1f6c001f5008b4a176caae9fb0ac55db514c62c3d977e9081809d260fa41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdb23ec5543fbde4c4add57d53d4e5c0305ed14202248466cd6af27c93741380d9f9a1fab2b06ee7ec817ea4ff7bc72f6e7c5f89f6ec25af81756b39e3bd3805bf59edd5f30a042fd8947201ada77bbfc120162b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10b62565d19fe6d8822e7ba754b9a2fe5d21a1ff3603a335d28998fba851769cc30a2afae97da758dd6f1dc3e9bd3e3a2a7906a9a7517e4ac3b78a54ba0a55769f8fa29529c5c7e2e108832eabc24aacb3696ece1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ba880699a01c8382b9da8269f91626ff2a59a9136c2dd8cc4b5b33e92b82864dd39e627399467c8bcc1fba228feded97b6fdc57abfc4432da21a054320b8a28fcfe79d5df41c4a692ed16c8519af8722c75d3e92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d78091b034d192514219951aca1abeecc0eaec623023227ecbdba038d9a6ef3dda8091112f5eb712487ff3cb8e47f7c95d144308b6611eed1d32f7a5ab208d008cf00e9a7078e40872d25732381a0facb94ebfe7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74062420e782dd5938444263f60306ea3f3a3c39986a35c0c7c1e0c156fa8e0a1fd5b2e7a678d35cc5e54b2a7414a2c754320371df86293381b07aae7f2073c05759219944ba83ea96cdb7ac2485a7bb82a5172ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h320c144160c7e4903e3e0fd60c72957a27585e255eda61cfb4c22b1978bbab0fd508146a3770c66922c9688da04bfd321d6024470d9936f709f1b1de45735119421b3c479c5586838be6a0656dec98dfffb3a1aea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcfab0a56c20e18b99c6bf7c65ed625033501cf15481ed0d7533e2a1eed1471780422beac8ff37ff8c44e62f265e7f4bca732b0b625b26fe0464d8af3caa08f48fc9640f1442d656bb18f763a2bc391384336b0ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf907c9dc679d7f04c0dc010535b81a8b8efd4c548eb1d4a8bf83a1548772b29e52a80e0f38fce2f71935c73cf06ad84b9bd946c85bed8f53228ae174bfc78bf70f69ec37eee0969345920a1e27174200d8e976827;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6d9d3247a346363a5bef01969aaaacb99033e9680e6e86ccc63dbe71db0c63e5f4423f47e0a8a963852667f58c5fac58c519acacf52ba07ba268aa424e621a58cfd6c55641b6b40aef0fdc93e1abc1fc42df2ec0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bc0787b2812212a977bec03fba9dde936a5e74c3744a51e31fae4174da7ebf431afb8425d1fd61517f0ce27530bb78c064c8c23e7d6f19d5bd0da099c9481d19f7f4dd5bae8478a02eb42ff7a35a0ea4bad033fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9c63456333914e59f3e3685c76220ecbb3d9f2c410b4dd1ab5a7bf7fb455cf94886d53fd45256f4b52568e8623636eab3a7fac2c4b78902f5ee800cdfbcc90ff7cb02c21e7201b5848d8a7901ee0acc998bcc64e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc950ec306e7c317dc3a0a98b99956155dd8eab31884baefe021f8b180afacdb0a48de32e301f574f8e3f05684fa94cc27111cb463502b622a4fbf0cf9ce2dc5ed48e3ec6f4f6623a0e95cdbaefe19b87835e5c97e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b33e448743936c044ff790ad80a4f0638d9ccf434dfdaffa3e12cbfe6b63b223510b2a9ed2817fac281c29578b92a53724822b3f2c4036ccf50148d140bd6f1ff4a908b30ec631951f448158c736ae511baa7aa4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0e8d46c1b49f227e8def3b04fbf128ec9b2ec1bbd7010a1fdf5e9cae5c1d1aede4af83accffd4ad97bb6d9ce7ecb56352ca9d0522465633981abef032c2d5b4c1353bf5a851464f34a0de01d346ff165d1531453;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5fd23bf4205063d40bdd27de263971410dacf2afe281611101dcc71d8b5c28cb185829b4b48913e83df8999df66c80e112fd6bda75342307847182077de358ea43d796f7de2acccfd796f5fc61468e167ade0f92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ec2e94ae9cf2d8da2d9496bd1b8c427a89c5bc826fadd3bbabb577c1dd1b5d65fba26f98e3ad9d86c32d4d49e5a942704788d97dc9570b5bf59cede565858375207586ae0f654e3af2bf34b525da237117da0d86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha342e673dd573e379ae9ce76982fc32ceb1c1904dc813b3eeef32063a3db82ae4f8e4e6650fc27ca5d555e11741d2cece3a8c5a5bacc2f5c5ecfcf008ff39a8b4e2e2f12b30959ef3c6c023a013ad0f5e57e02802;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6193e5d37fd7d2df348cefcf6433d54ba2d4f91408f8ef15ce7dfdf8df4c54fe95862fda75735af9446632903780618316b287f39e8ac5a4d4320c7b0d38d181c8695adfdf3bc3fd26dd9b80d85ebde64fa005e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h278c9016f823340fcfd6220f294091c9a15c5804bd7a88f9a0070eef922b9651348c4e7d8e08ca23eb0aca645413aa71307d785ea98e9f6b4c19780933e8a46acf4bec79b5365e513736f606a76a5b2390061f1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha58c949ca1ef9d7da1002dbf522979d8e7b631c5ed6edda573bfa0c58c4b511eb34c5564f39074085c5c2d66e1069da43d23e685f33d9ff09f3b102e769a330be935fbf602877cf748a38df3051d6dba0355bbf69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6da0806389c755765bbbbc4a899495dc9babf19555cc12dbbd9c6f001c135982a70a52b245d3d9f6e7af1a3d8ae5c8975d42689bd8ee93930393e5d15ae0f1520a5a60375d0f96ea2c4c555d1784ad0d1ef5e232;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2787d94086b825d986800bc5b873bd4a6558cc676b21e3ab6c7791a1dc2ed22e49b86de458564b08541612f03db6b8165757211c8646e7f64fc5823f901e6e571ae4fa0fc3a4698d7696d56552229edef608cd6b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5debe241f2696dc514a6613494d13a4cf6afdacbb1f93a18b421960ba35fa0c0df91c6ff896b8af56fa812a27d797ceb15cffbce57dc134e69abcb8022fcc18913c5f22caab3a5ac3ed29a79701dc1d4bdb11eb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ff6315e3e18c8b8aae4465efb346ea9e2f83b802d25937f85c83b42b4fdb29f0bd4891f7a8ae599e21c2f7791fdaea84f305bd302b672a53fe38c392f46ffb754342dd61fb1602330f9c5df4f1c7dd3ecf8f43dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99a1dffd064d85b0febe1e4f1552b6fb7add741b9e666288dfd45646e9f78be10e30bbebf641e6dd5b0d2e6a1b39554ae3d48ed47b3a54c45597ed12fc9a6907c6b0f67d03642dda2a3cfe6d725e74eae82fe28c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33f8b06bd4739dd936038c45d1ae918f17cf30c48ce9f41b81e0a1a9a61ed84a3673f2e705e7f756aa36f8240e25bb711a871d8a4c1237e65cebc91cd4636ad94258f1ab4e8ebb37010b5e20c2cf5318a61bc7b86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e46a0f18d9981268f66b9914313298c80b7a77508185dbb3c87a1a3c39c4f6cfe37bd74c2ddce841ef0e32d43f9f6af4d6a94d0d77a825b13a1d82cce50ddd948c41980e20b67811af8b7e349a2dcc2258660524;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11f7a3dd6a2893c1f6698c5f60be17b095182fb2fe4efa3712828f06c8374698cb87a2f394ddec80e21a0387ccc6cfc0d5a958d09017911b22d6c9d6d1d5b3c83dc5439fecb67f6c620c3afea669d66097ae2aa38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69cdef1819af2d97bfc837cf07c36ba9fba1e58d597c8c7aae51421cf4099ec07815a33e6b5f933ae17afcf38cd0e80c9c5bd17d1978f0dc8ffb6c7f60d083f793a112dc4d7b281461eb6b90c76cb72fbfab80811;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16242dc9e4285fbca68e84714936b0a8caed1aac2d242678e10973a8b837ae3c789fbe6c0d6888357a105a29b16ae0751aa54099affa3a28de75c331795c5408016e70c513e9db7b6483b72b46f0660c0941970ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7668a8aa0f3154b3e6d1419a264d7ee0f33db6fcbd2ca2df43279309ea0c5b1f34df952cc07037613b47c4f8c2b25846e0944d869e3099c8829f32935efde69f6fb69a5965ef776abbca1cb9c9b2cb5a47456dd8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha32f620493813dabae1b800d13495b8e56087b0c0a31fa0600838e53d08b42e1ba21ac385c6054266163999387f732079a065a83fde38ad66edb152f51ac68298228d2697d35212b6d7aa89d8a9487151533c6aa9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4e9ed43524febce9446adbeb1d1d0671c26d031a42c6e43801962b5dea97e600036b307a7f5efd65156849d13fb696907a440c497356ce1b219726800df26995681f197700ce53fbb2678246f6011cbd4e6e8370;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h117eead617619010dd41a958b8ccf22862a55fb07c0c5613f3780abfd0ac46310e213e42a9e60ca756a1e75aee92d4786211c5a4a287fd7a52e3138120bd815bb09abcc94d6de15b5b52f4326df259bb02e31fa12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fcb5c8b6e1c8b5c8def65cdfc64c3aa46cb030057924cf5868f65d0d82de6f4ba6c4655b318f3eec34f1e7e4c64c9fc603c9149301226cc72050f4a0dfd4118c11799a65900a96e987b3dbd82e9d361fb8599073;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ca0ba239e92a62fc047ff98ae52a812f2f62f8458c957b7dc691c8aed3fe2e88f9a8c06d58c4e2a6d5a60b87781fb2c98e45b4db3e4398633775a1ce615b4a0514fc333b42a98f83630de529243623cb2a681e7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h485d4cd4a1ad145d8c23ab9a667390c3d0defdd79d6ea7d9890eba82dd7fb482e1054e2d484b0ee9eaf38449c94b6df05a1ecd65dddc18d499aeb61d429a540f5d53dfa5ebcd22cdc4e084e6797c8fc2aa71d98a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71022f9172570c755bd925c83fb933e402ea949796412f01fc7733f5d9d239b3b52a4ca77fb8195cc4e9b5e4cea4a0310d1b84c3ffc5ff681b04b120f902d23e0453cc04f0384a5f1c0c770a3e19abc411a2a27ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3623be8cb873a72b205b040b5bb2edb54d63277eb376283318d804f478441301d79ab54b316f8642747919577675fc74207737445eb96784a501df7bbab90f34049ff44b43ca44db8330729556eb3e5a753de941d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f6f15cd705005413d0ca9f2f19530b82e894bed31696642da6860ba319bbe970dfa08b18255b3d8ec3b9c02e5ea62eceb636d087c43d992eaf7ceccc19e18b6f83afd39658fa0775ea21e4456ae19122bb70da69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9d6bffb73c8a36467b2510e9bdd255dac69485124a25f9f13f49a5fbc8c88d82a0e9bac1e329145098ae33bbda2365489999ab6bc600af4ed2790b7c11ceaf2276a042afb01a5b4e80e2e45058b76cb3ee7189dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h235b23f61cd8cf600a222ff4b2e9113a8e3af218e4ed68773359e5c0624137f007c359223ec6029dedce7b3b7a8496347705cec8b05f8554e8016abf93b445c999c217a6d6e09ac776844b5b9c67b868115a795e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e654389d1b219cba8d2d83f0bc9998523608d2d3fe51c37fe30cfb8320b76df69d074ccfe85dec37279b4170d2760caf43eb316b4fb37e4e3c02148b8dc1f78085a09323c29a683cc2407e96816fdedffaf1d982;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2438f8b0607764600e5d6bc6cdefaf9ecd78988b9b7a2b35efd0737632cfc85c97bb29b9bfc32b0c1a954f5216b023d81c84438611be31a435197a44bb7eec637b0154177f1ca8dcfe75bc9e38a3c65b9c5457e99;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h302f565bf12dd5d42969f7fa7215f797f73b0db0abc5cd079f4b583c41f1e27f3dc636dd052d6e6789a7522a5473936c0bcd081148882814bb9911a32d595e9535d469d798e2050b193a3bd916483a7b6acfc4281;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5ebdc60a91bb6859bb4f48aee2741704e1ab9f9cbe505480bfc7298036e69e0c5eb25f3c48f9639d2ffac27e557667d2a7c9a48f9c3c45585f61290df99188fab99853396bca5b8a007e168018e16bf647252f45;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a6ce7d58c2e68e714dab660f2f5ad9d644583774e2fd273fa77e3820986bcc3e551e29046131ce6a7bd8f6c1d07d4a35e9e087a4b7828bc1ef6a5d763d93d9b44dda455fd10bf16e9fd48439440fb54d85648762;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6403e85784cd114f9dcdd653264c8f1c685d12581d6719f521c1c4a471117063f6ece1f3d42ad6cea1bf31df6d24717eddde1fa71b152809aba8f9ab98c7ecca8d4e94f8b3b1fc278c6f02f9b1bd26ca3709739b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9eb199f0c0d6db50a909bacd190ef35443437907f3a6003b1d68914b23dec0afa135158bf01761a0ff067054cedac559a8fef16e655a37754f3347ceb5ba1f682709f1653c546763b53c018e5aad83c577f6783c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafca29f9baf654c954bf39ecf3ee3139d248222db61e2c449ba2616893d5bbf1aab44933e25977bde0ace378b9f9e977b81327a887ecb3d011dce6c2baf7adb775e76c7a16861ef2ea75b10a6d69eb52a686e12ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4e328f090efe0196f2fd97635c08e4902374a957308ae42f8f77285d07a898aa7b1af3870b41fa81e45fd7a283202a632f3bdbbafa2be85dce138c7afb7a980d509f4ee4eda4d4fe5735a39cc8501c2b96d5f911;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc648ae06f62a429bc01fa36bfc147b5f0316d6c4cca15c340aa1016a0ac31e08e90c8d2ff2e451284ae234a9fcbe5452899c698df66015a516985c5187d69bb92a34ecda46c88db12600c6f1c8ef6641c4ad8f70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68d474b83eb87b65cf53bb1405392ceed94c80c2e4bd00e851e0b5f1636f94fe966658b23754b4ab7b14d1386086be522bb083ceb054214405e7e10a1c799533f084b76df0c295db4215ab0f6eff9952efdeb1d3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff553a7c52df63f15ce36de0a5fe2f9444d89b073bcdfefd80b6a8d813ebc6a19264b536060a6bb871cfe56391656fe82a4ee72feccd65cd0c0643a5f2363e12e608033d27741c823dc286e5852210441a3a35f38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91c3c629ce789ce1d251747e48931de5e99fbef77f21c332b817f64b05edaf7094665e8352f876b5c4ace962af92db8d42a775c0f30e49939b20f7de1c491b8505839da1751ec232b72970ae88746060b2b5cd12c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5ea0f0600f795993c905e4c2e4db04cb7d93dbff1e3484e8ba28c03405dc92ed76176fdb3909bbb87c797475d434ad5f593258f8ef9a2d04535e572f74c0f6d6eecb7a6e040a195684bc4e3d1c1a5cb015d4c374;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb74344fb84f59f0d68ce3185cc161db157dd606e1bae07c148abc541e61e31c271b0c2d5f0dd8fbca028fe31d50d4a98c9c35191a7b7daa90479e7a135a0b3dde958bbecc6bb34bc6df17f08372326e7f14c72489;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha047e7ae195caf066e3f5fb0051a92f52773613c3d7ea955cdc4ce37e604246ae02ceccfd65d1ae94d76dd1bd2794edfba556092bf99f226fac6dbf29111184eaf0f64aaadf19e8b66b42d64d2c33673ce5b98e57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a5945a45584f8c1a46e1309d643bbbc13b6f6c18f2d035bab21e2ed88b6454bdb6da32c547f1c7595e616a9dcad30032fb3eb1402d8591cbdc675a985e70407db671d9ad2e527d7fe5dd5b0f9096589651d5fee4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab45fae13614fd7a2b9eb15f0b3ab5b891d0167da64abb869eb6288c7fb42c8e1c842bf90e82af5cae8bb842664b1829aee2bb51d6d9ec3754a10415926cbea2cd3d988a38cdbc1b200227b4f497cd8e619684b06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf62ce23fc5ad31c7d8efad76b6549f5455e2eacc46cd1738b0a1b09cfdf80dc60e4e06085393e8e4f4486e5bf9878dae0ee9ad3cbfb991b992dde92d105dbc393ce2096799b197b62c40be5fcff122b23a62bc4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12c7d0d8d650534aa26065f6598e4236b8ad0b4b2ddb9603dfcdf7466a473e0325c754811a30e5876364f320ed6ec0575a1ed04aa41c6a0dce23dda801a84713f0ccff86371ffcad9b0369afe96c5735290659f15;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7801379fc0a92a8d63efd6ab8b6acd097e2dcd2931a2f5aebbae6817cee3ac38af2d55b8d84a26a2ac6fe1a25368130da3ef41844203c43b2e469ffeb7b7bb8ed8ce8da90895ad21902504ec0742973fc163ae430;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4378dab19715cafc7610038820e2a8570afd02fdfcc4452b71b084cda039bc0054bb2b796d77d6965f1cbe9e9b9577cbc2b9d1ccfe094a95a75a124e2c153c0b72641cbe33dec1c5e1b404984984f98f8a8517df9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb622397e56e31d78ac54aa3ea0d85368ee9413380f21a724f9c53eabe06fa1fa6ca1399acda7d0b677ff769781307139aaebf55b159181f39bca4238b4f3c20ee32a5f24dee7289d453bb0562d97b4bf30042802f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b126a456897459f7204056031c95d6c15806fd268176fdf79d1c4aefb9d4c196daefee8b48e9c9104187c9d2e52638e327f2acb9bae9dee3808cfaa40839d8624ed84d79b8df63b44bbd7a5b0ba177d4a1ddf05b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1ba1e283c63453821c9df9b8858a892d194c932e75ce16e8ef2238a50b10a59989c1211edbf17f012d80997d207b86f2c9ef1d8bd22d3906c2b9f13d5f295cce4c26640de81940e1764eb13d31d865fdf0abd03b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84309c82e5adefcf19625753ec5441afc587ef9d327582af3c8b3dbd30241abc35d022cf571529021b23f323e0ffdbfb6a227727035faac7de8d61fae1094ad97dfa6d05d455f134759d23281cc9febe1dda69b81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h251cb9e817b7d502aa0fe323c457ead70c6194c08ceb4b9aed1a2a6d65fc18004e9c4ac7c59ae96e0a8091a95321bbc1315064ecde8271b56c4d9ff3571e768bcb31e6ca47565d32ddca7275c927161b0ee80c51d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2a23ebd56ab7b38d2dc2096f4e93c9f3470a8cec29458c869263c9d02624e167b98a845123427585e25e4084b11aa545f658b6a3b83214562d079fca4e0152973198a0b1d51f891e95747baeec61b0be7957ef01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h161c4262b07632f4258efd248999fb157b817e530167ecb2994a052c2379d4624f0eb81f8f7f99dcc243de85d1abe6bc53a10f0bd00bad8a41fd0fcc35dae6b413086097f62654f9347de0cad9715586bcc662dff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfecccfb9f56e8703e423187e76e612142b7143d0b894b7e1cb289b03dc8e480949b4fc659f352429469810456eb7566cba1d90446ca23bf9b4133f3292cdba24a5dd4c53ecb4c9bb6a490c22ee8a6a10d2e736dbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4f35e8b54f8c06f947020d3f54906233ea6a7769cb29fc58729434c3c4b82ba09fbc28b57546f9ef40b0e97e13b75721bd0c7b739519145e7e5131a7c2daef8e7144e91cea66089650fcbe287d622352a486d60a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he52562fa1e16028fe87d69791e59934b53cd5fa327e82e7468f5a300a4761b23e981bb783141b181f323d4ad238c7d3766f72420bf7ece6988408f290fd6979ce15c0b72c8df7e659473248fb2a9c0843034a8c25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he18f6e2f8f38e6ab6dc14247b626c04d9a07112a6168498f09a1cefba52d478a7517ed2ec4483ccec6cc1a583edfa289594e26cd761ddf9191d163aea2b77555e27e818a5edef09d865bcf01ecd09290ccc77b171;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf64008943d6090e59ff92a5ca9d2a1a94d1d57f02e5440488343b50ab7e15751ac8143f785f1809c70413b214f108b754a873e80cb5c2413ecd2b0311a00d8e70fb37f7b50950e05e68cf360859f80bbef13b186e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d087ac6f0107e4e24da31e90a3f10ae7a019538bf508179272cd9640d61b2abdbf0f129533258da8b7499ec285451d2675e8406859527f871f085ffe1bb7c44e895e47809a240bb0685fdc307af3306bbf7943fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf71182396df2538ecf3d757cf506619ecc0334d0113530b4290e25493e94650cac5dca0e14986d5cb40eb93f09ea886adf20327bd734dfd117a2990f924906d21d7dd30fc004eb2904ba17ce28d90d74d90dc6f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4426665146b0791ce199e51b6a93b434ff5b7798a6606e17edafdfcd6d80613544ae30b3da387fc86961f5b0daebc6ea9ad214a8c3f348cbcc0080dacc3ae35c5bf7c5ec3d8e9529c7e59bd1c23b073b76af93fa9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59d2a23a6f4fe1bff37211f9da4b841680c59f37ed1e7dd2847f52c4d3976a27ff745eff11fd31656326a931554c77dc572c0bbcda4de58aa28e75e701cda0b3558f23320641a3aa277bc21cc9d3609479ae3633;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h759fc21428f59b0133c74ad70f7f841ab35e2ed6c1c8056f2a7163a39af1b4a62cccb1ed7717597263eec8079058b625add71569f3a832ce8062eea06c5fc76a4140d041075504afe4f7cfcdf98e0dcb9872add44;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h531c6338e1d12605c9d87847b2606f254f7a83dffd138537091b65b8cb2e00c431f50cbf3e75361994d713a23ea3041c4daf1894911b225aaa1cab8bb767e60f7e19468a82debce17e4c3417caacb12c79acab666;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e9546a0cbe7147040a122eab736900304fb42193a6494cac92398c193a16608b469c0c53741a78046e4664c8dd37805f412905474bcc5f3ac3a81bc8fb9bbafb0b97d83a6d16d2e1c617d5c1900167965ab41d46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95ed71c8594f3a9d2599e20af3b9178246e06c6d9f7859e641c2af2a4328498189bcae2748e11fa61eece6b6bbed5b1742b55732cb9c312aa78220da843faddf15c3175424546ff5de3e65b25bb588b49fee30fc4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h684d1e952b33dc062068075a40d9e1360fc8f5577d87074f035d5b81de12e35b87a88822c062e205e27ea60147ff3683412749741498f41b8aac2cb58879d6f9e8a5f34f5ab8eaeeca498ea5086ae80663e16f541;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaed2e57eb2f3bdbbd218a207143c1fe689a38a4268a3d602209bf8d73d16cf8dafe24b6970c4df556a42f6c94fd0d7d89ecbec77174ca88301849f784b8241aae9fef774208c53f96607a816de64334a427319f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb1c5a122c14b33c47c2f17b071592bce3355cd75dc834824d49b18c626acd6deb19041e8045a69ab4912a13c37d92361ee97fa9876945c559c5f49a63fa8eeaa29e1ed6118d58bac65277d5529289931957a71e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd92a66513ae6612cf3f258575f43dbced0ef2809a10764355ee46a33d9d5f8df25d4dfc06741ca5933f3c6778f64c84f0e6d660dc034eba7a05a3343ede1a13cd04eb156151fe6c7b1958fb125a377f52ac0d2a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h817381c92ff408b588c97806e20085570fe29a3683a611101dcd628634e27e8b07d82c0157b2fb609b6cd18e8c6662f0ca5abc190a803eaa040a653d1e75e9977eae4e106e1ba74a99f4d34039ad9216ce7aba3af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaec0d6b96d8d725024982a34b4e49a6e113c53208c5914194696bd8ba636a04fcd3c37508f314fc6a51b52295a500a61655b9f800404d1d5c170b6c4d6fae73edf2d484b07b4a2ac142c2114030c60d80042e22e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e785e794c6eccd91265def900edb124e8a4ad7be003dedb6ebf2933d1c49b1c5b86295ed31479a9997b05d66570f330a6f1e951d755cc3ac6368fe3b81faa4825e6633f33130c1792883d0408d07a0b32425dd1e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b0e91bfef012094922b745a15c77960d52b249667e9ee9d9d91c8afeb6b59e59cbc5d4b1cb1891be73adf6790acf18e8c3868bf816fc9fe089f0a592642b3638cf6435cf8ee69bd007ec4a087d507a80fbe88e39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78c9a06154e9f259b0630b455c8d35b3bc55b64bf27a3a8eb1cae2515fbbfa58632321b84b6458da2d628665e6880fca9388d2031cc98d827cf573d5d787d53c8abf05626baaf5b03c5ed8532fc24596b4171f993;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h377b46611e7ba2aa9855ba88ccb2bf6674ebfc90186124a2f10e764481435b1d47169a43ce2f7749c226218c5324ab56f36421a86e5de05ffc2291deb0362845de9757cfe77fb5da9df212b9f249be7270b141394;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62d664d2a079aca116db81b5dd0394cbd827863dddc0dc86e0274b3d89fdcb53f0957ecf2de59da543aeb73a522c90fc0e8371dbef9e9a00b56e7231c71e44ed6a2f0cdb983c5293794ecd993e77ab7eafa19843a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h886c30ccfab9584723b62302aa218bdfd7bcf6ed832aceaf6bc45e324c9795074d031133877bd1309ac5fb222a614a08f112dbb25b7f0003cb14901ce28048293170f201112741173bb2e4eccf7ccbe050c316ac3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58216e36e82461017b66813298d1ce41a749fd5f17bf5ab673ffc62b862ccf17eda664f82b83bd42f53c53d49237192e675fd46b44d396cfc6f331dcc602fafded56a3a7ba50a2cc17e09d4914076056190e1df5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6c8ec0a6691bb49d6b6c0c8598817dfc84972eca399d03cb69f21f6973aca50410c726de381c61b03ce01eb18e1a01d1a58dbb76c09714b4a5117a660f7f7f26e2330d3febc39d56141caa27918d06cd0d66ff2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd795c3cfa4b1fc09739cea466cd6e62c3c11f1443ea5141ba32363e84771e314eb765cc8e2dbf95c8f6f242b45aad5efcce4bdd6c9402709bcb846e97d6b0ba8650cb1b34015be28ad23e3799aa13093a780e9814;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h488a548b1ccda32134ce48c837f2c1727f2cb4cc0cc8d9c2c75899e413d19a0d6929335429e528011ec66d18586c5cda0563fbbb0062fdf7554342a57868f2bb2945e1f8f592de9bfc0ff1bc6af78bdb4f2edf95f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde5edde7c27e3cf8d5a71f581e14f3643bc521841a5db22ba88700d7454b5137d7615ec32be85d97f695456d631e0f17429054a57ad4d6ba07c5ddccd9e8b9702998bce570c8dee298c479c38f6f61ee5657d9bb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca4272e7c82706bbf4911aaa1b7dc76f8c5d0284da8fad27e7f53b356f9f1465de2430510547bb12ce2bb5976fa4f287bc40353666a2a070e8e917b0af3f7932e401d17d34666646b4dbb46684f636a2fae98f627;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h698d58d20242c7c2260864e88bbcd3ac65c99a7fa98f4ecbfa86e873bb188c458e29364fd5defb50400a72503fc12272a12f2c6261677ffb56bec2bef8721d15f2a242cb6a04e198271e1582eac92de17ad8c6d53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha39d628498bb32806126495b30fe19b7e3b7ce5cad9fdcb291178dc1034582f24fd6de56568b47729d0fa61a1e7f94e5ce20bc87c960fff25da0549637485a184294b40c23802458a4f19b7d62e358cb252d032d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88a72d9bc341ac4a5f90cf1d8d08e3293b208d71ed57fa9690157820530ec2f12525ed11d1d35c82cb682a521864f9c955d5b198c34e5b20ede82bcbf789ae50f2cd3abee65505c9de4308b1bfdae99f6dcda226b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48bef9689a92d3b17cc616ff96dd4ed2c3be261cdfc6ee2c9a1d785368f0fa2e04def6614d73ad0aa309af808b79b2666aeb0d5f60b05dda71273f3ce735788cd8084718d64e1bbd594f20562e764b2d789501b88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3a15f64b25a41b8d4dbe66803f1e4a61e3583895c832e1cef172d8cc39549ffb8a6f98b98b48d14e71a50538ac8bb46e5f9334279402bf229085d82d2540b1b2a0d65f8590ab695351fde86f66c08f1d9d1ae79c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2511c6bbb72193ea8e4879d59b03e2b39384982eddf0553cfd9620333e3e22e39963870131ddbaf627e3c1d21f2a14b32bfb8a8fdddf12fea4511de16dd18741f01633df769ec8d2df19adfdb71991f1cbac00b96;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7af94e63058da6032d62d6d605d1dff3c431f752bee9c1f013344049592170e26b7be7117ff14e7b50b0e70acbb7d91bda2217ace7a73663a4423b1a342d11417fb0933b1263b62c7d81ed25c4fbc65bb5f8f84ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h584a7a1b9cb68744673426d3253ac83e8da3ceec19c6be8fe908704438e93e27e8131ae858b5b0645c6e9aa9544e640a4fb3b0582c3e67c2544d2ced27221b0ede9b2e7517b05a88805e95a7b225236506d448619;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54f34807f25b32d2a6c5dff571390cb473f225bba2345895bfba0476559cd6aaa10339c8b195b8921b481e84e2b4b7d37383dc3368721f8f9a11963d30e2b555f23d397a587b1bf2ef4de7f4d8a828a4f9b7950e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c0b70fd4d4bca394ca335571d267afa27edc6cbc5b99c15da99b2e76b97367fd0e571a90b160eba7b63c9bad6863942874cd1937daef670da7d50c626b3f70981eb6e8766f2a0d15d1ee4ed60b9139475138d1ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdae50212fbb4e5b3b9069c6addcda09b765b8f7099f64a0eeb7d7108331d5a9683bad23e559741c9be4c99a5d5b868d8086b86bb3a4ef07926ac517a96adc6c5c6d9ee44947749693dbd5476e3d5346d6e77ca836;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70234c745955ef20402c8d926e6e7752d2e1cade6968b97fac382244fd36855313e566c923364a9c889f62e6887ed62ae39cb878a8c57d993dc1808a55c443d556c17195ca1cb8312222a42395bc0ce36de1fd898;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h187cebe009faa98b309757b2e89dba9aff6ce5173fdaa2d2cf505f1b9c7ff6ca310bf893c4685396c5a2e0f2ec3bdfdaf3d78b80d5ac3cd993a28c32c850968c8a6d693efa31da880738a805212904636074ade7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb13e8c245262501ead13d3309bdfbb01dcfeeb5c3d0dc8a27a21ea61967c137b34f19f2a3ca9ed91176dc30b2e929132e1bb168087acc58af2f49358436cd91ab983b8c279dcf45a90cc65aa4df7a09d27c631736;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e466aeccdec8cbf25a1afa2d8067c8a6edec8fb0a23aa333c0d0b643e63e3bcbcea616d130bddcd13a7fa7a93cc6ddff1c74bfd754631e7ff6622011bd57a962acc51ffbb1eb43e41051dbcc7b76995cf6f8b666;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd021369fbde624dbf5d00a3d5302f06b75ffdd09704e38e9ac1b09d705d83862818c565a761c06b92e2d79acc93b2d4474310ade2a2924407c606d4f48ceab28e13527a921f3c372ccb2bbcdcf69fba57792c6f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1996278bbf387beca6316fc695d3547d365fb2703c6c2dce912897d6dd4c4c0844d638c426b7698aeeee288cb9d5f5f8adf03288bc225897d492239acebf7e60b55396e0cd85e78087bffa2035324600c5180ab5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7e56f8b9aed1c023e1cb87d4d0425e571e720756e0b0f7e2f7d3c3518ff510d7dab2cb2e9e40df3d7ee925a73165a8b2389200ef0391598908492dd2137815c4de8c36dd73180a20ac896fc8a7aa18c63fd025c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c0a23d747010394c6625b4713cd3a59ff2ad504d561f68f8a5f6bae05064aa164e3dff728dce2485bb9d48b1069d50271254134e3464c42a33f7554ca0cfb2acd75dc441577760e6f5ce979dfc1e3b11ac1d225a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7d2159b5655c589da1f851546572ee479af8fdec74000ffe66e179fa91c019c7271a88479907b4befd92b82cc63efad99649b95ea05d9190754e5a0e1dd458a04cd310aec2997fbe2c0f03a903c2edded3153658;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d886c64ddeeabc2f6872c3cc7dcb11822a9405d91541296ce5c4f6321bbe1ab9ddfb3e133f933ad9786ef2333937f023d88328fb4743a4ecfc1cb91101e37fc416ae70243682c2f98cb4209851d8a050b913a2cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cc9dda67567d8be826b52af5b6805aa71521dcb5223bcf4d9a7f9ddbb02f43825898d0e9751451f0d0829993bf9072e7286e0360dc1a25bdc841c7b1b2aa5f674ac92d5e5ce1d217508257bcc288d1532732204;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d914a670cf9baa843c471fe25de428ade70e6f608fb9be8c2507ece3aa7c6f4e9646beeecadafc613aa4f6d966322d4297068d9c9cd7e9245f5fe3289e83cc71db30770a55ef126229fee3a63da04445c43683f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34dcbff66bb8471e698e4e4c72b5e6bda287737a8005e871e7841a5aebe89f46503a1233c4441736f70fd513d47915d55e72ac970c43f24857a928912737b5e025a776ee8496fc637e1d545b6704ae27cfb82fce1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd406c6df8f33cdc3ce4570646c6261ce2895cb77537e7a13f54df856122725b4f0c3e340e481edad739d989d7b5f2ae350422403caa3be6f312b7b46daebf6014164d02aa603e74ffc220bb91d595b516651a8c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h600d270e0c0c4ac97da9c395e28399be2e67207b7d9be4024b9770faed7a02b71568a08b46264f9c6f94ce5e07f24cf04e1351eac084d4fdc4c96a2a6f0bc8eb9524769d6bbd569cdaa7e2387a78e78b70825629b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17bf39fc304525b417ab8a05d7b9fc59cc23c7732c43b2c020b35d9c4fe908c85663686e55d5257aa08249b9b27ec081228e8bde74edf7663f546c5bce1f7ba36db283ba32bb68d56f1a3dc317a80b9bcc56abba9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h154e3df743db5df1c540e4fc9fdd21a6b44b26438a38b22916e511f17e9c2199c31aaca88fe8fe03df57c882824e48fcc4ab88e4f21565049d822d5f56e64108b303e654fbef1f9b97d7d8221e1a632148ffb72f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28c2fdba660a4d315ec5cc30816570be64cc1f314dbe2f3103aa8c93130ae7a8c64a2f6db993807adb4a8a783c18a256bb19cefe0d2d61402153c43cbb2ba6fffabb3bc70b77df5b3efb6a5a335a3b13c2d537f71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfd5371f55ba378306af895fef0cdaf950a62ca6e56ec361bd9081b754fcb9114fbded42f850352f8cd9283749019d3a3ae3ffdabee267e5513b327cbf430750412735662cd9aa2b0f7f22512675142d3e13e0d8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdfbb58990e0a5b9000a61377097d0d16107811ff596dc5086371cbde5a8c7e075a190336b9e2377de76d47db4d4109ae182d4d63fc385a208dc77b5d46f4c11239f520222d6b7ba7c2c43c4a37d5471c10d72ddf3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha07572278c25f4e29f5503825201c0721c240d89920f871b15c32f5d70fc637372bea99f20ab4f3cd842adb861338423e2742597c290862a8495a3a795bafa1d99e1d8c6d099c00886da52075e96cee07c5c6faa1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h218c4d5abe43b08e0a54c2f0725ef6d8f9a44f495613460ab97bed866e0288f4956084114537a7c5f5026563f816808e80b3a2306c82661c8773d73827a229c5fbb8725a7a0c84249f37b70ee8738c8159729e67f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca49b51d9509a06b7186c111809af3f6c522f1e40f7dc4f68f5b5758ee2691d49fadc5957a0e74ff0b4b394d1716ab3993a7b843d1aa0446a6af1722c0800dcf03e9d8cd349b39acd747d1d54cf380356a3b48ea7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h300dfa43f641c790af1bb43a7c18db6867b0eeeb821453ede8e9b5616b487fc353871cf4a349eae9d75c94ddea6183d8d4a592b2a2a9011a9fd96811d4b77c2ee182cb44c0066ba0e639fbc0d3a81351102d10624;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha83cd8b215c32c2e1bede11f23dda189f3bda986887c52144f869911b30b4ec59ecdbf805f0f620a03a731679fe874fc9f1632ee3b24bd86463c0f3243807e6732d438b0f8805228011fa588d7861989613e4b0ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ca34b0215014946458c0ffdd381dfe4736e05d2a6a1018c5597bb0166af749c78b77709cc25af0df6b7f78bf5af46610452886309d9711a0ac07f5c795664b88f89dcccca7a59098d46a80f794ec91ed76006407;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d7abc35a15794198baad163c77f1791458e07816d28ed498c78614f418383496106e59701409a696fe4d64fa3ab571f9fbe3d3b1d69bef01db61c2f1c9497ba8902127e6a547872a2e4db05358a16b38d899bb36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf89955543f260522f906720fb6bf5ded24ad6e2a590de38a807ea98574bb5ce5e26d6859e70e46a113f3b8e472bf3032a4ea1f746625e0f069807aa9091af64cc96b8fe48c6df6a1cd7d44b8c702f1cfddc2a3b3e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21823bf5f9013c9dbc0af8c272c0a561fbbde4c2abfa63bb1f0de09b3689e899e8f62f6943762fc7750f2d7b330cb60ed75caa0afd00589df05791c9dab3c5a9e1ad30f370d12e9081c289698e75033ecdc419d08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbec5f1e218aea8fabe35a26c783a360044184df91517b7627d752ffede5ba837b0c703f1e3378d1e26b24e63f40681fe9e49bc594d4b3552b220c3f679f0ec74440381e6cb2e39abe2f37ed2f4da172f4b74c26ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4127554a0872143e6f491ad46f5ec7443e451730802531fc1a5e9d8d35937c729e75260ffc5025501cd306870569d25e48f4d5d8543018711d64436660050e673cafe5612ff4a708b836f02a61a7def4f9debabed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h755d8dc7ab0066bf39c65b1e74d6d3828a073a000ebac7d243fc7fa3f63861c47f0a85a75bfe10cdab6806723147eaeac14281a316ce590a2eefc0274ea316bbd949479cf4273b2bd915d97df43743146a74cd7a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb61463aca75284be306eb439206f5acafdaaed2edc21b61c5e9f5544c349a07d1327318909d2ffdc72e628c8729ffde1e6972efceb5a38dc6e31c8c0250573ec0de2e6a51356f84d836025f8fedfae8999a3cef95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde3924cdd2dec72140442be59364665c635f62341db12bc7eee3991235d465d04aa1a7bf74d6ba4208012bd213505607e19a1864310399cfaea00b635b1bb5605491348cd6553ded5eaa771fcbe5a62cd60270165;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0427f13eccacbf7b6014822c507ca3caf75880f0eb8001edfce5d46cfa718442210ce459a38195cc077c59451e85253e2a98de2053e5551fe1f8ed465f4f701f0061802b93a07529767a7329dc54315129d523fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb690b3c7e1875a24181cca6210557a800082d82958dbfd63e0becdf1bdcdbbec3630f5f5d32b44ea1a7a5715a573f8e0c5847588bf7a808f478d31377bc3976069e1561ee2c07cc23b6d6b3598f2e4d0290911355;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf2896597a25c3216d337b55a565bdc446e7a7180015e4ded2b9e56bbbac1e7047abd37bc7978d86d289fd4ff8ec1d800b8658a47759d47aedb08ffd79cb5f0b58d25a58a259a8439005bf553b27e0513a64911ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab66fc4730bba7f305e1130ec81d42168b3b776787a981d82563403886ce1acd19f2438447dbb1e693d7e64e1e24efaa05345fc007cbe5e82a899c446ecc2743b0abdbcbfb151a91ce6c3154283daa0190c960304;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h396eb3f0a07c68f45ccda4e04548036acc5bc9f7877c6bee6e74cc33aeefbffd6889877b6c6ccb7895cf1bba7362b837701a6383dc9e335323edc6201b18d8bff575d9fa4919b244b15e0d5a9510e05362817933f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25ff2c436f760f6a754282d9a7d10bdf6db5aae5385152e43050969b99604326790271b51f4c0208f5839ae5b8f2a2bd0d5a93258b276a6fba756d6bd54453e94b74ce4d0dff46300b10991ad275093227a3f2c34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h615c1b2cbe1495330cccfd591a110308366caa1d996dd0c15c5f776a2f4cb1ccb12d2ebc41d95227cb848ddcc822a5888d542d192119541aed8891e861a3b8fa08f2e2867f566d1697a1516b74ab5fbd6576ffb5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc00feb63bb8f583f8d9386b4e767fae5f124189698a3aa2fa853ff194d8433480167154f985e556a74c82103a0dac0416a7dd517441153424b9b53c79a6f234ba6b8a711ba52982739e56b2667a82d84b722d61e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d321af460b4183565e162707b18ff8aeb6b4c5d6a53860418a21b328d23a5a2f6b9eb46ba927cc12bf0c1d6d2a1f55a60b7b429d44286bd5a29af055ca3f75ea71cedfcb8d05502330435f900bed45a878a8d385;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3b5eee023ffecb542d755ef43cfa18afa41895c894d7b9c19c00ed6ad104b44347c0df2ada5dec93428b05e34427566229ddfe4f7b8d86855df24a3ac681324ccd5ef87c68016b2c5211a3ee08bf725ee680e305;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe8b4bd94c24a95a106ad0125e5cb5bcbdd0d344ca6ceb975738299cfc2df69e87cad7d5f58be1a4c98be2c4cf36372c0fd17bab96278de78fcde879f93a69f01db9305de914e32f07e790bd894eeac968b7295bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haab223321599b2c8f862265734ce6e41928f02913ca20859036588b695ab6aec2106229e411bb8f168deca0fbcf11b95ae3fb4a535ba1001957fba1024f917ccde8c6143b31702bc48b639177dc7c4726139c3ceb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66fb671b3ad44e2da8d2c9d7ba930085feb63ee38a7e2a44aa72cf5ef3fabbb48dc93292548a91e873b640e08966bbd67f99b740b75c4db9fcba208a193ae5e59d8b6104aa84e921b272626797bce9fcde18c7f6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h507f4dd6c96c81b21248d9cfe5d42d97d02de034dd915d09bb6e6ddb201515cd8d2406df956840d2b923b66cdf295002d04acd1d55364aaea5d4d118e743457e2c1a0e754e62f4fb9ff2e17cf72f32935aedbdbcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc77c473cf80dbf6aab2ba1c488ae06e92caaac6044c40125b8c70709861a05b6012dd04ff438e17ab364f3d86849c37c62093c17bf8dae167b1450122a3b247463dcd3fc6ce9b3c0b7579c4e05505db023a13060d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18115656ea745256df9929f565a3527b52e8b2b26b6bf73397e81c96578ea7d44b985bd2d6544f0eccb017921dd30dcb6e224fab25eb3b612ea80eeb3d433e2de91f2acce485a15c9ee7eb59be1ab78261e99cafa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb79e156918f6fc4b69f67d49014dc91df16be5bc496130d1fb8534387c19c3447ba8763ef977aab1b04fcdc67277ff161225d39e942ecac1edf430f0546a726b9c0127f4e55a23cccd9366bcd575a3c6fe6384e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84935455939d190cccc4f6ec5b31487a42f5ca3883ebca0ff2e3511bd7c2b909e962253bf5886d94f78d93d23d289d9c4313d80f817c4a0b8b6a7c88aab14bb3ad3e3f3fb10cc6c78d8c1c2e27cc17d09134e36fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5420da578aa9a5961324d8eb06bd04bd3dcc04996478fda8ec32c82fdd09b18483af66dfe8bf79315c02ccb812746c776f95e020212ec29b2882241c25441e72ec1182540838db8bab9e3e7b5b0cf06035105f3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a733eb8404fcae78b770101ef5e90c914e2381eac7001cc76170efc530e0b3b81ce6a601fbd89ca77d93bf65a9c6520644007387c3b37aaf23eba76d2c170a4a810f4a810a6cb171e2345d143634e22312419828;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc541874857ab2800c73c2620e828508e46cffb544b6fe498cdfe420fbda24ce1effd6b7fdc8349992f9c4dd74c2daa9858b405adf602810dfa247a8bb682b72eeeb9a3a945a1fc3fe01bbb8c895ae40a4623884e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3b616f35641c01d6b75e8df95952888eac72d4ff23f3ff5d434fe77acd465ef68bb8d03d8802a9db82f9899e4dc13d4ca4d6c56f2d01764f2a1c8e7b26b5ab5456857fe503ff2cd22a87abd2539f9a25569470f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd70b76686e7fec97618e5c28fa074790d9a100557de7507b6cca4db8dbe3c94fe1ea2559bbeb518c10a8e18ead931e953a0d2523e3386e78d6cfc2233f98e8914c69327ed0525e1f715a2df62d0bccfa04d78856;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14e9cea39765948480e094ca8e7712081833660073fa6db8e08ad8eee0a071ba09b81b33def7f6a1ec81eecae27c5416f86ffb6c430a510bb3a2d0dea64c85d0572e8163efe9c13adebc94c450efe2d25e44a60b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75c8746dd37c70975701a3b9919ec3f4d935c7178ab205c5eff7dabcff4eb3cde0a522bf0d9e7fa0954826864170750f4988e6b43768fd9367ba3710e3350655d702d7f79aff309d860e961eaa720b51d87a3805b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h565e61129d9a17a0cd4e6f217e71fb1273c16c1f6f00db5065afdfc880074639f3f7772f07f246208b07b77ff7860fa3575a587f7ecce96291ce21acc5ee5caf99de17a18b6a6653bbf2c583ab6dcc61cda3d5e3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b7431df4d5ff0cbb6ca6b69fc42fe33ce1b12b1f7f16b50e31d7626dbe2ca95394d4e64c4dc61e00179c7a74daa1221001df64e6c8f097e64c2e1281422db5965119ff5c5dd8abb45d0680e21f5699f2c7288d8e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6f6507814cecf56be7cb84dcd74ad12f1095444daa3ec508c010e58f644ea73156139e3cbad50c112aadc5209f7677e82b6e432f1796fd6e7b6fa7fe8af6e6268bfb49cd069cadbf1874272932190cd5f2ac0ed2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecff6f2b590349ab25203823f340aa2291ac898e585eba5369714aa3b46ce435f352ac53550f8ca1f431d89f94300a9d8c5b0479b094b5a36cad35d746462ec0e21d2ae26ab41fe118ab0d83caf5887031e4c5b26;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6933689841f6ba5844c91e65bb3039f7b4531cc16ec8596b07941ac98a7c7513f4d68afa83772fdcc06950ec106e775bead71e73a081dd440896c59207461fbc2f9c04401b2b9e5a25ca7b23980585a4335e2529c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfd99002cf5e9ee576a60833c85de1d8eba57050ab85fc92ad9a1313a6d01e05edf40977c9fb5409b2e28f35816991b6a18158bbf6aba63fec8fbee6482936cd3775cb78063add23ef1876b25a2181ed3545ed676;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fff027b096d65020289b40ebbb9d4f34f615bb78cfd1e24d8d2a7a9264f371ce743ea1a739d93958f2c8b95d6469824ec50dc5f405309864603f9ab04a083727df3db868ba2782050bf9cdeb4646cbe11d8bb782;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h330fc6e4d70cb47c1bb35bc25adfa9c50fa069737193d0f6c4195694082fdce4b25a1c27ed087ce9b6c468e5512e1cb502f221e54b85ca75696e83626cfd53e5488ca850bef498bada2827e601b90fb9a5ae9fb46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9aa328f2f17c5a49aa9ce06fec793feda771a2737572e00f1a479ba451515b821280a75f8f00c80f9e02a5148011b7301bcd0aa58fa5b4b66c58b0c48a5b9a6d2177dbfb625c8346f1416de5de3594d31ea2b086;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb1e1e6adb0d023de0b5010ffd857f7ea6682ab1f4c4d22a5437315091d8fe3d0275f343f916242d2e8c533b1cab2e76c0fce233373e42a25d20fe2833eaa996130614e2e294f545a65741d28bc41c123759e6313;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48a8f014d74051ee841752d796af3036a70d3f649e24250dfd3b9c450b67fe2de4b63e2b1744df17e48a18fb0e8edb2c3562bfbe2bd0c0ff40bc0ca359bcaf09d8de1528d778c6453ebba7929325e4cda31050e3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd70d432ad2bdda38f3393fdfaf1cff56f36d31d25f60772f67390a2e16b5bff004d9e8add7ebd1416d3d0b1e53b844395bd0122c47e71a0ad5c993c6b98895478fd9f0eefc9205ffec2e77be7524413d783088c23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c70fd3390ccd2a13e05d288acd37ad494a02edbc70dce644e56dd55d3b94d44e8411af35773ebfaa72f5cb96dbc87d8a860ab916c6e9e600d82562e4c91921ae077fb1c5808769db254ba0447ee52e4c7cb96dbf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e41a7f90011120507580d45b37e2aa380a49a447e80a7983b4c03d81bc774c114d1ee70bde0411f3386eebba7a3f19eb1d865ac82dbeef704cf1f4a9a183764b78f95bdfe754359f4410826e851fd67dd634fbe8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbd84fc771158f9154376812606cec020e6b33833ccc5cb4fec370e5f098e636ed85e49a208f52c713a3a71c0cb3ee8736d158f6a6db4060cab0561ab77b84f1cfb714e9a17a7a53c7d11d5ac5529bf0ebd0c1427;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87077b9448ee7c9477ee9dc2a488af6c2ef11c7799901c0900c283614939d2bb1a51ddc6d8543e22cdc121e17e2be0eb6bd4762daaa1c362654fec57380ea4f114895b09f9b7a74b6c667a9d3dc2582a2e4903116;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h915c4b80914eb2b30d7279731800eaee97736cb7aa0c2da079d8997f987fe9e8635fdb8c878e6fb8058d00b4dc310ed122bf8d09bdacd19e9764b2f960e7b59c600c44e6e49749591f93e61ee097c3943e76cc2e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44ff4a410e4a8ce4d89b16e32a2a7b76b48b7e7333f563d1c7ebd75f4b2a682e9d19fbc74d631303407d16d6da2117b30176bcf0cbf3e44aee0365b7398f52e410f1abb58d8299522938a78e312aa7b5f80d42883;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c8fae5e701640e61faed0e69083e29936460f2f4d9d3c3357962fcc878bdee7a315bf6044b8da33ad09cada59ec6b12cd9946119ec386f500833f597a316d05391188db04ee9f3bc8a76bea5fcc6100286564538;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60ffe56bddeb40262c0d83f1c5e06ae2b36b163d799ebefb405c14d30d8e6aa6ee0300e5df6a522a2f0336f690034b62e229b0f008140869ff41bf4f96b6f2d2143552a67fefe786c5cc749743bcc9c87ec065823;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85486299cf9d3379595c70c631480b4100625439f46c67205b191e0d889d7a580ae9522c5da331d90532f4358675d84bc3cb4d4519fce29ae11b89e9ccda95aa3fdd8dc7424b6237c533b1469fa7351f3eb1c1341;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eb4918537d8a6c53069c34cf1067250bd7a8d277e1b6ce2968a0911890f00a130ca8878ed5dae86c14bc6bdceb4316968ef91e0dda3a120df56adc36d87ff82fd91161c4a717d951fe741a2745b4cecca2aea100;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11762c78bb08b6a7e8d3fdeb10139a9f77fac19a66c85111cbf742cf638430a988751d6881729fcdeb7b44050840d070a1a8463403ac59ef8d18f4099b67d0bdfe2312c43e5856d0346e5a6099c66d146c14c18cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd86e560593b7788d769bfec13f2171075b25e3ee86bafe0ee670a18f68efcfabbcce632c4263e3e02e2c6e5709299447d20ad3da7f3a330a7ad6054f53f03d3c206ae1dbae9f97a5989c6e2d9abcb131ae2572075;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc39720cc3946b2ab8631888696c18b26ae73c054f2b672cf2cbc6d2ee8f5cff66982a039c85fd7b68e4411791fe032af814bf41f55fa81e14e6e68657d22b79d85c66932f47df92da6a6ffc07dfb2b5c46b991d8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff51b19b392b3ac46690f3547978b493dc1c2703d8d8436e52a09731f16bd221634317dc1f9ea68891265087794b1cba0f4a14f662e26e17b682ab6ce1c177c7709772756d72043b64760c7fb84a4d5f18ad80303;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92cdb3444fd8df79856a0b59cac4dd96f32d28abb60ac7d636ad3d0d1c5d779431a76cdc68022f488fc69b6c9cf5712ba8abfc2cadd4c421c1b80fa255aa7510cab5a5b59982a7d74df593b675e5d2abd734fb089;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h473415af1e3400ff8d2bbd78567fade8f45f21a405bbc4973bf26a21b89742385b07158aba8630e24326d0821ddc1f0e34bc0f5c99182914226d905418b12a54f6750ae983dbf6d613b5466622eceb42e7ede03c0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33f177a24d0f78282f46fcec43757a2e5f6048a2324e9c23326dd99b76bb04d927c38bcc86269d35e07cf08ef0d0d49ffd7f5a3aa658530c06c22ad652b235fc7fc6f6956839a1f45c14793419c44f1a78a6e064d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7073a08f93fe88647c23b511c1178cff4aac8100ecbf83bff8bc98b549a4cfa74511c18a9a52891318490977e8e12ca3945c2b7997d6a9e46b26e618f3349c86cbd1cb2418a769ee869f90a612bccd258dd12ca53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7707ca3282e3d56f39dd61a87be70f33b18bf58338e1a91dac17f6e99ca8105dcf48cd0ec6648b061533ced9a5cc4bd0c9b378c38034a34c7485e0758e92b1c6b1f23f7c2719f7e7097e0d4fc9e03364bd1ab4c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e7a8b3e7f91b4363733117f53772d16fd9c72a6fead1970cd895e8dd7b1f86f7e7161f77bb7638cab6589aca630367f9ba398a8a249c4f829a99adf68967b6d80fcb2a0feafef7ae5409d1bdeac63f28d7fde0f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4279d8bc3cffa0db09c53fcee844ceeb5e9521d9b8ae05f9a1ab67a6856d31721ccbf7a0240e30e16d91aadda8c0c94ee7db2834205ff487770e28b6947ab3b7ba80c6b336bbb80bdcad97ef7ece296931d8a9c46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd344d08840246c35c21361ae2c409f7b78cf8af6b79d0828e4717deee60f7a50556af8ba9943026efea772fea511ff535bb16c21c46e9545cec9541c97f539453b7164805d163f46b507d124b1aefb8105b78ac06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b5a2af75e6b280990a5d5ba1f5dfc84d871839ed952ddc9829b6bb80227ffaf48aceee9e0ab423446ecea595e11bf1f959c7449efae9710e07a922816ff632aa53eb5165f465e1e96d27fc55efec1a574bbe61f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he676eb810b51cccd3981906172f2ea562c5c260a773bd0b833da5e5e53511f6626280f4834dd5829e8b392f8b61f509b427fd87c7d0ef20732ff1ceb629000a35b112af6b500e4aa1afdcea8b2c057f59ed10654c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f92a70c4b925c26e0593828add46330743a0e8c66d2fb800567fd973f2a01d83a234750d604efcda8b4a0733b1be3230fdb95036e39039613ebade6cc2db47ebc048112835f7c6972e8adb67ca4ae3ab7e6d8049;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5e7613d0e0538a6aafbf94ab9b0d5c0037df472d8767d9923a2777b42d98dd45c1b33a2d5cba035b420ebc36d27f4a1d5144bf5d34ff4b5eeccb50033a5ed05fc14a6ed562231ffcbef15b77366e88282c64de75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d2b3ad79c5d33589de646243ef3cf5e1d231f0b7529861137f4a0b7ddec8a6901bd173ebe0b14fbc5b0d4a82570151fb77b49d8230c9eea6a264d758a3bf3ec1eb6c5b1cf27aa843005e42c1b8ab4dfcbb0a2273;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb5f301838ad362f8992fd1230d99f6e0a6c9401615dfa7b8deacfad42649f7e370a1b88a531f36ad38ed1de53f459dffc38e78dbf72b5a6854781bfd75184d3883965506c66ea04b00048b6187a84a90ca850605;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14f75c4c9213282da28377680ac543ff42e1f41e8c7c85197b70a3042cc449a7cfe3efcfa7db44b5fd613554c04b4a9d361a4dfc6290c75d39443d0264f45032b6bc6184ea50a678814bf6c0dddd849b423852bb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h450a7499d3528b2766e4cafa361b3c4333e30cc409cfdc8a7d6988ce00e0393ae92cfe1db893a437ef91b178fccf9c44317730e13b4addc99b0757818f15d8ab17cc9c8d74426e9ccf14dfe4fb86438d1c2b775d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25b6226c1ba07bd569f52f1528344210c861ec8d98811e1803b5ffa207eaf2bef250d0a8227d4cbe275b555c226dc84dae4148342482b4f276776267446ce859ffc9a5c1eb4260e357b54ba8d31e8c39b1b9dca40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9421b8148e7b3f6f6ab7cc9b831381ab1b631c7df7e8efe50711dbd8a34167a57949d0dadd23e5f1e34dd1c48b2aa6bf32d52febb0b5010310468777e656a215b39d34b0d9b58fca17e20e4288974724db3107b1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf367ded667dade2f2e84869ab46fd5338198b25e2c3d2b8072adddfa6358a21da145a850c93f2dce0c1816fed8af051d015455fe925c42435171abfc7147e85b27708c3c37f9569a634b525628fba32427d49fdb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h830bc06857c7797dc796b55d56d406997dacf350dce7b00f2871cdf1213dc1b60e0f9aad292e44b1816a29f609135dfe679ec1cb3ccc1442b92fa8e74b95da8fbf1ceeeed7457cc41eb29d72f3e850ab2b29f727e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cf9e1a4f89c37459a8a592adb363f1b725fb52ccd68c139c7bfb921daf1e642b5cb204ec6d3db858f38bf96e289109379983bc6611d9d2a032dcdac6a00e8d431b6bde32c4be2f379c82bc9a6f5f08f258038c7a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c1210c01bc549dd440b6406143c1887c29946ac7e57d8485003e82004da03651786e5630d7879af6a19af3fd0708519c385408ec893ffcb30afe97f78e4cd2b2ec7b5220e0d703bf44ced9ac169d826ee16defb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96335d564537a86d29ff906c1aed4212aa865e474b3ec965fe1684032f74aeeb0a89158649fb625ebf5dbc20843a474be787ed971f0fc09cdc96f1011c45b3f717f7fea2a0207705291f5453f42b0789f78b317d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfea32598e1e6f44c5f834e52007ed86c6297750932ac7be4c8a4c879d730810d07ec5e483dfe750e47c99feae456a41b66511d36c56c817b83f3b401b220c1c3057544120ae41c569f63f243f306184fc509ce21b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h998c40dec92b49f5e7638391121eda22894a128806af5f7c44e547dafd32474d12d8db1f930ee20181a6061aeddef7f6107a9b371f4bb05f3dd4ecb1653936b6bb746138bd0860464121571296f62f4dc9aa90495;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb6aed33535646b3739893f824d999bb1a2a91d421a19fa1b295b5e1f36c9d7b581004a5fab1fc1e6238e974c9766658459eaf24179187505920509475b2da0a1143cf7c8fece74c3cf41fe3626a15b32d40186d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h897771aeea2848dce18cda46e162913978d2d934766bfcb40bd992b83c31f18d23ed5c1fe5de94995a47694d5714948209e84f0994df361bec1a26fc998a9ef822e789c9b74bae2647f80c706d6b46726882e8f64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0dd40ee325c534e72a9bab2c7010c1ebb35aa3efdc39db039f44af7c05df87885b05fbdd5e473fc04173e8b2d5c010ad551bfde8d04e463d7bab65ed509a1a2ab1245e22d8c995af2e0d9de9b708ee5207c7c3a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a398b09565e629db00e683db8984080f2dc746088c44e897f9e4184559f8f036fcc49e48062df0b40f4952b2b602cf69b3f457c4bb9f641a0c9a48aeb76489d7d1fdff183db81fa7250e49a87ea4de3a4c65b35f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8eabfcefef1978389243e8ff6311243620d4b224bf69562e89f5e46ec2c0fc8885800548387db0de9ef6fa098a5d68f67a16c73e8166496c98cf7f52e402591ac19427ae40913b5dcaa815f57f287aa7869c772e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50d3ab86753333aba08fed3e0f82114cf9372f5d2b84afdc67c66ec4a4e34875131e15a063da42fe9348fe9fab542d4100298a7d70b6b6f384f62a6848d9601ac47d6b55f10bca26f256bf5a682ad12350bc7f05e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h773e70beb0fc2598d817724248ac73fe4f533e3d8ee77f8e08eb9065a26bdb329ce25382bc1ecce846c3004dd6328eee0c0d7bd9bb21955310980e56a11c7720587ecfdd19b1248c1e8b090498bafbe13aa4b0c0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb52e8ea00146c9afe154a572ba844720a909377aebfda527f74b7eccf2be79ddefb558de44cd72f8abdffc72934e96a9943eb55bd4c7c1e45c6368ba678af49d17b612acdd50da4288e93951793c93c4fa0f71ab1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53bfbd6f7317b4deb3b3b479de1a8960b5d4b028fe4aec84fc6ef9d7e6be93685273d05635c84647747876c39d69a829137362e8f1fbfc148c14e322e37abc8fe1a6b7860febea2af4c5f0c70be4e3526ada5b61e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86ca356f5bfae570e471152b043c5bdd5eadbe5f0d9658715368f95200fd287911b62b206891f103f18be3eea16be24cb4be240cfbc15e83d8af591241b229dfd9bf372ef2c4d90b7940c4e7c4e60a5348a8458c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbbb30b249193975ad768cd05bc4b59451a990866bb9e18a9daef8cdb8c488edb893d8afeb460ad52e2d4687a7a17177fcab320f7647d6d6ec13a5419ced15325c705e4a42ceb50a3186aca08f3414b81df26b44;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42418952d32d2f67c49054625b1d37f4770244977271952af48d68dad2761749612b46e30b261c1bb677c608120a6f3e15b65a425d9691400dbe2a1340579566cc87bcc5cd178fad4d5cf3724ff5457a104cfc7c9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he919592c7b8a9accc6e3dd067c9a93d1776626a74465d81ecbe55d1efe19af2c64562acb5829a5700fd59726892e1693a48397bb54d6bca2bfb98c117f0f5ede619e900b3ac931a9f0035d81c048d86e23e4892cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8141f937cb09d95720d5cc59701e253157041d5cdc69636877b4c3edd654c612912c9d76c83f38534b2a43d2b105f2c27cef258c2469183d54dc12e4ef118f604c54306a382e74f542bffcdc2f3b3f853dc443636;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e959e19635b7d50fb8e871698a454b8f6ff09cf26601e516e175f8034fd935303679e7c235a3abdbb3f379829f950082426b5fddb71371d0d33ad1a350e8605492a9f2ef251a07d9542c4fb6e7cb26ba1e5e26c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac5ece7c316180a8d1562ed222624986b6a8e7b1d6fd3eb070e1d847385db6c5a46e5d0ac06afc0849460d514ba527ff97bcd7aaa354ada80fdce6cf98df98efd75f9396e62a68c7ddc6c833c8d53a074c21c7e1a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e499f2bc7a10f67f252fbe3c705aea23eb35409b3d53d95c87d843cb4712327c4f9880f85cf7015d6e54c169c948c6a6ffa2d3d3e1b4d6778b480ced87310d0c548724f1b31bbebfeb3c10fb0527f5e16b7c5ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf8b36ab7951771a115541f0dc7d3360788daa236a6edf0d646346ba60d0eb6514b912319603a8f792890d94b979b388a60e4c1ca8ce6831fd243786022bf8494c76c4db951736ce082815d6ecf5730425d088c9e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ffcfbf7ba2c8cbb318c7e53a0dab1ed53c668a46466617c97680322c249ddb12104dff5ee6838626d6ac6323aa1b4bf787a2dcc656c5cb427a0b6bd28b23dd156334ee44233cc3ace34e89c88a8f4493ace2a661;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c99ad22ccf505094a6707e96e3d449dab644ee6bba4c537377d16af31cfdcb127c169348ec168719b50d65fa72af9111a122209f63bd0032e69a2b67ed9aaa25a6409938e1203a13162c00f03f12854fb9dd413;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba0b7ac97c5306a6a91557faed88126bebe51ef77e2629d894a0b9a8ab1ac576b0725052797d7c7e48fb61003fe55ab03dfa5a369a5385bfa5b02443e07d1d11a39d6dab00e8576ed6649f4ceaf1ba3eeb677be08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8605d66de86829ced655e300517ddb210dd65eaea40e56ca2ff8c7883d26a7dc7ed3f9a837d6c5af4213ed7442db8d9da07303cedae5044b0180486834da7d552aeb65da0a788c4407f17cf0d9e7148ccae3e334c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ae0643d49368666ed572a871cc77787d31a4dbe0b43cf41e5744161ac50e51c2ce1dac0f0027323f6e456d6377f8a37dee42db6914d0ff6f586fad3390427806f5790db0558af6fd82205632c59fe8f53b092a03;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaaed6a348494dbbccb022aa86124e1c0fa5f9c47926a70f230d654ae3879928c00a949d5bd4adaeaada34eb2357dc2674e484895ef228512b9cf186474fb368d61debcf387da8878a7e7634767007dc258e99266;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca59240849b161b66d905d10a71837e63fb19746a8496743bf9b3717900ab53b7d0ce52e0546c7166914027444c4d4d05e675b95273456d4133aed0de360e11fcca0c2b5b3f4cdb81670b7bf15ca39400816db715;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82651c9967b3ea064686f9e5847a008a57f0e10b35545ae1b5e24657a8a359a70e40a2dfbf52a95976429cf8e83a8ed4b43b509195cc9925afb09382fd6377084fc84832ba5293efea0f739eecec5af24cdcb21e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2be2f9c606f2864c17ee43ff0b7d81eae521390a4f5441f2026519745bbf5c4faba0f5d070fde07823cebc024a8d3436c6f1c55a523fbfcc25e58918b358da9612119f168445f7eef5e6e109d3631a6d200605e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4221900d58f914f18be95c3b652fa277887f999e99ec0765efbbf2338b512397f72a83f6b69c3f46d3f7836ec7c102d72bf25606b3a8f8d7a0144aeffec67f61e80a40e108ff2820eeb361affa6a699cc8cb04d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd32608864d98092f039c495023272ba113cc9fdb0e83dbbbbccf8897d4a6c7f9fa33c52c6c5c392a94fed536eba67d7a68ae700526bcbe4effa2890fa902766e299fa2cfc996fd58344dbcb9116aab934f985a10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heda0f458704f6cd08b06385be9635ec1881ddbeb977aac081cb4b936173c063a29d459ae37db9f8ab518b17cfd2a00dc5299e32bc4647628ad8f987afd3204c8030d4b0f79dc7ebebf42c155c4a6ce4e5c1990a57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8345a201f35130e0687cd61f48749d7d1a37c52aeeff765da60f8d09e2d215585df8689f80da55e7fdba755e82f174b2e51cd3b37ed40a8b422edab0e5c1f10d4a9c2b7ac454d618631f110cddb6a1c1c4dc876ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff3b955a134dc5fad045c0e2b75b2e7135e0f14873c997c9dba68e1b574ac2d3862053a9384a0ab47965a6a0f8114b8b7fb184ad4334bac8ffe10cf36269b323f40381bde6d55b660349dfe3b70115cb6a285b9af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc41e5fca8d9232b9427bd913bbe9ca021da11802c9efa44a59d11934b1701a7dd1e118205407292a4655554fc11aee631b63a4570264e7210a020f83fe60f386dcae929218bfb7b17fb37af7cdc25a219a888628;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6bc465dabec6283066e1e0fc8f8ad463f1579c3db9152e3900dd61d7ba0fc0273a5f7cf096f12e6a49e6c1cbe79208d01c441ec9bbac748b5b2616429e15869ebec12862540159658279d9e50b8196abebd59316;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hceccb5bc0a254ebca599c45c83747f36361428733ad22dddb73221735716fb0d49a80c5d5ab2a20aa1233d9064ae9370c54ea7b0abfb5718c85cddd99d96a6de9dc5990486c4520482dcf0111ebee9745af015f91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7beb7920426ac059daaf494b857cec882c15cee0b55bc2dd5a02e2f1db28cc901aa9df469679e75a9464f23d2e2d2a0e42f177ea6dfeabd60bc51e91a1cfb6bc565328e9a3d8355369b0af51206c8505ec494316;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7ab94e350a127aaf1f22e75db29f1cbf230cf3ad07557703f5c5a04d9074f8299c4a395c92bf2748018938b8a0f3b57516200978463d62206b2d05290f44d65e604003ff66403a245dc90e55c65124c271bb292d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he51591bc536b903caa381b45359f84ac378942d4b03e8ede29404eeb17d225131b308ce42ff4647433af443864816bc8f5fc165c36d4b883b811f004dd964c5b278591b38f9e9ab962dfaf9eb4687eb02238797b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3b8fe102a2ae9cf1f2e95463b32a6c65dba020e4f8a076a77e7c434939362e5d47e024ec97857648e692149d5fd3e0462b80f6a7bbf07501d2111d1d4e210e098517df9a93c8eab394a5369b22bceec300a394ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cc976fcb572571eb6b4c01836c938cee1158d1b3656ab0dec9dbfe006d383b18b9a561b2953972e8cf726d03495495f64c9501d10d9dd5c54d99fafe1cb148eda18e9f302bd20d536ba2868d450be5077801ed4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d910cd5d40e10b8f735cfb60d4ed35ff4a4654b3b16a949c1356be62bae856013880b05d8967596fa5ba1e5d19a7aeb3db73fca595a8916889d74f9dd9d29784bfd6a944495aeed992e09fddc9ff309ca70e5f16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c1347458ccd9b8a83a8c311a835e404972dce6f7813bc560226b7885443d4c5e35892a33e915ddfeb72c04a169b7b31fe86628eb3d18637e71f0126d8a20262d3efee2fa5b1c7e9c5db58521f518fc769482ba0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h421942d35a96bafcae78be3d263989d4b455dda2b627fb74822ac468f39f867b59c792d981cfeb9b95a5b94fe97b3f692195b4f034e553d9d3fdd5d9d50f16b4024cc4c7cc60c6d44c584c8cd9dc8d98814fabb25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3939f3ea293a8ea0de6fac54592d6b27e4c879b8f675d21c181478aee9da5d2eb22692b7ba3416724d64d404e16e47201ca88467ce8df483eff11ebf96288799bfcd54638d0c0aa2651678c553a14f8c717ecddc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha75758c6686c60a45454416901a295235077bd9fdfca3cbd819b857028604cdf90ea6ae9ce6fccee6bd58bd4a32930b4f0b0459b2d025cbdb58bfef920a4c879a00b3b6df6457b3b114cb1d88d8720ab2c02986a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha70d7b913d823cbcd421e5866979d3d3bd91c40b6e451e0df6b1fe6393598b71b1ddc1867be37262aa96040664f42c3c42ec3f1e05a3a872863184018d68f0bdd4ce305424675bcb4f8db7e0d86c0a71086526c4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h220ef7284c8c65f4d4d3d8df302b79e6b2146bd27693e5983bb62302367058723b8ca7d6be734904b7522fe5c2b94d981047ecc8e7aa5b6d58bf9523a28e6483a042b8a0b8dd854651d9cf5c4edaf4b66c5172558;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e646d1bf8906fcf73f61a0db531276f0eca283802a5ffbeab85a270e6c65662a68894668aedfdf39458d32c61edc2d9d807d87f513d844835e741b6dd461663ef572bb5268bbd4205f88faa6de1056e8860751cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b893c4717c8ce95b81d16ac8a65f080d6d20e09f4a0d620649aab54a710f58e26548028d4971ec3af6badaa604ff6daf13fef6179ec92cbdb20ada74b240ed1b462cee111c0cf9efc0d94a465dbada4f423f872a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee413ce0023bd21d33b2e34127bf313f44b4a62fceea0f5021930486ad6f05c84e8394b7bb749857f37b214bea23499744d740f2b83d3d8badc05de06adfb631cf0b8ddc8702c4ffbd526b7fd2ac546e2286d77cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a28f86d678b68bfe51c5fc4236b71d4f9e6760d4a8689fa979f5ff650aa15fb378223bbf352824d6fa2411897f626ff347affd7de2455be0562cef73fcbf6d1dee0e5b0cf95d2e4622e27f19db70aec8d161f224;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa1655ef4c3688d4df0be18bebb038760fa7b9f195d7aaa9ba1760f51a2d14353ecd32212198bdbfe7298a4ca8a76fa334f34449ba0c309906c982849f319977107262afd4d37295472a8585f0835783ce6bf4e52;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he35fa1823a8411c89170aae4e00cc6707f09ebb36bfc9bb40eb7c040f692757b5b4f0d8bf2bb19a5513377056c4fc88ce1a9a799e139d715e23ef9d8865dec8a0a4799ce03fe0f14519654976110dc23bcee54164;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf70b66d88507398a0f05fb8abfaac711df5be5c53aaf6fd8c16746c0f006df8cbc19f1cd5c21defad69945289f72055f6987b6443c7c17aa661a963340fff34aba3cf40c27f1c08f788ffd0960ed7f5d8717b319d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe96777f772f62289c4b335b9c113b1f181d1eab31bfdad2091643ead97aa32a7581c69d9d582293f94cd94badd542baa89980ff2d63d6beb7d7f279d48f045d678c7ac8ab93a2c30ef4146b935a7890afb3d293b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fc7e32029fe927058f7a20f9bda03a4756181040d6c92d67b9fb4134b32ca130a39c823bcc9781a461c6a16b1aef91d94af0c85bc679e2ccc20eb10b71932432002883745b26daa07b152a909474b3eaf769f648;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37f1037335ed6aa1fd2ccdc5ad3b59d355d0bc73cf5ec2b8e549b429b520e220493fce9055782009468a0ad64f11c4259a4198d728b32b50fafd90a3253dda55b13948b11a7c22778ff3e395186d3e924bf506355;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9211fd23dab14e3efb386d22ef6cd08b76e1db80729ec682b23a8858f5a741e6762c2ad1007277cdc9b8dfe236e653ee585b8448ebef5ee720a4a83e917c1f3fa0bf5f14b2763da9764b9a45d2e740a9356f5243c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7b09b6fa73f058f8c4d02287a3db00383ff5c837765461785e61c295c6206d9d3bee7bd52a5a7f943b1d25a29b4d2e2e6ffa7d03c068f579e961c41e8a635efd19e93d86b7f02d7c64cd119eeb8c58dbb09409a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30a6bfa0829ece84ea56fcb5b52665ceaaf01767007b3949ac3c0582e677d88888821d84d239109363c4eb7deee5efe3afcc8b145fcc75ec23e4a58ced40ae511101a57934685b9a3e608fe98c7e72721a0435324;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc04c978aa64726e60be4f301bbb9b5e3dff2208eb5e1b584ba02e88f8f561c2d549d8e4fa2239fa5914f13638695fdd645d2626ac815ba67c4eed4561e29ed0a7b82153d4b1b1ef15d5b512c177cf274b64c6d70c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb881f45234c6b9c667717e04ca2cf54da26c87f94cb91b603ae51363114411fadde1be0cb58d5743abbc0072b9996c7bf5dfcde2d9c5423d95e371c81b5278783ec7259fefd564382f449f4e610f1ac87ab99b3a7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb25eae075bda5abe7483aeca4d193e41d7a004debcf2e25e11c9561ae9c089b90052f1b63cb37b7a37103f74efd817f1cbfdb00b28ddd4841d17444ff7b53ac62e2dfed2d80dfe8f283fe774f93161659f2e19a0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h486b8be5fe203c18f6b9837710e1dae827b8551bf9aa6d842a45fdf1551d9741d0a2a4ee0d6438790da1418b15a2c9678078693b406a592301d546d4df3b92e54b3b6643e747ed2c92ea0e5e26f1638d1034e33eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc897de31c84a4192cde0191933aa799ff9beec79912b86b29bdaedd3bf23481f8028a420adb13f35978b110e52527dba3c24b67152241e8b6ccc735d206f1095ebc3725cbc201f3685399fc348660140b395e97c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha97d8940ffe698e2feefb9b0511f4bc721e05be7c4350a1ed124ceb7b4ff41bbb26576a6df97391be6c54549785a266cad1dc8f19d34fddf13fd2521dad4d5ffda5f541eb57928bc09e48250aebf263b1384d78e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h444d302090a4e52d46921a4c9a9f28cbf9c4c74d086207d06c24f38de91a62d63a24bc951aee7fef7d387e09b6ec35fbd78a2030c8cdda63001fb21b944d5451551b7dbad47b92439f4a49293921d2f0e5124d637;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e3479ca0519db4ddc2a00e6ed150ac68ed54cc9332145dae5f85442e490a535ec870ac5669d56f5ab4289d130682aeb3fd9a2fdf3c8b307204b295e54541d4a629f668ab221f2d07ff1afe22acc630b68f454f66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5653f63a7860da2ddd70fd079cd6d17c9c3625fed57af4884b9fca6c72c8980d8f44e9e7f026372b15db22ab7bf5d321bc566074c0dd4164d99fd2f5674718f12fb6e13b08e99e3e1368b1db917b9af85334ce0bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he33662061ff71c65f008fea05e98ae1d5b16e38d9a17abe5afd0d58655fea47664f021dc73674ebb36b0328cb63e998990df888609356f5dfb01f5931973278084bae349da7137674fb226c80e8c2ededd4a39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h572df07fd30119d3d9f7f9ab039b84c5dc4fd6b0a81aa1a785c503debe92f48868992e8dbddc5c9d2e7b3080c7450500a085da3c5bc5042b12d67b57cdfe55d7ec362c62f5c533fc4dcd0255745f062e5f0ce57ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5f82d22b292843d222365e196f67f48f2af62945ce7e02cbffa264990f97b1c0a0ef263d2c98ec5805ca816ffc031354dc30b0e9592cb0e40c3458b100dc47dcc5988d58ac09b29f426ecf581df2334e56fc8a1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h167b91bae2ff24c61e98d4065aa12120c2c42d623e27ddecc40898f547238d3eafaf838a547ebeb8ddc71228b47e933563dcf39e6354f9cab80dad6dcd0bce17e798da1c0352cfd841b415321b1128aed83d3b92d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2c223e7489abdb4011229aca575c25c7a81eb8929e5c5030a2062365e4efafffe51b0a018359c65351fa9c8c98f719b9db7ff8a13a1f7dfca131ab540723a8398a46de71a53833c14a32470099fa13601b20c0d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0a525dbb9e5f85803c58cf8340b0cefe9c26eb998b10ef018012078f29fc0d3b1850b410245d9a24a386600b1cfbe078cc3855be262bc8e4a545a14b738163eec92b2d677be5a9d3afe31b2d89e56ef26b2a0dc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ddde196e764c472bbcc06837394cae570dc4d64c020353fd1aeab1014cae498acdbca810571722dcb8305df5819581a4c77d53ff12aebcbd191c2d79ec01efd4c05c5f679eb3fefe6072ee8e85457dcdc3b18ee0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd8e6b9d3df53b47ae9ca452c85fbd51f6bd879b060c345ccf503426da91c2f599e6015fc38753abf4990a08250bcc7880dd36354319d47fbaa3fa03b023dae36ff89903732ed736dfd3437e8e5e9fe34acbad36e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb52bb8f080f5350a568936230c76fc814dd1220b75af703ad2b85cf0ecc5b9bf4604c04165e560df7820f1e3a0bbc718689dfbdbb4336e8bcaad3f9dd655615529066177f4bdd97c5c3138784920d20e18969b1c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79b2d239872b5b7682db504615e1ac9157367904f004e868980c7894aec3dde24d972c346f6f745ff31cab62ac0df2aef29f7758f65a49571a67f01b7591d9c822cc45faffc76eba51ca1bab682446651e9d4dc17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe1d526438209c0a550f27e3704a399805371d7dab2939a632570bbef117b831a7920ff2e4f9009aed6c786007a9cdd4dae577f0a3b55b2eb409372e33c3f2fb26cdf9d509f079659eab6588d44678487b81a5b73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b6d90908a62a47936e492f2fb96b24dd7837fdf76773402687e5cc4d7659db74011c16f1cfc3983e4f7ae8490369f0e61c2ec0c0ebc5d1fcb6786fd0b30b4216cbc7b225f4562fb21227ea959568e44ad5e4817d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd11b8bc64ef937f0bad9d2aa9d11cd3b0b639072f8d637ca2b81e18f4c204247751bd05dc641cdc8dac883865109eaaf34085af8658c8f4e7a446f958d1a487217bd9fa2fccf4a246f5d795ea219e7a8e1b06a57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5dd43fa3c9a1e652746f5d88869b88dd2e70b79e262b6837d806ac68af30ab58f3fbb9c92977012515ffdb544ae885059a68d61c216bc2da93f003c646496a6068babd7e90e509fac42cf09caefc49d984d884632;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78ee8f26fc5831f9317ea76506a0c2ec48a7082acce9460cce37817d6d119084d5b83c5ed32c7f7375962e6203b96e47fabd3c93c94805a5b8b9112f440e461840bfbf3e0f7862ed8d97464258446020a2d322c3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84b631b657bda784a5540ecf4d76046fe54663e30f43023943be96f27e4e9636f66f419b3c04c74afe279cff84cd91cc28238cf59b82a5072a58c1d8434e15a199d1d2bfad62185eb114545aad04acb01ecc32a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h921a51fff2e20ee61b9305761f75e3fc17c2b52867a80b7f095e2570a8d1c76263a2426a6ac60c2c4e6d0b68d85c7072f9156b3835286f3a5d1d767006057c3cb2cbc3cd2bc43ede2a311ac27e9e076f7fa439a05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3e65c4e733688fbe0893f62d1c9046e7e47ff8f767620155942c5c51e7d8d40a572a6a063730ec6a97edf66ab8aeceb926f3447fbc4471a2fa9a6ac4c0284c15eb78e881f37881a74140af8636460fb5d21e39bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha575e29383ee6c1ff90186984861f40a694189ac0dbbc879ec6c58ec4769ed81300e24c334680588b27f14df0e6e403bf6a03034058857dbbab09595889c6d22ab27a68b68b754186094a146e7b22ed23336db998;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcff99047a917f5fa68a191019341ef125f53b32d494d0b8bb25a11f2b9eb312ad4f6a0cce860f47c8eab8c17e24cacc4d1afecf2e9d782bd438409a37c6ec227cc2f23a72a58c0aa4aebb4e79a9efa568b9d1c05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6859f33edb0cd2d2fff7d1eef18a0c9c0ee56d1f76c17f615944b1189f56fce8d24ed4ffbc722fcc671c3b707c9d28f876b06f901a85c1c31653baec41dcdae400daaa70f62162ee913651a86dec5c4b5b6fec8a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1808dda8e12072b63ee51865285d272deea0c54a5e20eb025df79a8bb0d0cdfae82d71cfb1b0a20e2ae9b6bd56a5bdd1ba46226b4191fe436e2cc8cb5070894cf89d2cb07e7148064219dee258f7d1b1935086eb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ed391022928c8dc2b4584bf0d0e1595606a92be63501bbfb61b7c19b26694ba3ebc2da1c1adbe3d02d9f6981b4cd6a66bc84c76b2ef6c155130b2be91b78260c89f37c06d3f508eb4d3830442c3408f21149ebe6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90b897b4e924f6045416ed88d13c8576bdfacfc05142f3c51016626bfa1cf8c3a6b3880954e1f5ea54abd7c031a95ff82b915d21c5ac63278957f3c990682025bc86622b150b19ca58157e0b4fc5d6350ebc2f42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d1abc75d5cd7fcabadf02ddc838ae48fbdaa384f57edf942060ebcdafe40a0843e6c73382d010b0fab92acaacf363f556732b92f5ab9e6169beee11429ad551993ddb6ee0e62edb31f121c6abed3b42974cf8814;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cc501e64f5e372eded038154b01ba440cc41d7e0415fbd39318e70d40bf916391bf224aaa091b901532a5c6ac6a48ea259874fb0f5961bdcea2d2bef40f5b91ba4e53f1584708100402656e00506732d1792c4f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a34a3a12ffcd90af7e03fbd597dce96d2cb02ef150db6d34b04e3653fb70a2a9d7227e98adc92495b13d5b30bc0060b07349ffc4ebdbfcf1b158c986d74cb68aecd669ea6dda0a677d498de4f30d2b159679ad07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6f5318115a9f2efab5ff1ab8c585b12312dd5b50a8008b0699785d401101da0b08c978924726861be8fcdc980c914b2d5e570adfcc3cd730144baac8a8dbaa8934e9d1f299bdec6d7e9fd982d2c9144d42242da7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e74705d198ef2b3842c917149868a1f5e678e530c97a3f6258335896af431636640b2c9261f5516f853dc39a94c7f9e68caf3be90a964df7ff67d697718fc642377e31045b143122da6051d3d5b51fa79e6c6e90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h827644e52ab8bcfb854fca21a799a73608e432da2b91a517b8a9f37af478a02120677137b1fd9f1dc993102a9d82eda2b837f22e01ed7bdb971588190cf40d6811d4942f67af3dc642b3f8dd4eb03ca926926382;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd059c6b94a192abc55319a2588755ff43cc5867769915b8afce2d7c6caa1e56fd8163d582dc3fadcdaed5e538750097b1048006beee1671055aecd4664f0efcd0fa36e042ffcc88bee5570e6de840c3599eca4a41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bf4c9292a96177476758fff918beb7f531a64657791afabeaab267acf5196db7cd15cfce6f12660dce5f781dab77dc2ce7400c638a1490da618e15e06a4c2e1c2f2de8638c9d235e3fc1c321d79fcc7572398309;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25be713f04033d33877b7c57b07ac7fa5a80fec03e981043ff42e527df41bcf22450de59d0556ccdab8f5ab9449fefde4d5c89e648d2d3eeabefc4d394c94272979743a58944f0c0aaa6bcb7e368493d641da3bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72cd2c5c1753c31517ab2fa1260438cbd25398544aabe085b659ac63116c3c8f92f174ddaa3e6c378225b7ad082a0cae6b7b088bcf903fb51e3c5f71a8f8b30d5a9deaf0d24ca9f410e31740fbc22557ff51bb6d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f20ee6ca2bfb5bc5e7b87d1f3899d39dce26f2a0abce4c2f991aae05b644e9a4d894ecda2a3f3da67bb5c5685baec508d02ce66055f0b88350d30341309a51b8ae07869631d29b6de94be68824d22d700e3aa336;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dd698a9389d98fc5273cc327ee82796ff08ef134b25bd4371ff0f5336d424ab77979066e9e8fd715c97c0f9c330f58704134f87266b26193260d618a588145b32f5b0ad9c42a95b7276240caed2528871caa65c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h217781770c742d01853467705f138f5a7c34523b73c38f24945d455d2d6dec63dcad29fe62fde4f6369de14086bbee4df229328bdc250b0a5a0aa66b660e8c4d5370689e614ca5ccd8a0d17bc97c21a965f641f6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde33b66d10be81f41f737b9aa90cecaa5fc6ec3c20310510a38188e8f4a1ef44a51fe378a38619c021fc767c299031bfb607b84bbd1457c92ab7c7baffaa1af4f4f28739ebd5687b6f1d3d5e7b1bb75b662eafe83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8e6fd74a4b68def7f709285074ac84ffe3e52b6234a3c149145b209e4ccd313fd8c23df06ca21ecf7f99ce30b00bd30a93e7debeec28b15cd34766b5bb610075c668251ec3e6ae6de3d2633a5f096e3821ad5d36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda197bc4535680d5abeea7faa81ac259a77a54bc946e43af38a1c2bdcb419b84d46df40247dbf2f018588aaec47b6745ca995eb54838e839b8d5ab965ae8e9ab26a9a41477c4e643b7b0c051b45fa75c7a4cd5a56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha577700ed74266cba959f27946770b57cca0e356eb91608c796000d5c8fd1b1095bd1f44f06adba50312ab0f6f0637aeff159af1ce9eec3684d6bcd8cda9ac5402f243538373af49f892e16ccd6a6ba62dd72c27e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b32d9fd483e48cd7a7eb4f51d17655469dc23e08a91b5b3bab9cf12167cf6f3dd47a4282e8be535cd96af7d2bdf8830682576f3cdf95fb88aaf74c1025fe3951cc132f94ceb65e1697ce2c94533a1d3fb8afbf23;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd03df2244a539b16b9a5034523936dd5bee013b5047986998f1399f60c6b4ff0f341a2639d46b24979f82e9eda18ee3e976f4c69b12f55e809c2c40e7d3a015829ac0054b3f2d8b78bf1a45f6f104ac46882de3d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb620a1d1eb3327489bedf3f5b0cde8defa8b581fc2a6aec524613912c583ffb7dc61a0a4add173a86951312a4fefac2f95d895ec62969eb3375c3158c5b24a58ce706a1c9a730aa1d32f58d65f07668efcf600b16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h134581c2f2083a5b8ceac5c50d9beb05a4012a1ceebd11557e2e4753a2480f93761c09ade8777ea6776819fa50363eb9e5d2e973e9e79ab9e38dec4a1475653ef8981c4f34fe6e8e2ae97db60cb8b5444c63e760f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcc77b50b03a9b2db8d14ecb90b0ff0768bb3ea9130315983adc5af5f58ad8c5b2c1dc329ae0534a739d9117ff98f40d3917f1a1281d27e7fd87cc3e9191ca4a8ada13f43bf79803ffdb4ce79aecd3013d2c89289;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h657130a2862d8e0eb8936d49332391c9f6d2d6bc997f9f7ac3643e0eed526148b8c71e613b577b08cd8137714d8904c2c6ffc204e726319e4c68d384b709c73aefb0020c6402f1accc5b0cdb984368afb837290a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff93861076212a8b309c9f4b2cc5e9a1bc862c8b9b8ae6fe2b32cd4b882b3abf5d05decb14b94e1e7bb18d1bb1798478a313a157d76c78739e784b63329a1e23939f9cd146690f5d3b451580f8ee39d2ca3e68d80;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29b1bb07dd7afe1300a41ba83273dc61beb14a6f3ca744e44f86c269472db084e416cdf94863e294ac0580c1712ad5bd4d81ecfcbe5a7d662b88675012fa3949f666993e7b89731ee74c3e58dd74767eed0e3981e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e7461f5081b577d0e65786d5c4763d321fdba4916d46d75fb3c8e033e7d930e97b8c97df24560e46e211c9e4bd257cffefe45639d76ae5e7f108242e022608010d3a223054f17066c99cad6494b0b3751bb4f327;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfe8f80ee7c4a384a866fccbc93d7df3b056cdb2c95cf21ba90cea30cee2207e4fdfc360ab07579c562b3cc7b3e63f0f9f3f48c302420e79dc440691c6fde8908f581eccbfa65f6e480640146045f52292aeb6566;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a862141245a7595f92183b32f9056f6921f4d0542c8a6cb0684c55c7147864ac55285aac0dd5f61906e9f14589dbb36b98b110a2596599d746d782e554fd596254b27ce9b74c7c10db3bc7afeb3e5698ae9b026b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a04ec9c83174fafb45f5e87f4f0dd6d437a7f01c534ca5c5ba022a810957d4a5f548e0f8deb71c3bb269a7dae5b817e431d7048f22f3dbc24fed5ca92629b121633d6831f4b91faf783a39d1811ca0d0aa0cd3ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc494bbad97ddea5109805bcfc7ff56ac089ade12587c1e691be6d044e0eda04c9d4241099ca27a9c0194218ccd8b2c088f951b515f1d1dbe0d3790e456de555f246479ec8f781b37a49b08d90babfcb4a48b510a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e3c96bb253f024c9c863e677d224c419f40cbcfa6885f37d034be3fba98cc6ffadb2501211e975286bd8a71f06d45906c7898989df8498cfddba23b0c9722fbc9abdeb0d1130800c403f25ca30dab71528b51853;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e20258455f0370f24152b14cc2e3b3199780df0f63e2621a79eb5cf4413a8cbc21ee911cab9995529f7f7ef4024dea71c7389ff5124dca06dfcf1238efec46a68e61d18965190d20682dbf7d2bae738c47f75011;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b2068e9dc70f15fc20dc9f468414d179bb7f90b643d30c74ae46b58cb6d4bbaaf068f0769fb4a58d67ba2432b814442defb77d2ace791a85ba5fc80dcaca1f699048183d073383c13f38f5ff38528c8bd76eb4c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he74dda9b68b30a97cd3f67b81d0b484ca1e6c2a726136ad6ba3a9d15c06ab6f86ce966549a0cb384b4d7cba17144fb6a93b62558f2954b0dc882aae06e3f8c194d52bec1b7157b6dcaf539406c06f86bfaf701c58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ad2182c866fea8f33241246e72cfa14a45b9e5cefe38faa6536f4f51832403ac96156085ed8bd2d11d2530608f5cb0e4e2cbaedc31500dd2f44d808f660ad20f0b7f5ab026797f91452514a14d0bb172f0f93674;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4284676f8df423c9df72ad3e36ff5ecc398ba8cc794cbe2a04dc6eb45a23a14c90e984df3015a159516cdcc25a9d56c12376cb263b4fc0a0a11b23cae70e0d4543a781d26b45bfac88656682fe8e698f0a7cf69bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h531427536e85f9457a3e9319c996bc68ecc68b66f3ce12233334c2932c3376dac50fbdd4d564e1e52ccc4f7281aea50101aeefe1141ed3cc755f41fdbac7a2fafcea0d70a8e9410a09bd985814005206e031bbbb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h864c630eb42bf0a8f9dac027745eaacd9ca88300d18e0f99bac66ef7b45b3c8538607fe11ce351a56a5727cd0b17537481d6a5646d1b3107fc7736a0ebc5a4566ab7712070e3b87a9788c16bb98b4297d246ef937;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4993301bff49ae1d00106bb208a111da6aac178ae16f42323081f1311b7c3f803c93cdffc5f534787a51ce0b188540669c82b9f967629b26c1818a806f538ab7dd2d7cfa07b93245ae374c27d16e9b2dd18f5543f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b67af5ce9573459787e0f1ea4add50f6a05e49d276e64b08226d25579e6c1b4edbde7de642b7e4cbac618bfdcfa57d252d0939391ce2ef2f9f74691938edad91d05de2a7eac2567d6d5aa1cac0b08466bd6bb23c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1675a8e09fc66944da4fda6d3ae98a0f3c72c33bbb579df6c2bf32b3e0abe83244227e1648edb6597cb8ee0357d399010584454771b458e93f26c784f50c7b0e9c0726fdc627d449877c17d710bb6b775d76f8a14;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91f160f84eaeea83928a5688397f54cdbaabd7ddace231f995ee475d219a2fed52041e4385b28484dc3e8d44006e26743d1153ca936ca92d0bc5ff8635e96dc1e63d8462cc88821db2abc42f0d00d6647156b882b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h659405950bead289924e005e9fa1a893baebea876a9a157bc92fce8c02a251e22b6ed0fb931a34cb1a520d3db6e32b35dd09aa971008c8a41f6464f393bb1680f24c4dba35fd26c4891f9243e232f1ca3fcdf903c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a6aa6e87aece1f1d0ef3c0ba4ef64289af5c7431a430d50b01d4af2d375f60f3e77222f8da1e2d08d6a762c860aaecbb11e22a7d1919e183dc41f319a2c17056094bd0831b6023336fb5ecfafac4c1c7d4f369cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b464baa779e8d7a81c0dd21408d6e84f3f39ff7ca7ab9ce145fbfe99c1d80cd84159ec720900d65b9444e8001460a6cdd717bb37e19fb59ef51f0a878fea8ac18fc01275b03f1d06c26f618caee625310cf81e69;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1892e7be1bf0efd26eb9b21c53eb76cc2d533626d61ccdc62d08a78a31da7c3923b79ebe2101409dd160b479ca4263088e61ca02ec2b7e6d26067bf60c414da1c59c6912a16e1f4bc861e322382d8bc4cf9db3ae4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb519175149f0f476c7132dd664c954dd4534c26e4bf852eb84ccd4ec5195e03e70f1cd75e0c3110b4d8a9b71b71e20c8b2fd81b7f5f8efd67cdbc496a142e7891ef34b430363db2fceea06b5571a11d711bf0f075;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb2370f7be459eeb8512b179afecf8265a360393c26baf6194b8e5e3e302ff2f25b0639d122e80847c10f4e2e86b7412bc8f1a8a1a3957464ab1b1857a57ab7f7da17fa2fd35a01c21f164ceb06fc40e7e9a06368;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h905d549dddfff1b9f528bc5461b397a4c5d3c294d561ecada53345de27f95eb63db462fc890b147aeb21b1f2fb134ea4f3ea6ed2bf9840acb249eec386807752147a9d2e256484108a9031a0e1a6db193ba5d757a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a5325328c6e26c8cf15925bfa04ab96f93b56461aeb004582179a73833a5a98cbe3a0b40882412056765576a574344c88254a53b1d13790b3f16e31306df21adc451590dab90961f99148e73dcbe7db529d44de9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe9144e18435165e0ad0d6158ce435eab2f10514295cb7a7aed92a8cf49df4014b9501aff3c422103b54b88d01e295802faae3ef7d6c31f712949ae5a8ee638b76d6076fc8db218452a25d80ada2c876fb1652a84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf960623fa7607c19a57efba08833373098259615a5b03b5e742b1aa6da0687e5c35477182d8787c27ae49db7d275580e21162097c2d7a2d6cfa18147c596ed2750c831dc768218d1619cb754405f57bbeed68f4df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0de64d56e241a26c0b1acc419d52a2e697f551e15b5b103b744cf07c6dd051d63ea2cd56086554e9bdf4b20a6f68202eab49a7a22fc03f92183fd78ddfe6148704a91417bfc58650d43f5dc96972edf7a98fb5fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40d9029379157e2a6daebaa6a1917d3762e418190a3efdee77ee58be712975241e26d3837173cefeed3dd15eb62f2d5557bcd8b8738599c719e214d51116f2dea75c88ea3ad712443a035e1a515bc0e66233ed59c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a43412d115a73d92ab284e8e3310e288b65a7106808956f7b97fda94ed1f559f1ef2bce79ec6c6a5c2da96baaaa24379e26402a3289c238fd72d2e6010084346f2a2fda8d60dabfd2f8d36443104a60b812ca65b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc93ee1cd613f11b497854c95a65ddabff35d76b0ec555ed20fb1274f77e3e4fe50007a1756d67dff6e2077b5a079a4e5746a404079c4cf78f24028879c3b465d8c710614cdfd599ae54ae6717d14c085021005430;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82807cc148e65e807af498737dfa46021b9f3a5131ad630d5935cf4eb06a76f3606a09322bb020b5a08a60e0d8a330aa325bbe187dc610c4cac1c99a3a3edad61784dece6f5dd8c6a0d089a2221adee8abd95502d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92d71563082b1c8feecda92bcc0e7dcad89a43d38b8255399d673972c9316cd146d486629b1a9f5d549f3a2449f66f9e8e6c509d74c3e4bb982cc58d666ac88c175d037cdf9a566f9699b3e0eb333a30ed186b901;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96e76ac9dea4d4a70e609c75ebe8a7c5e0976ef61f83c742ee1764d78852a656a050835a8c84f25e28e36c30236f17834a73d09c0cfaa06b27f1d779c868d5ff053d1bd032afc1c8c2955c8f05b50e3f309535322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81a4f4c34ff205c808f80fe40e9692e8fc7044d53f6ad5d21fa00de43b82ce8e3f111f956e5ada6ffb02fdf20c9703fd32aa21686e3f32944784775c4364b12341e20c7527b7a42014f7615c6ff19d7168a01c1d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc259608ceec6b8ef23da49d8fe54947c71204864b684b473390d0c1d7ff12761490e5c94d85f27c3b504d47674a942f702476b537c5058ff6c10d778f7c922ef80ca46a898424d2021a368852a5dbbbde35c1c1aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4359b9c6b8492f73cd9798a8a64ea13a7b4f27b1b4a461973b2f4b54b071471251571c07c1ce3ddac259a27077920cc2afab0fa7676dd25ce5df85ac23c5f2793d45ef100e5c919bec037f88a6dad588bc3bc3a84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89111332865560ef90295abf69323307f854866aadc5ed6ac8d177845c24be70b3b808e4667cf0427667b2dc567ba881d44963953e99711cc9c267a2fdcf4d2e23bc6439dda6f8524ef4769cadddb225c80c07bb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ea391076049a5bc047f436993ac197ae3a7bbae6cb6ecf996ae67ba385c05569a37c0cc127db6ff6559ca02d1130f3d7fe03fb22e124c7720634d01ece042ab852a78cc9bacd626893ead550692a13820def38a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9743a2251dcff641b441b84040715dd109c01bbcd00d47b1041cdd9d89567fdf2bb2eec96001c5484235f272ca5e6257f6a92d2654e518c600d7782af7c69d23a08a26146e6407dd15ecceb504db33068ee62320e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25e3dd0f791c67ea96e1ea9efe041877ee598099022b4d6ebbcea6eb56a8c630aba8f1a49751413f3020ede022ff6aa7af70cfabd2975babfd3f1f6f5b837e58c391a72a96ff22ab60a42037377695b350c61cc48;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ff2d8ab690c587e840347eefcc880e59d675e31ae5b547d252116a09ffbd2b797527a8a1808e03bcbb0eabf5db6e7c5766e06676f01abc29556a587b903567bb97d31994a8c8dadfce98bbf098045bdc132a51ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3565e989e7d7dcb1520bfebce8e85566122f8e197d27ec513eff347b2a7ed4947088dfc11077d94256fed3b6f8558cbfd8357e2f429a8dae7abe6b0719c03d7d0a88dfc512b2a4c98ccd1785fe160ee9dce240452;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef618fb46899a3e1c58f4952d3615ed3f243d95fd21a64ee64d2109e1eafdefbc0c72e7a4079caa95ce835ad325d9b2a70ade8382a4bf7206fc7a860648d3698d6e770748144032fdcbcac0cd8effa47e73a17a10;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd595e1956538b1df2f8d1b498f861ec71cba616a96e14a94b10a0f879cb6632f7bd5553fce618467d2f8f24ccc3bbe7162e25f8ff99572295d2db5079d2f171e33cba92d5cd87777b708fbb4cd5c75a2ac7946782;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7bb52dcfd273b9d4b06f174bbee09a35dedbfe998057a64463791716758db8952c15caa4f8d86eb724bd72f2e4f2444240e67c35a69608143cadeb5feeb6f75fe4f60ba6be54370cbd5615bbfc3012b302c5ae75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65140bd9040e153428f08bcb1ce50a7a2f01ffc0544ffa2b48d19322f1b72e7a644bf383524dae0c2359edc58ff5b0801defa7eb572cf303f0193dc05aba721f8ef724bca1f800fa5bb31e4c2fc794e666eb3cda9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h320cac7c25c9d8412704a49244b4468f9f94c5775d3ba6dc6815ade35e9e58ec9e3b8b6438055b295f6855217e0d5a77949af1460a23fa0c7f47dc72cf3338d7b56a476e9ba46c05943898c2ba47227c39b44dc1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79e7203bf14813d729e7b3adfa4f15927c182c43d0b5ccb072831c76d5448b186fc75ee38c9ecd3166ec3ddf9fc5a835e9267b2cc222bbafbea1c2664c763513ae4d0429953e5086c27a2041508d76ed8fc054d47;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h127ca3558d92991103822583aa15c23526a833a3d07d009e4de80a2a91ce55c154a95b9facdf7d94d189bd56aebe68ebb0f1cd3ea2fc54e223f2849f3c48292b2d90b5ef6da13baf878678613e04a069b25b5fe2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40236fcb1dfaaee35c512009bd47172269326b87399ccc28adfd44252d2a5f9fcc84ef14edb730f36f5b9b76390378067e3f0bdfc25afc7b0bf26f2894e1fbfd293122a9641244091721d53730d8d7dab2fd1e608;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0ab11d0ff67e3acf2ba0d5ea24cc6a3b55ffce68db4bb427c879cd48cf7ff7d33e50bc289d1211a0194180b03c7335366b32f775078545e93da186668336277a53690b8ff0423ca19ced749f9ccf5786c1993446;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17b916f98f324126280c9f166ba52688b4209d18b212d6501dd615e5798563bd7dd52a1cd1d812fee3aaed096821eefd6d334e8fdf2b72b3005744ba16ebf20b2baf0a5d674051046a0a6c23c402df1657b4f994;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19afc1a5dfa91e1d06e1d5a532b871482f1dafb6bc91120534c63c78f339b204b89cfc1486db862cdf89c1d67ab36fd983ce8d72533212db06de3de43ff0869076a5888173ec7d382d4561073c41f1bf555269cc2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe39f03ab8870453db48fc24a3669dee571112539d7c32f80cad3cdc89e88b4fba235d946bd56ab2bd7510a94df9ad272206fe14ee775d4fb9493ac52a3de5421fec7418c00584d74a38c7b94ad6cf644a86bcb58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1890ac91d392093bada36fe239d031777ab21316af3889538f538dd6dec9d4a5e5c0221557ab698e23bd744098011d42e1763c96649f7b65a12b621293818d0fa2ff9da19cb2962dc0743ccd915917fda6bc8b6f6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92cbf3abcc6ec052e8daea2ffc6070642c82eb739cea10ded39e2b935205adca55e5b59d81ea190ef46d0f14e28bb0d652c55373d6f284d6ffe56398b91bf5532c819692b1fe16445122a8cf1cbcb756fa3c753e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f78257eaa0c198a80778afbba86b50857e69f0825c9a5e0b299d8a71543441617bae3718b8013212cf7763b84bb578757b2dcd86ec8a254b0251a59f517899588943cb50efe97db6d0e72de2df4fd891db4bed5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28066f4e02180dff303610b1d667eefb1ce60e75f098a4202d1d66fa51ddbcd4cfcba6f2bd3c561a26025bc9a1f4c987369fb3ad3810e87f3c5a15c1d17dc5a9b805d46ad218b01419bda86ff4dc75d8517929393;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93d0f854898c4cf4f5d4effbad28e8cc5c0b9acd5c02c92a5cbc2317c762538d33d0cf5fb6625c966b409842bf7f7a1327228ec82fd7d363d05e93459b8fe06eb5fb83c54bf12650d1039062025de6151b225e30a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64bade20abf2196487aa44ccdbbbbcc9653495289c34a0aa3261a4a2266fa8e06076a5ff26c58b7321325d4162c516835c4540a5c005b8e5f2a48a9b8579cc838e1fe60ddad7a652870a5200e7d4f840712b700ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87f3d7fd0bd597c955dec79401811df8bfe546bcbeec36631f925696b2c668cdbc27c734eb924efdc3eaeb6fb118201a102e6ab7edfef63b8004eac75d99a0aa0a7bb0e3374fd9cffb9aaf7269764df21ff87a993;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84ec63332df9c20ed239a61c990b8cc48986c72a33303443619e0dea1b3749497ef42c469cb40202ed5bfd5fda63c3ea77aa7c696b9b1472f20c782641deeabf20446277a2379f57e780c3b4a7ed86689d1dcb19b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd968b73d1cc1f54b83708730f609b33cfa1e8b545bc12e7f58e47228915e243ccf96a83f29fc5c1b63654a7554d3f05e048252e428ea97c31c111922629bb63fe6a2c95a41d9f66183022637137058d2571aabf36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1dfcc7f10c14cf30042abdd14a1501cfacea77f70b9eaff4c5a61c42e6d1d82706c9bad5b70596a7934eb01920489d5d8c0e71eb948296291c61c071bc092160a544336c43f1b296787a098653455555a3de98f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51e8388c63240584ab29ae2e9a896646d3a8c6cc939cacad3d46597ad0fd4a78c69b6d87b643ccf85f0d5086df8a9e7f4617bed6ebf1254ab1293e7588ea6b00e81b1145cfd5051cc85084f3c271c5b57b4890921;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9088ff87b868b1ef6a724269feacf524a931df11bced9155d161f0f3162b26fc1fe4976d2917b5fe7ae7427bc05fea7f0754045a9b51389190013aaa78cbb09ae3614da2a345ae4c1d2bbd6e3fa4cdea4a7a5cff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h425381c1603b1b60a9ae8f5155aba119688c0c0baf69e2c109ee192ef9d188f59f627349c7c601032e148d457ec5bcb41bfd50b49dc897404422b6c9db858618a662f25e41cedf60256caaa243f7f731e88757bd4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f1b22bc5484066a17b82a74002f9781b39b3f19eea5b59b20abf5bd285e211420e6b889a53bee40935024a0f86e3373b8ddb4221b33205cd3200f9f687b2a1959b008f2b3d3b4fd8739db9846821c3199b17ed53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82428194aea4a37764ecef3c8d0ddf9872aa3418cf87c763fe38611d0ec5997f96314b16e4a72d366e137d9bf9cbe4526f6f1589ed304d6a791eb8fdbf3306fa3648c87ba7b4f201f787d9b76397f622cdd815da3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaefc9fa2632423a749994253e74022b75565681dd157e157f357952cd3d7978cc304289848c5204226a8228b07bd5ade1bb5750ece841ad2f51117564d042828a51c4afe4262f356b46e5f1bfe3b795fe22bcb32;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d09ef620d35a64152ff5a52ab41fdbc60a400f11166e9a09d3e63b3a21bffe0929ce2b7d25138cb5dba5e9dcf06038042ccb99613aea45f5a773f54c5cc0cb9815f8d8c96dd92045f78008a0b8deca69ef3ef50b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab123d6c3fa2a67948d64dfc02624bc294e53669b20790683df39e8f46b9912bcd325eb02351a38d7af5355d2b526dcf0a0bd413fdea20585770b36c0dcdf7ef06d6a7abb3c2c470f4202524e0c9018254e93f4e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h797c12ad3b1bc520d04acd6728732395dbe85df3b7116460a78b993fb65a73dc4b50f264ca2329bf2ba29993fcce67637f51bf832a89598e6dca6956957ec24397dd0ac21db11f48e40bbeefce20e3dc168f62bf0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b928783ae48994bbdec8f2b051514ea46cb3c9055994ba4750c66d04eabfb6daffaa3ee31fd9e115d1fb8a60f9c4353ef56abfd90bf67aa3a346bb7c292c3c13bd3da8966b1d192dbd701b0cf3189e7d8670c9f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc36fdf621ba016db4dcacc52623851daaadacb09ef55fd0352289e84badebdabf8e7d07daf5b452edec4a942ba7f9e6776ad0324e66d1e103a615b424335ed8af13af9c0b3bf648c2e41546641a98a9c0737300;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19cab8db1f28d5d38761efd2b596091f029ce8fc41010d787d4e0789bb8cabfdd65a6ecc0615d0a7ea786e8e8e45efb3912013d300d8f880b56fdcf1e418c6776ced02472080d9de7957b5e2459135425733ab53d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7c1cec72222a3ccbc11a38313a97435f0962e86b108c57d6733976e3e2013fe40514ceed92a724096a13a7dce395b688622ff06b948d15a2bae76d22202aaf38d17c9a1788e1868336493945b018cf8a24f61ec2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40e0b98108c14912717f5d9b8544a588bd4867ec1b3d615d1dd2e2b3167cd1a8df4abddac805c7e41b6c3a3cfcf7acfc09a33567c8a11971453acb37ff71189d5838194ce9ff458a7752170bdd3e9c8dfabf98394;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb0a44d404a8e10ee7a3730588f1f0d2f1ef472f323d3fb3850d19178f1ee8ec7c1db332a621463edc80bcec5f5c74aa2d5b9f2a45f432955e56171924c6386a620fb17bc77288bbc7f6f4d29c17821cfd59879e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7705f1ad591077db986ab6015bb7d347c7e9be5c5a0e507ed09cca17cbd1a5620ead8bbf3e34d2ded0573efc067379dd205eef9d339094fff59a64c75c1a60216c8b7c695cd8d4e7ae95d665f50d3c3300d22ea8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb325f81a9e63eebc8754e9ba908f5b79053a690282c0797c4daf366e866fab3a2ff1db645b8fb41d4551821e02c11bbfd0b7572c4f07d7b96963cef19093d604205e8ac91cc4ae93eb78eac611b1940845a36239b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a550ffa5c96fbecbf09323dd83ef90c5f40cabc86b856fd3c535c70312ac8f69c453bae3e29862131f1a0461563d1548755d1cbf93a8992bd665243510ac09b9823f336926f0c28e152a7cc82abc9b3f2dfbf55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd79b19d5a93fc3131378bdeb59b612067741524d2ca25abd2f8cf8422eaafd814871fd636711965231b5d29dadf1d06fe4330723c24ca8ea922d411c21011b800efe8d741702f8f32062aa9ac532ba11b2d27731;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbfa9709e22daa757532d20b02709bfe27f03b6e0f1d248c4ab5843af96f663caf3248c1e7ebd9f510a4abab0bb1eaa42f23f9820343e88f2cd1d1cc09616c04d37f1db2af2a2031b29f92dc3d356720d9abdee75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48ffe6dc4541ee994a9b2ec2c9d46c769964665297e1d64e2014b6dd47565f60cb0baa09347e65b9184c21dcdb3ab30d3d4d4b1baadfa5965dda9bbc969e50b11e12509dcaf204184499820aa409def05ca1e97e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8bb7ba858dff27be36a857c313d21c11f74f77831e0bc8c88d135f75bc57c9a13d9fd317095c9a932f04853e12baa2b2492ebc4f43bc256a66a155e810c0df8957779dda5eb665d6ae0281e305823014449fc0dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb0fe1c6edecf2e0b070a508c2e925ae7247acb4d2fb10b5881d02a3311ebd129b25c12e0c09d0e73f413a85ff3dd22b93edff733bc12fa7bcd4ccbd5c8269383bc076fdb111012a4bceabfe2fd1f7d23909e01e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4562112c66454543ae790e949ee4f850413d631ba59fe3a48a28818cc2643fa9658316a88b0a69d4eef1bf69dd51d52f1b6c925d5b9e13123ac3b55a14f8252ce747dbafe5420a8ad41e886a5ac8144696a02a264;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd512787fec59ff519205ecf4c55f8e8f2d1782d140ff5d5bf17178f60f49a13da17c74aadeaa1834176cb05a6cc0a08b649c7069a64429dd1da99e90b6195472269e079312e5ae06771d60bebcfc5783ad88021bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5fcd95faa967a81a580337aad3b65942375f348c0009547521ccc5737479d789334a6299fae8920fc8b7bb6cc392f664dfc83d132e711e36afc7a53e62cf09d1ec7a0871eec7ae79d19b0b4f928f4d46e6b4df91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa25eec3900125391a7aa8a9bea5791062380989fccc34071321f44df6ece7333dfdb15c33a4707f2f7775a64052a7833ccfa5c13485372282ab5189097a57e59f3e067141a3cbeebe8a1a7dc72b66fdf9b8a7b53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0f4cbb699914a0e2c15acd581f62d302916b0ea85231d9bc62ac30ba4a03c37c3f07063d6de4171a5bddc509b171586a9e32a0edd741cb1cf1f2f47e112344cdbf4558b9b55aee054b61712db8915139b25336ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f4dbbb3eefc8180fbea17a00e248fd4f4cdb93e64a7c0e3f4da87400d4ea03f57fd6dfed541162adf2409e38c2b1bd70475212a12b5eb28fee66fa4dc7a18c40f3ce8662e6d0dfe86cb7107fa581e45636a18f8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67bb225acfbcd13ec1954ef30b1de9a86f8ca70c2a8ff4e95b5dacb7d17183db68706c73c2611c132173177cdb419aab49b7c73ba3046a3370434015a4678252e1c2a5ccb935a15c3a64efe6deb3b1632b2eb294f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ccc1530fed0de5995b9f18abccdf64ea7ea1e2781590e624265cdd272ab4fa1814b9a1b4584b0016477714cf58c5a02066b8f380aecef905beb446dbfa87a2947e32f9c2259b42cb11e6f60ce9c1a57261ff653a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha303fea5288793dd4cace7bf38a8ad348b4d504e88df0059d7ceb28e9c345f17c74b61e146972548128a138f8d3e2ec7cd9e192b6eebedff846afedba3f39f71c4e5cda0403081eeaea9622139151ce6ddf514de5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ab783afbd2ca552d5e94c609a78fff47396336aeaa55ec047d1f92ed3ed7b13e183e087453e660b2d96ca847b24d49589f1d8bade4bd5c65feb156ceca881826e205b5ccd1e9718a14b2dd63576d520e02141e30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb911baf7d3c503436472d240adfa7a5306111310895cba7dd0a03f09c5878b2f9a0d41829ea922d94f9231da4ddda080e993e476c53d4197ed1cbba0402f517d76fa590fa7569665090ea8ba0845a6200de5dba52;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a1d1a986f6d39009fbe428a6d5b70009f47d8d15178c1ecea3d8e0f7fea3b761752b18c01df37e21d1c49334dde1a185eb45f66df28d79d0aabe0b3a658b5a1becc04b93b2ea4811573a8db12a4590d35b7f7af4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1253ab7a23dceb6b8a2c6424cc5e590007110d7f625beeadd32c106a3a45fde4bd6572d8c9097284127352a817aafb894e71d25d518316f7b5549901e5ba86b953a869e31e7dd6a29f8bdfcb3cf4884b485fba7fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6802f44e386ee72a83df1e4559b047ef56cbe0a1036e31624e5cde9f18ce6c0faf93607cf98706c459bbdb9394a0dc8a5ace9edde1ef95d389f52736dba9b773647240e4d34039266d42421d315da0299e1b2ea6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa147bc5f44fb8c50051372ada8671bf70ea179700d5d31573787f47b47a6f620895cdf7887e335e1be1cc0c0a5fccce6b1f2a41de539bc47a384dbcdd49d72eb59eac7108cca5ecad173b091901d900e37ddf8ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83eb59e1ad2cce34482f8dbe174f47fafd70466e1ded1ffff5974f1dd8a9dfe63f4d1b5df61005be0b2cb63d12525bc3ac07745a0160c6171c81694a56b147a4ee2185950b5680be68e347eb05f51a40a72b840de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h735f99cd980cc111937e7418a49ebe5b599a5a3640ee619bfa22094b272614a562f05e6079c8d6dcad1929f2f1198f82cffa8b21dc7cc4d2fa86add1ea0f1e398d064f10daeecc537b7f8bd616bc6cca4af38d0e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa2bb7906f128b4a239a7e04de2020db53eb09febc290c83205a2a8c2ab00fed1b52062d335eb5f541469550458897625a2613ccdd0cfb2b8a422f27e754ac69cf0f3e8890f4ad185da8f5047b5996f2a8d35481;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0b6a87c32ee703e7de779f3ea963966f200f8cc77846fdd339ecd44ac99f56e93b91f63e400e6124ec750de50bbafd5513fab2ec7816483ca3ca0f165e82c5c9cbd1eed34753da994e241d03d54ec494fc99faf7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a583e514dd5289d33bfc545e269b4549f1e611b9b3220535e75cc7dfc6b54906371f45397499c4b10275bc00dc311aacdcf756eede763f38b18278bfa563141bed10b125fe68ac2602e49138d097cff42265315c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff12649bd33016cb349714054408d91af4331de3232ce622619090afc1281a89836e9ed9019d99a47c00adbc77d028c211bc1e5531e3e46c542fe1cd1dadc3acf3904e486ef3c34d32ba6d6c1c3f33f19341636a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b1653b3d3f9abdeabdef521ac09b1108ea1268b9a961bb9ca3a1b6aa3f6461491588cf35b545d3b4b09c52a8d8cdb7ce96a267ba4e3bb4ea4ae7d153f00897e7e06c0169fe2088a83b8b60e46ea700b040a1b737;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb3fc04e127141bf0f886826c9508144ee0e95a33b9d7ce847577d244299439340f8b0cf94fdb9f71f6b4badbf78cde9bb7b074a1dbd0030034206066027ebec357245d0eb59180b9982db83d99f0b88baa3d221c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h210db61d5886bedccd0ef59bbb1a6387390d0d8f80dc8ab77848b7c2b0b3070a2295cd08b1b563f2a79413ac1ed4644245e063be7e673b7d133c9668ee4c30f3dc766964b890e977e36e530193aa7c84ac134e456;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a62d0dc55fd98a83a4739fcca951eda29ee7a53230bfeac8cda752a540d5676b688c77f2e2268367deb479a8bb01024ae769cae29209df6301fd52a573de259779018d803fd899ba6239670bf8c6b739509b9332;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e007ce8aa62c3aa2473eef45ad8af129bb4e6591cc003d3222182951bc6b7e670d46bc7f2034af34fd1184c03aae7079af84d04b97158bd7f56c5147f43ba04d9ea5aa4b0881c746d0626938939fa136195fd1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d1cabbeee7b31bd88fb411906967f7ff6d7f6bfb221d421d350d3b846f052739642412de44961e9e676881733001d647fd521fbcff5b6fb50822e8e1324b9ca80a940176a930597ef1d2ec7e254f9418fd949a99;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f3109c0245e73d37b32bed951af97d6bacc3fd660639e7215db546a7be3bee39e86b21b5eb872a2f67e124ec72b04ac512a0d99def20b6e962a1c104d845259fe88224a45e3a196475171fa01128b471ee4b1af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde284d518df45dd635bcdc560128f6fc39d20b02ed96d0b11d85f13d143e6ade86a327a77c89953250d32160f801fc7448088f740b96dbc1a47f9a80eadc03e9864e69946baaa91f2e7a66ae39af9606837395334;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h174652707c5061c616d3585044e783c73834a8c23d30bc5e4f0ae68e28e06728c962524253ef949e98b75e72051583deec22f85a565b6fb6aba44eff435ceb6d9d873768b1c2e10fa2c060e43248de4f4873a1e9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had01cfe552f02dbf6ca8e96e046099c2c45ac956dfea15fbf7920e31a8905f26f1531dd0020083fe354997e4781ab88d4bc3694e57905ce7b4aee409d3e16e0919cab7272ae8b9c0db9bff4755ce9ef0cf912adf3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf906116b5b64714b0076b3f35b2fcd7e71ec50cee15421ec50d794efcf148c278e1c02a08fcfc3c31a4c78ebb2d8a52dd2a325ff896298dfe06b6966eadd28e521a5e206ebad96bb200243b9c3cf64c32bd4074e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd645f0bb32cbc5b6ea9744bfddcf681015d591043ebda16727040b40458c00e36dbf2ab8deb5eaf8c3a5e8bd7f6c7eb9e0c35aed8f9786830334a5661681347fcb9f07ed2dab82b8df4095058ab7e4d0fc2a135c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75989d9566f23e1f45f3c0c2b7b75a8be703783a5e85bab7ad13b1b1428e9abc3d18ba953218a60b294f24284c40d01240f5f4eabf33120d4ddea39f686d3606d83166fe12e4056f2bf2970a536cfe17802f993be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42700bad43a408944608145a99a2c8b6966a1fcb28eb752b40927a10b6e8f8991ba9299e53e8c2732b25b71b87ee4495035305b219a135e4e0927bf77ac16e1d9151fb20bc4aa0e22bad554c3e0d4c82714ed4b36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1dda8e948e7d9c51ad7d13371f44487284772a65884dd7c2e1ef913382c1cc4c0588d48330fb3e61963095ae109b20471737f7d4e2a9feb78b9840a7657f4f81044e4181389a2f0ecd0244ff34c6a5735c06aa93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cfeb7f8fbd97bf8a171fa83a142c303a1d4b458eb7cfdc9720defaa3d75a1e61cbae9e25d213c976f736d44412589334b486e60afdfdaa10d2d79a68414359a50746b754dc237c232aec196ef488ade8672f936f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b19200afe6b14f028be7ad1cfae4da785b205d1cad46c598fd88ec7d2205d00a4bbd84da8912c1e8b7a2a991d93dfef3540c0a107c949d4e58c68eebaea9309b9876d4df9be0cfaafe0c034766e88d795f40a813;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2409541ceb031e749923061b7f0055cf310e630d1bbe860b24dc2abce51f2ac3df9c57e18480f65074255be15b9860818d447bcd0a4c373737a5f5fc0b210ba4aee3b88023733643f4b91eca18e702a051707e706;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h581abeb3fadca4eb042cc7a537e71e9cf36363b29ef0fb7ad42d87ab8c16b01cd4b58bedc04417aaac0daa688e06a5d3443d3c76a74a7ab30a0fd27ac64700ebf2851909aa8689271f918a868756874a28e0cff08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee816bdf7dcc6c2e3ddb3e77f3e4187f202229b1e988f936c26fedfd4866a35352addfe48067b46069bf9c9659b9c98370c7468d5ff848c3e05c94acad56e31c636ad6e9680ed4bed2c825efaa6a025e001d5156d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h533eb4248902bcf30aa2c354f1da572cb8222bdf5e9421923c0e60f474c26c606a143e27cfca8934ad800983b5312a1f4decb4414d41e287418d8a172d31a34582881e07f47569b706750c159eca73747f377eac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75ae732773a71726a9b3ec7200165c42e458b9a8e9bb93c387166c3900c545bb0fdb249be6e60d8d640882e69705ab07246f66e46330d84ee81dffdc33be0801089f083014a325c06048feae9a89491405b10712a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65590c56425648d3ca6651193db946dabfe60a369ec5ac97c5a594412bcccd57aff53cfb41d90634680e40a45ccae99c1d26bacf98048f882038faa42e3e8f19e02af40376b90a0bb371a2382d6cd4b63689ce57c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb99d5d5037504c3e4b30ef8dee1576eac49c9af327635515202a19397f779131fb2c8ade9345feb8175052a2fc78e835d3ec9b72ae27aa13d5a69559b252f3acdebb8c4a5b0fa3cdd918beedf1a39e6baf875929;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbb3dba9367aa217cebfc8ca5e298499fcf73bcd9a792110022cf8465b3d2398bb4bbc9bdade4e9b0c85a955482c40349dd00b86471d2bac7ffb28c5e3e80f734adcad6095a6bf470e4272cfc28d04cafc5308bca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc2a17867d0d9db240c7eda43028dae5c94481e363d9a77d13f4746e6f6e7cec4e5f2ea65512abaa23475710398a226816b03361c84b42cd3020d4a2920cc44723b709a19043e232f1dad14ceebfd017c1b12a9d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34da0de0452ea8d41e57fc88cb6217edda0b12e6e33b9c6544d24ac079282c2257989d97c4844e70cfd2aeebc9736167009788728353833c3f2b587380f60f34b41a17f523d643502224ba2bb3a1bafe63cbd825a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fef8157841fc690841ade4cbd98b0378dfde4dcbe2da486880a245ab25578d75f21c945e58fcfc236ff89ffdffb409c100b61a5499dd7208e91e37bdaafe89230823ff2f10e0169d959cfd4875a2b89f2cddbd41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5eba4dada34c1ab808276a3b196db28d65119b66c8ce0705709bbbd2dfd2b4253f7166ecf41c72c30030fca34e069e8322273c667bff42cb164d48283c2d52834d8f90aae384d8a2e19c8e82188f46d356bd90ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cea1e9483821ea1b6d1ee9273d40e38f48227005a45794b49373f4c4233022c1ec5f57909560634c6114870c5c966a82352d0b2f2288f0d68fb5f96134115e9793897f0631f3c24f7ba0cb71cecc8abd81061bca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43fe099d33e785d76c99ef4d92b612c1389ad764cc0643155de9cc9749710f4e4f8e7a04460cfe882fea3926a84e64a87336bde8af42174648793461591528e690b6b91420813049d0e5ea16b4547743f98dee122;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c48e129d6bf99d465d19615a95af6854632ac0725d416919bff515a01f1e42e056592dbeb1f4bdb4fba9db1bdd1230a3858437f22fbd84da8601df2e7c8192c3cd3b0296c96cfa02f2eff6d138f5695bc2e1a8cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b380601e23deecdc420fafc6d3be8973404dcce28af4a5329aa419e870feb2eefc7ec7b0bf78f75999d264e4b91a95e495b71cc7e139fd0834b66458e417e44c1819def9ec09caf1041a1d9714ed22ccba9e6738;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c6e8a8b73b13e182a0cfe5da7d8fb44ba351212fb41913a9f7f4d3805272ceb1a949806d5af1cee88015976aeb26ac263a33b76c4f85791642e67fa50da29ea9dd669558492633e39aef34b97a4a1df60b4e241a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b3d948ae035938aac704c1b7418ca1e54aba1c183277c08bb396054aa13276b6d654b0dd0a8f2954fb02146767e53ddd1f5c40a6ad5c6fa91fb3dac99eb9ce1da7d8342961fa6523ae05aa6d24344f67bb012e57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb015b23d0d640219c08f9529ac1c380f9d3fbe363c8f4a2a7dc11fe016b44b0b3cf881aebf7d9873717b3f57be73f549de3de87e3904fc0ee812822ff6d7b6fd75ae0d3181ed87fe8b610dd514eba37ec2cf0f84b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda76765cddb56c01729ad65e5e740019fa773a71449a021c9d9fadc8fe7c0bed5fbd1428a5dddeb7fb203a7842019366d08cbfe0378aa43d1ff9b36105bc9b7ca05b8d9a22347623e67e887274c75dbcf2e26814b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h712cadd1ceeff35990f0d7f297588899a1c44d14f268bebd32f8344768f2caaaeb258a89594852aea90fc1c398da4e842696ecf684755248966abd4f99b9a044a8f31fc010bab7a161de69531f573c50e504bd57d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1342718c84f707808190beaf863d23c60e5664aa48d778f5fa751d62eedfbc3951691a08b01faa38b40a2e1c95b3b61263f0cc523277c7027a69c0b00f8845c4f1bddbb1892ba95b51f9cd1e014792a02941bfbfe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a0ea04c2dfed14bc0288349b53cdfe66d6db450c9f1aaac555749aece479a9f8bfc26f8381c913f9d489b4db1905afb05d91d9be8f6098b5f4f45c6863d78b0b4bc2ffc9e176c5042dfffc3f1ef39f4028f9a1e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f1603ede9f2b6ad5ed2b9a68a6cb2135d48e1a07c1df34682231fb50f44e313a5b0a92b2f9fdff779c35b29f4c8e6a748acb13082ad0c4e13c50e1a95f44e05872241a3d8abf99c753ceaa1cda342ec248eee7b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0b1b2742df0c13e16623cfef2617656cf4864e7d5fbfb088df8b6f800a172f479e60fbe160b61ce20c7c114d86ba8a32d997b78eae65230fdeb3188cce2464e6e26fc2a66f13627124c294d3d72371726b7eb9f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h374d654b104f67da6c4a8680322289252b4d23557289c5ca37a3588cb5afb31f060a6f44153765ab45596f8313a21def28c0f92605075475313254b07dd03411b040aca5ef071debb30a192ebb82037a11ed5a9ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d72031501a460006e26cd16e69ee98f4648c8e8ddd1d26acbd21b28c2a06af8054712f3d1508b4c9012bf3f849538797b843e84881aec47a300a1f1f685dce786d0934916d5f0a6d7a63658b28ac15e445be714c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d3558f44fdf6a8d9fefc35b09e5bb3e24cf770fd29dc5fc0eb2765af2f0bdfbdeb13b8572a1123da69fc1a405943ca306f293937d15389a5ddbe6b34fb9bcfe78dabd8a34a881cb67f635ae014e62eaf86bd78c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d4cadf3982c6d2e2603f420da56e748dec9e6d7ace5c303b3c3adb56a2c2024f2f7d35514f8961db95ec9b26ed87d6c6ddec7ffbecc190441c33323b21081b795458adb4b919fe9e93656d3054a2b21aeb6cac40;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h783513b7d42f0c86738619ded1b35e80ffa1f0b2d6896ab964961ef758ecf33828c4ccc9f39e90ed6ef7b713d58c515c8c8833e64dbf06a8e3486d09cbfe84ea95f374ba6f1b606d9088c5c48798e67dda77ba92e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf49f6a42c50e2d5c63739ba8d8b7ab8b4177b8713e48c2cb089570ce91dc13a301ec7ba03b30196dc948d6a98d689f7a98713b596274d71f408fe83310b08022ce11fe3b9d23ebe7cf7b575ec51fc89b24bd0cf9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea47549c112dba8c48faf1e8fdc51d3b26015b32509c15a4855681b794c189a8b2599ab2817adf0394900cd4c366fffdefcda1ee03f69b12e09ab09add0e8648d6133a75ad55ccc84bdac0f34d14d31b926c31c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he19829f0fda5babaa146c6b44f81b1b7160e5bbc5f4f86c4b202161660f337a282345291040f84f9a783cbdb7a8a5d6c30fe155198943e92c692ee4593532c5b8e8552c8fce0b5c36bd5b57283e5d468c7618abba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dad5e4ac222306a32d48f271e4e6282ddd5c72e214c9192ca764e60b359dc87c80c0dd79119d904a6e2dce97ca5c03d357a59499f7bbc91481b132280583eda003673c684ed1c40a25460ab4c74aa447b685fcb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f5a551838e34a6fe3be4590994a713e5bfe0bd130e47d7a27346b68f03616b3aa7b13b87d0679435e3797657b4e0f67d21df712c508788b2305b0c8a5ad29907fc32d7aa952c1355c9daf92bac31fd607bad56a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91f97537670ea4500269649b1d936225cb9ad91a29b0ad3de569d3f34174a0c7b88a674f3e16c8515f6b21fb9426a2cb08cb8a97772d120a3e97b0ca473d7a201983001716eb5f414cf7e87f099251362d5c858fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fde6e68c0461d2b42fee6814144c6a18e22bec3c509fdd053f4ae24046d9882be113101d0fb25f254a007177d78de26827c746b249531c4380825d0c6090c157c3971d5954a1fad1cdc822c0821e28c1e954d9dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21ba92c90b62bad22e33b9464332d00c46af46ecb7c22dcc6404c3d4aaadd7e278ca3da66a59d8d0242a474a2c2ec0c8eea07086b52df85ea55ad7598200235e85409eb9d4ce60552ef50c874ed4d20f60c26a24f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a022aa0b91d0b40550fa6ecbe689ba7befbbbccf3ccc584d92b125224c29af0a200d49f886f19d0071b120736c608fa9abb5578ad9dd12a87e0866cf4bcc6cb51c9cca7cc3377ddb0ddc4648492dbd63cb9c81b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40415ca0782dcea59221662ed9e909b4c64d9dbfedac03114878aa32374a980d4da7635278d45366d943b319a55517897ef1c7a4d681fc772cea07be1634d2d9768a7065673b17cbd339cba64aceb0e75d6699995;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he516efa7b451b2785d6a890e1a0744a18f69c4ee561b2b050d53d8a59287485604d907e67e14d094e1249fa7f611ea0684a87ace49448850542555a396f9dd044935cb510814ab8212274b1fec76a9f95fe04b91b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h189815d7f158977e47ea8c6a28babee3fb2101d8ee649168feb307ab012322630de1e08790f3f20284b0e9f96c97d72d60d5bdf059c0e371bed27fb3f784a5e6fdf0bc6bcf95cac36fd5b522e31f0192a8f935894;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83f5353fbe8f9a8fea5cacd02e1f2e350e06b6e752844e9f2d5982c814ff6511ceb45b72dcbe06dffa5f936301dd80862aff82f4285431ad21b8ccbe35acd318895e45d1572143ff06a7f559d3b91046d187b88d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49a35ae0611131839374eed9a0424ef6d6cd137c441cdd24c1c7e0b62385ca445a22f6dcba98352ef25d8361e97f62a4e57360316219151fc91098b85d6268bf1c8501b369ed38b6468e829fa1ca1f5faeb80b602;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he665a203059ccd6461480b94afa7c97baeb805fd6fc493cf34ab1fd608de39de698fd5712dafebc3515d5557ee8989b50b9cb5a628b4072a77f85a6636c7b8301c4890130680d71d3be36e96dc0cea83ba008a751;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83234e092cbd36c062280ddcfa68077259efeba396a21b8470bb2d9a3ef637195937801655dbecfa8378d233600d1978f84cce882ad492fd8c016ec8e19f36f17ffaadbd6eb4303693405fd919b9e3ba114717ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha169daddf300a665afdc8d1c86d3f8d5a261e9f3ad4c9b6707c78ab3e248f2ad1137d2270ff6ca0ed1762fe6c8738d0ef3f9dd40737e90004492ce8d05ad051383afe5c361befc47aae436c02c74e12430f35dc56;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h631bee2c8648c96f269a45bbb424767f322282572faae8346c3e91427287ea1902ca5e34036224abaed8043adb4bfdfe72e4f015aace38b70df31bf89adbb61064c03e2188b462c7febe4cc1e62778569703066eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaef7528d215c87bb57242fa14f54055831feedd7a8e46fc166d79d1c8dcaa00f280294f697714da1ffccddf980ea3baf75c3f2c5e152b93435002cf1ea58c85ca770f30200cb548bea06245ff22928b90f1b1bf2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e30fb749bda9e878fbe23c5134cee5db29641fbe4059320315be2de43829d91dfac8d3064e0a5e65412654ce44699d51f4e89efe4db8bcb5e58f214f57f957fce6c9f93ceb3a561ee7ab8e67114e90afc02a1d55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31a9f017c0c5516356e4cb3e18d7eb92ae1419ebbe2cccfbf289b1391c587d17cb3e2e7233d9d0d88b8bbbcfbfbe919c309e2e5385d66fe478157b228767845a27273fa27d7410efc3ddc889140bd4d67a76caa4a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aba5cc51b1bb157e4211f12e4290b7c96f5b1887f0714c2f0192a1a2c6cfcc6674bc4197c372c0b452a0c8cd03b4630970d3e2a102dd60aad410d867246e1faa7345cf5e64d60e0bdc55b9b89d5a2ac044df8cc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79d7beb312d710e145d27051990fe541fa1c5f1ecfdefe4d7affec11903ee1ac0c0e67c8bf23ccbd229530498f479a69155cd27eb6d25afbdb785b35af1d6157e2790a14b6898558c19b3c5804268e72fa0a18d9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha689f92720b3d0304f789706c0b732ae27dadf69ce86fca85276d69ba9811d27cbdc826b57eb59d0aa455f064bc79f633108cc361c798d022c9b99bd35bc04cdf3658f63f146664f1c807d0cf0bda51977202021b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2f61fa50ae651c59402eafc102792497481e90c384631e033e98a4d9ff985282c7042acf46da04c31b0909d6a2b08636eecedddd1b58e2bd448d84eba080490283411e03ef33035032b73afc09ee242fdf88c063;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9414ba3e6846c59c7ab507ddffa6a356b2b4ead04ee26bc2b852173beef1a6f02b72db2a0b95fb884ab3b18a5cd39ac01afca699efed7d57ed012945d0be38f65a8bb322b00cc6c2423cae64c36832ffca10e5bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc35da8bb5e0c7a15ac9cae311150efe7c90dc7403f8295eaa3fc21259c779930ca3575bd8a4c35d90d3a636d5f1e9b56df5e2093559a7f2495858c233a322c25bdea054440e2bb258be4eeb8645bdb24344734252;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h645083c11124bced3600907c36f87a3305c5c54f4e8611770c77713292a02cde2feb56368a7629001caa9897bc0b800d7dad00f885897ee8ed7624f0182c59b3b111e6be341b77c24d135ff811f0eacf6c985cf22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf56122b84a430a6c7fc7cbacb0c1674688c70da1a433cbcab8533829b8ae1c72f205157687cb17a9dccac2e8bbf9872d78b6c3c450eea1a1457b55e5e52d53fb9f42c29214e6b894e24fdb240f55b03731c440e2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7530db095c0801c01b1998992046873840244b3d92bfe540aaac3bc443c70bb614abf33f992fde971c99eedaa314a6b77c810f761d24dc3f4bae9ba9b8873278193aafcce1bc8e2c61bff0d9f2c6a2931fd09ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7fc313296a85bba90efe0b9d0b8631d90679e5b8aa266c159d62b17b6481b08eb7e1d3b23035c9626c8d2be5fb11d83f063ca7f148f0cb0bd229e311fb6a6b9f3039e04ec4822223d93488ae5eb523b17f2114bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadc7eb315a689bfc91b868d5a86735ec46452ebb5a22be00e82349f0e1e203909bd37f3a8b91b40ddc4e9aee1d1df51a9b4adbaf0d0986c8c2cbbea5db2d5b44e68b52c31b558ce6c7b965fc6b7dfc1d60aa57787;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5cff47321f996bad97d57b55c28371da56524705f03dfe5595dc507e8b7030deda203e04fe8a2c2398fad68c9da1612458a8a79155790b7070f0fd7b0ade2af8a0fe64ae8734ffbfb0e9ec9fb430bbe004fcfd58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c89c9ac4860fa59dd9412ccd73888ff0bac4bf6242cdeae1b898a60ef38c9b66a67910f0424b74054de7670ba6caecb09c7f2024a915ab361df660b45fbddb6d959c5237cd40775bde7aac5aaed035c006a1ada6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d85dacf598171ad62f127d7f990fe1ecf6c2713e442eb0b656bbdfb889075aa03f6ba78f2df894dfaedbae2d5b8b15be0baed40f9c280a00f8f2f377cd65acf793351a251ebe4ac1b33d3fb972d1007e1334a23d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15f5af78bf37c8bb5f6dd1f365a92c57fdc040ab1a2b8cbd2a6b894a61befa66d7534a6d7c168ed187e1dab0b4c611e7d3316bbe2d24d4a5a4dea3229aad4ad357bdd92ed80050bd501a35abb312499570862827;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3bc87b41243a621b125fa8033fad751bca794e546b4d82f25c9457ffd6191470ab58176e1a26309d36d40d4fdc2f4e7a3a1f25d67209e8ea88970b111f6b1bfdc3e60ff9c739a46d4fe8733e06fcf3cea6c30508;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc6189b1c9e059c6217438450b0e4c356fea3a33c7233bb76fc4d72bad6c98485a386d5bb4bc72229c9998ab1c3b1734130a3e5a1b1ac7cd04b3df76de59b4df461ab65be0f815826d967964e842dcb7e0e7595e5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d253e98d3bb9af9b7b3e6441d6911315b1494a3c4dd82e763cccf6f4cd75d5d7d3db33d04a73aacf3c4a1560699131446db0d8ac6c0fc9f8bca1b39789355629ddfd74af37ec3cb3da37fd7e4cc9e60a0c475688;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h783bfeed0beadb9d0a9d4d1f42aed900d8572ae6f24522c87f099c4ada99ee108ba1b47a7d81badb338e478f434aa83394b019785723fb2d31ad9bb383cf3f1c8c3754a30d559a638a3e73084c6c6abcd6f728868;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he76f11e5f052eeca77f65677ff95776aecae35f76000ddad328677189e08c0e220d63f09d052a768de0120082d29b0d6f9b001032630c599f8b7cce89ceb0dd82dd1f601b88fc0c50704483440079f5c7f4fd6fae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1de92499439776239d9112bf4fb9b5f61d5a27a697cbd3f4b025d767332191dc9a5ecdf1b310d3ebae8564a7bd69a6aab6e3460cd3fef160cd83fc865200f9c290d83cf6eddf1ba57bd4f24795ab9c5cfea3969a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd8aed64bf5e78399fe8173844bf48c995a0d4c94649c039050e14893fa60faf427bf785bad0ba315015e490bfc21f743436d1006827332a00a47a16b7eeec723e812d2e96f48c2162350a5d31c58babd183afebf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94a7e3c190531b0abd6d23c5191ba5ebd03befafea66187bb4154441934dcf3eb9c237d3c3193eb361a0feccdb96d716c083100e6d80d88d94737bd3b3b27f08dfc09b0f152fd6bc0441aa1618aa1cff12c7716a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6237b9dd38139f5c91e143248362ba7f7a654d6582e5aff5661c5fdcf9d559c0fbf578f8e4e843ac85f5fa60f3355093567a811b419de3d9b52de10b43fdf955175aa17cceb2319d07a4304eb01931f5cce95f47;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f1af05582a235b043e3df03ebf99a6a741e7107f23a49505b928a96ec5692e3186b1ea0867d606a7ad1dc802f7b6434bcffccbc1c14713c0acf76947398864dc4ff42dbb05d49d008b2390c2d8b32a588c66af6a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a6bf44691606c8b5fb86c6213d1fda3f985c37c1bfd187b9e445420486d7bd96c616bdd0a3d847dc074114764f08484fd90c4c18a84494d611e89e7b399e924c490c2be2cd1780b691026a601aa3be154407fcc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e93ba2c3eafcf30ba222bc373b179fbdb43d0071972bf381cac8f67a3e4d990550b5c26f96f19f1dbf460f612429a78350455fd7871498eb0842d683b25845b0a861121d1bd618c813696683db0f949500feef25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37143c000ddd1e7accee3a9bcad71aa1c91b842f9fa0aa540f92d52d8345450360ed2ec7daa7680b4819b254c0ecab6e5691f853f70ef03d4a22389af6c1a89325a3ab515bcb0e0000425a314860ed8831eb2b872;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80a728d39acbe4538c465d1db5231ad86792595d0b8f8abef86cc1c25e93355968259adcca0a900addaeee3ba70c1786c0324863c8a6e85175f84efbe5b42dc2272da1600b11bd7575e656a20d99f2385887f6524;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf71c4bd25ab5cb0f578b054fdb94f13bca56fca08abe755453ca41bc2db11ef892b680491fda1f00ef72283ef176f86a6e54602e4d94a1da9000d17d845e705d5a70be3de5a8495a80ad426fd8c3d7d35716125f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd91ce0d0bd8bc451ec28ff3e54a5d1bd30de9b061d7502e42b4e6b763a7a9fcf3bf28f8619a76d4d6e5bc56ffe244837ace9a4361a786c6532e9b1a0e5511a4f3254764ca50799100422d5bfa8ce5cca7dfef5273;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h268ac6b77b5761a312683fee50bd86c7bf0ffa5ba0181de5d5c6388ae43254d9fc20a922f6a28909389d7337bd22b4ef3db53e9e910c97559a848d52559e50a7253d989bad0b76c2df8993060b292d638898bf01b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57619f397032169e35e4e20b4f9acc397b82d3a0676b34b70133ae0513e2ba65c1314e599ce0bb0b708c476027920f8a67cbeb9a91d2efb40368cef8e01f7f26dfea1bbb569ac8b6e283ba3d4c8216b38d936924;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha59bb72f9b598a905eced0f0ec3f05b61b1b3a255e43910c25548501c2818621a7fe926cc7fe52defe72045e5ba710efc885b9c7671a95c123d5c8a560afb1c9b9a4bc909014f6aa5224d997fb11f6ab99608a7ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0f60161dd99f2d0ae870c320b3d895284681f3d70897eb2d72926f4904f2acb829f41ad9898de2a759e8d501772c8091eb334406a2ee96f4d80fe4e9fabde33146d680c7dd401f07312342cfac3a1825afdbf3d2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c8b49bd5c74dc3a8e04a806004aec17c842ba5ada4e8f8d738d0ce9a4dedcbb0dd6101e86beaaed096a7d0277ffeb3684ea7723e64f00dbb85cc63f1c63258e7c6e3ba19b5269f897e263cb620f39c34d1be339a;
        #1
        $finish();
    end
endmodule
