module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [24:0] src26;
    reg [23:0] src27;
    reg [22:0] src28;
    reg [21:0] src29;
    reg [20:0] src30;
    reg [19:0] src31;
    reg [18:0] src32;
    reg [17:0] src33;
    reg [16:0] src34;
    reg [15:0] src35;
    reg [14:0] src36;
    reg [13:0] src37;
    reg [12:0] src38;
    reg [11:0] src39;
    reg [10:0] src40;
    reg [9:0] src41;
    reg [8:0] src42;
    reg [7:0] src43;
    reg [6:0] src44;
    reg [5:0] src45;
    reg [4:0] src46;
    reg [3:0] src47;
    reg [2:0] src48;
    reg [1:0] src49;
    reg [0:0] src50;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [51:0] srcsum;
    wire [51:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3])<<47) + ((src48[0] + src48[1] + src48[2])<<48) + ((src49[0] + src49[1])<<49) + ((src50[0])<<50);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1318d85ebaf017ac3f9ec689a957702525ecb78c246afaa55a186c23ddfbaf5ee4a4a45c19188219eac1c95f9546d57d74fe61a8bba1ece74bf00060b11ca5bceef408bb36534ac9cda455f2458f274011eecde7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6becb0bb3f6cfe7cc017654dc3e3cdeda382d8b692c1b597b5ea889d758c1a8758ceb765410c09591099870b3e87db17d22359e5ac603f7ac272de611c90191c9248fa7d168c8efc12e665c6c466db336f21fc31;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h543f5ef9920e3a04a8f6a7c1c84632f44d5f9c62aba15850fae3cea8b745b0b223be382e439bca5463a1a7137843a10b1edb4c87629aeedeb056002a751bffb36fdaf1ead6b4ab235570544d94a6044a64a7eb4b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h862045721d47c74c26cb76235e70593a140cb8a284211702bafd714ca4a2c990a04aa14a5146bcab66da7c12b4e6ac3dfefa93c0c71b26ad0d0ccb20b3441e49fd26f42789dcef5d8853465e96e34e775a3cdc60c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h593febd2566562d81799e3b30db1b6f874cf1edddfaff2567e504566d75d5431da349cf6a981b2f7289b32a8e2bb572594ff9b0dc511fffde95fe0cb25af101b267dbe45019b7920f29ed8079b524732b6f0cea26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h486cc504b0622c9558f267c50ad3f7d4233a26fe42b0d78bd3ed3bf1c343991dfe8279bc8d08282a2d0cdd0e020c7ee01ffe0470da0ba03fe17f1262f651eeecd39ad98331a6df9532524bf14d0f51d85b445f090;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9872af67e833dcbb456416c61b1e7ede8717601859008c45f4f95dc9ef58b014e0cc126597d32f17c43a78d053de835375ef2da4e39a4121bf835aa6ca0f9adf9a72434a48b357f2b17a98a2730ec9b48b0e52ddb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ca921e2de3d742b62b46a17c30d1c418504d1f21f5b7903e91269840e2f0c9497f6d162b7e8576331d1851a98aaafe5571bd37aa27f796d028b7616e11e09e2c9c0bf971695c9f7413b5c0f507bd866d9306c36f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3af6135e8e3a70a3f155adeaf54bef54a217f98441adb1b7fb79acb9dd2b37730d4ec5995d60d908f579d6e03196238c1916b85f21c9446cd55baa3660fbcafc4219bea8c854b7ac25a28d9de0ae384849d1fdfc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha832ebac88bde67c86635710341119108e9aa256f519326850d0b50dbd0606daa2018e9f071eaaae9b78621c1c7f7cdfa76975a4c90840d1d9c51a744ce0b43d17c60ecf4ca03a7c0730dd4eebe42f7bf80cbae44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec56dfa6424172b240993af857ad5e7f2810bb573afa8d2356ce53d77fcd4e87a04030ee6ac92722ebbf8f1c94e760ec81f892fc91f0528306602a939c01b6258891db488749da3bb11f7414b2eca4de191dd0a73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf81d0f5d6598bb518d9652c0f6b144196912e84208091a3ff9307f0933da9204acb0a66b858279cf0221a35d92024db4ffaab83d956519c2ea79946da3fad9dae2d8beb401e192282f8183c3f6843dbc41d728e53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0007674b4485a74d910b289153706afaef5b900750adc566dc332f12d1149a61da926448efd7711a21a7a2435faa795049fc0e08a0b8d621ff86b16edc9491539044ab3ce41133fae19391831a13993f12405b08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddf9da712b4847bb8f7e3fedd5e4923827eb553346a88695e3d24fcdd79cae45d5335190e7bdba074aacaa13902a83d286649824ea02bf28706866e1e307ec97d1357d999e3517af35a2ea642c74e99def4a4381d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha78055d595467ee833f1c60eb217c97119ec098269f796deefe2c20ff9fc4b07e6a389fa98ddc7e897bc5b68077a068a042253d49cb754ac0535916e01900dc8ced86944bf7f23238d658b8ff5705672a56d9072d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h965edc07259bf9a660d05cea3e702e9f6ed1bcd49dc8aa717990758544629f0626a59f9945143c0e79e0740a678b70fce1fe16c483eef4b82d370bbed33a3c9733497d7256f9edf743fb678f1162adc0897012de8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6aefe41adf1a05f9f6f5aa7091e396f7c325ad9a450722d9d330ca61f32fe3d21383705eef5d07fa741b801d4b90ab20c2dc6cb66614f7d7dd88e5a51271947a29e14c0d3da2565506983ff0ce935cb1cbe6aec3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef17889896f0cca54037d57a571d9b1b4ad5eba28d13a240ccadc7b8974d63413de23bcdbb5cecda91f456776042a3fb92d505ca6ceddaa80c65c98e3ec905ffe213a877be5d8e8690df559d8cfab36878f86693b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ce59ab82a5a2e2cec53ab744bd39aee03bd14ce8dba0c7c369d7f70acac5182b1b0b8bc9db3294f41f22f07dfe8cf81b141c262b49e5bac4d087389a1a55b81ed8fc19f9a8063965718691689666b94f310b2bac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b7253019cf896fb2f601dd056ea6ba4d8a1edd5be6fc20ca2b0adb76aa5597ff8950f834579cc7fbb6e6838633900533cdbc727db0913b4a996876d459662edfc9b25b55bee887ce3f1b8875624c5fc828cfa54d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50647f4dfd6aeb8c8b3dd3cfde96f8230e1e02fab0e86b94741c8ab1751856bbe94ae2e45c1ad320b25f211f6b21e27697c9d9abf1c94ac9156a14f8a823bb1230ca4e8d683d66338dee64fad4bda60d4894c1c5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbc182333b974d9f09deea2ca61a4a9d80abc10f02c7f11a1a7277c958d452f58be172650e614d356c9028f68c213494ca18d3d686e1d46c3afa147bfa58ab9a9e69f4b40e70ab656348ce3ac715a0c65bccff524;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba63c4c2c68f213318b0400b583eb5ef5b4223cf3b78815086e919bd738d5e65ba4c80028f81dbec2d81baf8a91ff12a8d1b05d6b8b20e546110ab5f0bdb9f8572e458b2877069bbca164521ad19a82ed71abbce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ed7904f6a386e56d4c03dd38e28644c56f48422d5fb7b992599fc0a222933a4d8e87d7a44ad14aa2080a9ff01f56c22f5c2702cac9bbea155aa6248ffcedd2cd9962d0223f8668b9bbc11c779fa6e01c9136238f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae9fa7855bbe06ee5ecfdb465265fcd6f5ccfd72d8da491fa7e5f924ce1c8af9b64a537f00e0ca4336373244eade79f940f7be4fc7e0935ca23363773896c457bbe45cbc336fc02738fbe4e084a23cb43b4e0cbd0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3337d6a47014bcbf4e1e61f65edfd2b50d91622a64762bda913aff6c7416d4df8f8ac543cf17cffa2dd032416e60709d587ffcc1a8d6c2c5b4796788b923529ef60542581a3ccb02898eff0d67aceaf71b0171f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he14276ddbbf2b6540731a3db8bb9ce4e33e39edfdd284112a89d1904f61aa84bda34064a35f3940389cb57cc34a60c171e70dae8aa82157c09288d9fbb9cfd01c98e403d1dc12a0788b35cf15129bf193160c3512;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4967e1ee0b3a9efa633c3a9194d6eb8b0e190d0d903c53a92f4f2fbc7699b9db250ae93650e3edacf0d7d238acd9bf341e5b87bd20c63af1c8c57059eb739838f7d22be2fe264c8b585cdb318c8b9725bcfa550e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c849238b6c1fc576aba7abdead45cc415947627707ef2a035c7dce241327d7a2adcc3dc29ae787a68ab0f1e182925d3540f95ae234d087fc7c721d6608c9bc2954bdf1e741cbefea3460a9c9be4f71700519243;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb638e400247be410dd58d74236b8d7c69482467c70a8d98e67d8921eb0d9de46030032ddc6e2b8526e2298aa3d9af7b9d76b0892dc5ff2975a90bf239bd7d4eab9a5e9e65a3973893e80d1a149bf25a61d01eaf89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5ccfaa23cb7a5e21b1094c298194379c06883dfbe4450965bdd005d5035b1df943c804d535b9153006f56c78dead9566426354eeaa2fc85d22aa34a0163998f0d241321e6f189167d241e0b3629915d75e269b1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58f0bc5389267af643f8c1fed3050b36d4af21c87cbf46959f8a68865615270d025e57b6b89b6465b5842f43799dadbd9872222ecb64cfd599288cab7a2392d19aea002af5e412215c11bc07c591d4db29d925c21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf093db85b30ec9c8ea400f341486dcce838c385169a74e5656c797706f802efc1f2c68ee1697c8877361610bc7ecc9bb62b2958e8dc3bbd6d3a6f5ec887694fd3ee0e0bf245563ea913736f635878df3554d6d30f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9673dabf8b91c0dcb2b1a013691358317bfca6473c02272f94ca684f279c572cff2dd6eee21932ef1b51f6883f43cf55125820676686e3c5f41f6f79783e0a27b1765783042f8738a4eac06092676492caed8a952;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf97e90fbfabd1765f4638624d64900181aa139b7b18f1edaa0270aac67c39c981c10ee530b0f83453b4a5328086038b9440daa318873390a10b4c01705bd1e7ce47ccdf1860a60fcf2e8281235057988baaa3580e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59378fe78af70310cbdc3763f4349ac0050edfd0615e225eeb6032df8d193e1fa2fbd2b77c0114f5900cc6d662550c235df4e92bd402e05b92f6bf2291a5ae0ccf89fbaa09105ce447888d6d72e54ae4b38bbab0d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h965d9ceba8242e54a9f5a110c40821025697f5af9d91571c57e2b6f63494670161b7f6fbd669a801bba2b508ccefe62dc7235ee0177740ad8d36f17ccb61e4c57f9f5ce3607652ffe30aeca02c66fce1ae9283678;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3424b7c96b0f8783a6cc32664b2d77429dd3c6c0055b887da0ba6ea4bd5e84874d14d7c8e849a69fa11da3d140076fe80b41f63eda82b27d7dcffb9645d4873f51469f7126edb2018a4221f1f714e83a0d1246a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf53a87107e85d82ac4fc4a600af381235bb70316a2a417b27fd9d94356d87129761a45b6c31e3e864ebc009d8709c0de95ed05603dba086d70bc692ee524bb668cd08b24092f8916f3b6cb6a46303a6edd3a795e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc027aea8a61a01eab1d45ade6020593967fdba0ef2ebf49cef38839eb59d99db906452947f1a3fa84cfb84c467d0a5ad483bc08b37035978ad246ea955958ba57212bc746bb76ad1b8d8fd66b6a02eba0b840f973;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc135327eb18dfb53b2485b7b365fb4eebe6338478aba8334ae53c487d2b091213f64de9301bf27ed711233605f33ebb53483da370946e5d77cc4addd1f8d5dacb207b394278b1d92b22321112302f94d00c072a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he48be97feba7ce911bab2a15b7d403f0d819c964a67f57276322e22ad600de739c58455d388f0835eab60b0fde6490b5daa810b1d1d628f169e15ff9c59b5128b8a58c80c43a42078602e822c69944b35fd3946d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c9f3b8b8c91ace11e4e2a997d404978a93a754bfb05887c4848cb88c43b802a8e5ea634fd34b0fb9db3c281bfb12618a773f707eff500ab37dd484799288644f3b5cffd06766b08b77a399efe834df905a5f7c80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34fa96739fe53bb34cc6412f955b4b33478ccbb110dbf6e62bb57169440dfaf7c8f5dae319f7fb889757e006d92802a55b2e56c2fc101e787a179547837a36d505ba50f15271c3ec505d0cc866b537aab136559d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacc1fd01aa1f45135457413a09c1146f5c7c05b14d6037f92a383e576b4497f6725c7333b885ed0a6ca9ba24d52dbb7f71fe674512ed6b0fcc7d4c9f00f275759f491232bc61305d0c84f8f18a01c6875b13b5cca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf035396e610fd91dae6546cc29fc80422b6de73b35d3ea928e809e28d6e76c84d8ee9eccb83279e8546ec531d20ad9c369d27a182535319efd9e9a1bf0e48e20bbbdb4a8fc4e5168219c65a43edbd13eed72f96d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd72e34820dd3d910b53426c495a31e080d4ab16cda83f205b12f22444a53d95a4253153f0c43dd33dcfff73343ccaa6db285ea79deb22d2cadca0940ff53af1c59f52688bfddfa79ef641ba1297350c83b7ebc8f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7cf5e7fc02169980efbbe0ba8adb2ebf8d2b7947d62c9d64e3ef792323850fb5ae8b0a1b41e09eca105b0a7ecbbf2620bd5ffc4c797831d3be8502edc286366a53c9c6abc0468c53986c84cf9d98e9198dd65d2f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf824f0b4a80ab0a3e3590cee88de1c3a4cca0cb9f6e89b94a8339bc1c15d54a16a13d4beaaa279c7557eb9bf32c313a4239b5582c9d3b4cd5a2e4087d0444ef2444b683e040351e008bf370ae19922a953e827424;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41b2c1d61e36306ea6cc0235347b9d42d781674245d799d4147c4e220d13f4097e933ad5ccee62c05a44f28f708aaf76ae6103543f46e2cd213cdc00239a88cae19607d82c2e54246510a1e55693651671bc51e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65eea8956c1aab389b29360e6772ae349b4ad1d784d2c0a84ec79c0978efbc99b268527e1b589200d2d77089e2c9a074ef97d656b402e9dfc2d19d030ef27d47baeef4f63eda906dc03200bb10f7b8e4ee0f0adc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4b36c68730c741ed4af3abb4832906e1dcb400dc9e86358d81812d937e3e3372364b7546886aa453aac87a038ce1494e4c1f62caccc33028b5ea50b3d9625a9314b42c11f56e42877392979937310918f39ec20f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde690e9f025b9692f90236770731e64e1a328871e4587b28d993d6bdf163447184b64fb23aad6c60b2dc21ffe7c4e38cbfe8e0fc74fa870113db35dab8ff6d02e82e7ba4219ffe16330acabd9e107745c1ed00dbd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he52aaa391141514b0c2f828659ad4fd7eb48bc1f031907ba4bbe6c28d11d7709cb8797230f78a24870249028a21b30d69029dae53d96624edb0d6552d4e09677d7fa80b396d46b6b20a3d46eeeece39b3b02b5de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h288eb1674038b6c27c31630f0787f4dce2fb7d2788849976b85ce7fb892ce39ef248569ad20869ab8deea5c423c2dca49dc768c839ba3a5e1401f4556f07fb4d4aaa6a00d695e199810337107f2e70831666cfd4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb00b057a89fb20b876e4d7eebed803fe123bfa8aca5953221124070a1bd88d88db43516cb4d6f111d92388a5a7e6bac3e52359c78877a777c4567ed83d46b5d84d0873acba0d8258e0bab34a5e65064e6e7be4a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec4ede38c24fc40f94ec76df2c6cfee8509880abf50ab31b6111db503f5ebf887cf832ea1cf9bc16a26359e563be1b273f91d6be6d006e39568b0d893555162621f675ce3a399f9ff103b586bf3a3e889c41897f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6cc5d14743bb75260832761d01a3e9af5f1fa25275fce65c86f4783c3c399a7805035df3170ce57297292335217d3d78555df7d611ec2d312f1d8f4bd8cbc353c3ad36dc87dc0c21f56b4af400b29a765963f054;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he39c4690131ef06cd55de1dc5949b0cc716dd0f86d6610bcdd57a0c745bf0f43e1895c7fbfc4b444817905d2a5502af7b0283b9d749c41827094ba94fb9f2d7365de290f86b485528c2ae213341bef87e05e84a07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bd96634dd79c589711e4899c3c87c3c056c96da795654791c152806803442d4f40cee232315cc1005baf1d3285d819ec2505cc631b42f2471805afc200cabd20038e0cc59292f5f65e730907aa3beb9c420df4b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe89af83f24724607b1deaa52eebf6a4ae206c8aaff3ba75b742958072f63d0c054de4e4dcd6934cd2df8523faefc666f9b4f5930a1712b28f5fbb1cb92afa78f9d649037e364e3e105501e32de6c94c61e9bcceb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcaa0e4a95f348ad2b6f122a9e1a5ca5ec10e807c787fa8b242fa66e2560e3a26d389f018c096ec3916fc00924f43ecf423edccf40a83c210e690d233927751da264df72b041ad1cdf98b314d716bf0a11ddab154;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h982e4875cb1f6a51c3f4a813de09cd8e6cb1b1496957d9b48be7ec2732dd330fd7e12a8f3bda890bb08b74b99a36eeaea3be767390fd5ae46350a9e07683046f74d4398b43bd048bb70ee390b1734c523b2a44c56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31736ab5637449e70b6f496478dd33ec958af0e694969b43079ccb2bf956211cdd34ab0cda88731f77fd42f64a1bf52a93daf17c50e0e73aee00c892f7fcbc78c1c1687005b7fcd49740904d4633a5590e763ff3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b982d87fbaf1e830f7d5998cb939dc459984843552fffeb64c31bcc4ed6c9db95f4d964a89f94366ca9008c2d8551de0b348e92d5e9dcb3efc7603662b923f1bedf178fa91a1a0f3bee8cad2441139de011fadf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2dca14c6c369b881a0e70ae6ff98b82d43abdae6e323b380065fabe0ae1b82c49db3cf22296b102af657a6c31fd66369d4a20329cfc3396857de323a5e99ce8c4b3bcbc427709a83c83847697abecba32384290d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf4795fd4e7a859ecdb99396fd13d6d2fd77d6f61a5b0785c8a7466b8129223aa1dd91282c2e8ee09e71df74499bcaf7bf3d6f549c5ff0f0276b59e7cd208e4266682763dd9ee8e00cb3749197f6d9ba8dfefeb22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebd4c2a3c22c30fe992ec50485637bd9d29dbef1dd9f1a039ce0b20339fb4c5fceee49e3884a61a9090e360a7d4261291e55ef829a0dea40ec0f6a6d961c61676cfdb9b64e49edf664d76b209aa8aa76c35de923c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fb04f56f549ed5789249ae08f29f1b43037a8f8e8b3f78f12ed4f853bfb05121f7314150130fa4c1154a84bb05db0eaca2788c60f95d93eecddfe45ce1dd935ce177f06b077cf376bc6e3df6258d9bb692b2efbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a38a47d9f7b6fdfd6c484dc8d8989a0240d1d8d380d4d59d98f0229c0118bacb883e2ed49fd6cba2bba67011bd47398bd0f1c3260518804f240526a5e2127f511c1a402a0bdc0d9e2d652a468b2983f57bf47e54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4effed806eda49898342be96f3d24f98a7ec581111098811a2c021bcacaca5b58ed51e1241c151b5ec38bb854c2455b08779d84ffc58339b62670e725be8bc30a102a59bf96550d1c4d23abe0f6cf9d02ec6e49b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf80c1e43fa127d2bee86a6907ca3e1f3cc7f137b01d4e4caf478b13e89683a27b19343c01653d2b61b703814399b8cb40495029232f66b415ec1903a4f750b714f148e961ba0be9426afd13020771c03be6a5d0ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf365819e4c1538ef25acf83d725f8abdc0bbe274df05363b9571bb9d1aba63ec707eebdd7e32bdd1fe1e6a7e7a38e116840c56663d2121569ec15cc3a03cdb1b81002e2390afbda01879589e41d217363120096d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1bca8d44690a668d4432d15b1fe057c9e59387149764f4bf2fbbdaf4de68873811c116cf416736170fe89beffc011a89e7750eca36990f77a1a153e5d90a7ce0d3c47a02ada8389db30e67595782e09d2d0c62b68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc84a83d1da1138443dfc6ce650cccea42efd464bf17f989a46ee58f73da0b0e4d677b3d18843186cc75d3aef6bad2c35be5ca47d5088abe2bbc91d73ca0ebfdf05329a9487aceb5f9dde082a5633eac39c064ba92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d27b06c3f956a33177d3618355d5775254011a529066b276787c4403e4551573c686ba09ce90a9686e983b2091ae1e2c56f689b19bd9cb9424008fe45a351fe816ede8ebef622fc789f3619d797873171118d215;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he14e7562329b6c4f8528c8b8788cc6b621e3f0c6e10bfec1797fcb36baec4d0f15b195bf856a7f1c92dcc771c39b68e36f4204bbd77e1df6d67c49ecc43accf4fa3d18409dce7635fce048eab265ed4bf1c0eb2ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94799579cc8e0270a9a6ede7a80fd11fc8fedf58d7b38d012489d220bee7a660b199eaf59adba2b271b51a22846aa73215f10b6be60ce1b95df88373cadfcb6ad8c96bea13ab7e5f4e4d7f1bd6b9210383335e40f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46514bc7d3775f3d1d7777fc86f1b68dc9425978347232868ed46632ae1b4beeb51d860851cbceae53430d409ed7cacde94f1c8a21752c96d30f666b499715701a43f9f772a5baf0c572fa1d89fd7a8fdc94cf96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c6449ef2e9a44949ec057265255dc2dcb4b1a1579e53335011eaf96173a611bc5fd9324282d0d2580827eb99c4ce750c46d74c26a89446913a48414ef227f19c1b924945475b96fbc44afb3cea699928b86ff224;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fbc1ae3df4a6584a92732ae54ad4c39b11ccb4cc007d835396ebe6feb9d788cd6263b340ce9e04a16d652d03c7609f70736a5f98eb84629ef99c077cc4cd7d095bfa2552e8b8af51fdd82069184d87cc6fddd806;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha856252423f60120ccb66ac0a7d6ce7536a74dd1cff17f82eb98a739a631242459bb77415b81b55047e4494457c09ebc896ee8d56cc48c3d968b91bff010b16870d033acbe0c1ed9824aae6b372bf80d1fc16b371;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b60616de7ca96318f3e96f0f5b8a1bc168fb21e46b1629833a654510f18b4e782eb10939737b522d4b1b66a5b0ac5c290c6dac45d2cd41396191cd13198df04fef3cf7559f7f7f13c3544f0cde72d576510aee50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h347e32549b2441d32cb7c6631f670ff6622371e335d38e1e47325a388f13ebcc86ec279edac369798cb25ff917fb61b5cd3c2c58745df5cf7eab77c0f728a759ba8f0e69229fbf87d77fba6b26d206187bdd33e81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he34a762b3f4d8cf91e496ef226d7bb24b26e86299ba7dcb84d0935f963d040661e716447ccb4aba17185cc337bc4e55319a220db644fef2150dbc416048527498c822a3f8f9cda660b47dc87259fcae08776a1271;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc984e405af958828f95aed12a68659c9e77177e5c64058fb876761bb4c171156c8132831e9598d7a750ad75c51acc7a51cd47b2259d42b059b76b344ebec87cb85c7d478e85c363c76bba449011aaf3bacfea3d01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcc541795c652727b37a16f1df7662a4790feffb9aa0737a59784f788ca6b5e4bcb8f52bd1dc55dbfa0f0d6d500822611e969a4b9c7a42d555a930219fcd71b39ada168fdfd1ade30628c1411ff91781c6d598dac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70c2e64dab57b7f71b080f9571ac929c665c452a2188413f7447cde5267e7e7c88435c3a25ca88c65c99bcb050e3ad6ef526bf8d1f5fcd904e9a789fa5878654791a138de89a6519adaf4414e8faf06bb20bd4c46;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc87e5eafe0eefb158b06c0f8e5dcfce6da1b7cc5334bfb46c3b95c0949593fd6213e29b66c2a62fc32204a57c513a94f0978ac17d91e652d26cc00086fefe0c4c812ae4793ed3e7767632fe17ede6d90e0409357e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42a0e2986b6a580e842697e7b040836390972b1305440ea526e1163e63a49854f4113fa7f6bbf5da69504d6e1765921b36c70bd4092d81045f539dd2069ad8183371f2e176ea14e243e4cd443429e79cae88926fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb3c5c27a25a51a611e7a5a3d8802edc8886fb55895839da13898e2480466be980b5ddb2e1b51e89f6df18dc4ac993b0a299aa5a2eaab7174f76ede57df51249834ae9434ce0b9660f960ac45bb55954cdf1efe40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c20186d28986075487094ae573738d8baa636165c5adfc9e313eb4e53df20d3fdf2eeae2c12a551f1bd9e55fc07c16610895c2a291792d648b9b10894909fda120901ad4843ba002add4b03e213045b1b10efa41;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfe951c0951d716be8f568228b5ff874b84878e7a5de3499ae1465dda17e89c8ef5c1a290673270c1c83367ab62dd4af9a1f37c43d71a063cdb8e77005c4d6bf51a9f56b27622ffd9d2f0d3a965a6101540d7f534;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf441e7c54cb6e5cb24aa1759c7ff1d025d120c15b73cbe177acb79ba7c571d6a4580f1f3b9904e87c545d78523e2d758377ce424ddaf71ccd37c90ff0d34aecccebbd0e380176b5d126852276bf094ff24569d05b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6eb4b3caa3dd5adef47e8a2fd6631054c4fe1d9359c9786587c174692e5df5e4cc05cd96c9755302f4cc6e2165aa0879e458032c62c86c13bd11996be8f9d9b4ac0dec6d6d0bc37424806c020c121607fcffeaf31;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30e77acf97d62a146dff0d34900bedbefecc6b9778d5874f5c43c47056c3cdfcecdf9b2aa6ce90ff2d306256263c6b0b85998d96f6e34ed12b0f4c6341909034d1af23b15d2c35fcfde17e45cc5f824510cbfae51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he36410fdae2fc940944a8123493db5a37ac1c390b6a82d549b28a59e88e79ec15d155fcdd5ec332c2e4abd2c9111530556616bc6036b58638e17b4c1d97d3490d0b49e04489cde50f5d61e513c828d841183e3f89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h662cb7ae639d35da54b589f9ac72023e9c13c8b5c87beb404dbd0d1d7aad7f9ccd0ad3348e9af0d4a478475281bb28a269a25e8f61edc1850d07995455e98a3b6403d0e5d924bfa512a3234abc6f2ee27179f59ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf255211e71b45a0d24407e5ee4122dd35ba36a0de6e1b9f991b049d8f74928e3df89497d8d3c8567db1c81deecd0754c037546ba8eab52d7e6188b626f3bc59f0d72cb524d834c2a086eed46feec2f855b0ff7787;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h131c39ed513bc9e2669ee1a56fa9b773fc34eb125006a1cd6ae0333bed9134b2458e6d6939d0a0e16dea1ac2b416510bab560fe85adccd5cf2fddd0e37f6750f34a91c7e3a3a7fe2819284db8811c52c0fa24a55d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5e5796ada095af0e57ebb365f16a71329d9224246995caecdea7c50b727895237b5fefb8945c4380ae56a0a229abed5e7c4e877c9daa2cf78763ad1d7132ccb40f75877f67e99f3422548fb0c64d7267b3a7d57b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dd18244422b34a569c0a527ab5b0a043f41824b76624ae531797607adeafe9695c47b5ed1181a82797af161de53cb4a35497082496dc5077c5ed4f4dc2a78e2601443e8612572ccea2bd7d2c163caab57f08ec00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h676d75ce2cca50f161cf296ef50226fadaabe616726a417fbc484174cb9d161c50cff8d3e2cbe3236fcfbf474b81d3431ec2acf67509e4b770215e5b930f382399073af66841dd7914d0707410444f66afb2c54eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ac09229e3e49fdc02454760de91de3e43b87ce890cb1bf6699b10e90515f9a7cf58153598d13ad1098b7a56e231fc6498cc3a5b899165d13779102eb10ffade5dbcbe17074e98177171677fa92a2ee4d9cc3783a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdad94dc794a51d141b2d13f8498e0d910247c7cba028e87b5556a514a2c26ead745f1fd1153673d10088b3dafdb9c6ec234fbcfccce5e7d01ec831a6edbac711290e7992e0d99f8003aaf8e1fcfcbebd929593a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ff861ae90c2ace50639aa34b2988b3174f1dcfc6d390ea02a6c9dd67a9e8e254fbae7936490726fa1a95f7a9a00daacc67c6813f25b3d37441e2ca8dfceff61c2725abb82570e4729f39016812ca515fd443563;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec9ba9e5308983371147a16a77e69bdc205d8f41b5a4a25f3de9bc3978757c7fe6a14e9d338bdfe51909afacc98186b05fc03987bd5bb2aff74649b9813b38a12df64a1756635540dd566f3974730a2ba94f2559d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3517844762aa7539e8ecfc567e13f93f7a0f863df839473e76029cdd0735755c47b499079be4a3fda1cfbf652a9f77297be40548c88bdcfef91ee618075b7801cc04077098221ce80a0427731b137a4061eb4978;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d4bd3806e827330331bba1e64e30a08fbd72ce7450f7b750e7921333cdef79fe4895c5a2526104892a62ef21e3d99b249a004c528bef5ba48d9faf278e6f129f8013edf440a03d5825aca8f97da42c157041a4d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b133bddfcd6bce33f75012e5bf1061491f615e2e13b64902cfab13dd06dcfcabcb1420783a2e79d450dc00aea73a7b1e43b0a504ffe89e24cad80f7dd579767f242050b82fcd9c50d12ce408b514eda20d2b75ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51ba4bb7f189825356ea3c8e6d8718bfad70c5b443c77abb3e5855f472ce725c524ed87e08ab678d9813e7bb952f574a8fd5c32f08fb32c59d8753d2d5abb7a164786ec337745a7dab6896815c6a1dc405d4e8a14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he23d26211dc628d0b0bf399f6343bbf497239b4b23a4a1ecd985f6d9f91c2bad2cb707d5ecbbf435023e3e19e194f1413057529887bc45db7bfda07e7dcb1d260b2f8a60ca7569956fbaae41e1d429827ae979fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe4b97e46f90ffe7c0e71127b8742ee8ebbda1e8026d6fbe33df566b68cc753e4df3aa10ca9b250374669d05a29f676f6d6ec71bc60e671d1512dc44e18fdaa9b1c42c586b2a0dca6a25f9131d235b2099225256e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b5a00846c9bbcab8df76745a5880d7fbabfc7013dd516945045f444b103c10f7ffcaa28912caa5e731cd4401fbd09e291904b2621c660f69777db27593e8b8a348e9f7c4888acd19d977e523f47d98da8e28b095;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd84fc268090ae597c49a23402874ad6c9a2fefa376ff56a53c2cbb8dfd5f64463f34af6126401dbbe45bc620a0ee0436509efd5e93dd294f53f7c5958621c48c03c07f11081d2f340ee072c9cf8f21a46046b0302;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd699fae6f5b9e5f4f22512a793c87cae1e3ff6fe40ab9cb379be3ad3c0ec086dfb40373e16856c30fdf6b7d9ee6ec6f23a5e966658d27ae9012030039a7162b44e05523f4e2ad8be329b90f20ccf77caa9267300;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h574ac16707196dbaca30af13c0038e3a6270b87f6a6950787ddece8b48dd27ea016c022ba35504be1d1e16f26bf7ccc8a1fd2e1bdb9638d5368d45ae072b2342ab58e0822317dd833a11d040370d4011b2da26c52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfaf983924208b4df820bcb7b574993db463f3c5189c3a0df3e875e079285c0d85748d819efb67a48c05c10544fecb6319e1467558e52e88cb6ca020e2cac058f046c0195b57e7973e402fa682dfc392b00d4c568;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ad631c3ca79a53adf02ffb85d0a4dfcb7d0221733aeb1224177c90ba266785f2ef57ccdd202376a56a5648e046b752399819eec52529cd76eeb63a9ad7362ca8cf2cc56d2f012a0b59af1a550146c2892808ffd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ca74b15fd0c8ff3073763125495f3d844a1c6cf01f32227846d5a34e3ebe480861a1132df424898bfad2708480d383dcdb967d43e6c18a1ceb819e310e1c39380c4c469d233812393297e0a06415b593eb1d0eed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7aba7c9138051b89d3e88fd642390c8ac8cab4e9fdae10f8eceda95a87ce4296d5c71c514ed2ebdff34cc15da3dbab837b283688acf7e5055fdfc4e840edcb5138468cc0cf993128d36188a99f78fc45523b6c10d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24929c32b071ec898fca703fe11fae0416822b8a5785df336eba571e17e164b117d28cb653887842a6de828fd557876b0ac5d8dec3246a25a19a6b2edb5b0e3060cb1a216a23078a018702ecb6c3234438fd52d78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5bce295f533ff52f639dbcfd86d35602f4aadea17f76253969becfb6b36f952e7daaeb31ebc75829a646bb7d167094132c013d6f2c8a2b263e0df6243bfcb00226b6cc73dfd8c5ab2a7c5f6ef090ef6835f2a92d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5378910907ad7672863bd51928018f3abf09c87c91f934c7c69ac2b86220776f88a644abc6c94725f1901617ed202844726a06b22571fd07a445a249545d0c9099c9c0a05173e536c936f1f568def36c2361c1344;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h292e7589016060ada216127fcae0fbef62375631471c1a06bb868b8d9ea8fd05740a0e3477d721a0aa90166efb9fe4fd2b1cef956d1be577ef9c30b26621893c789f63d9f205340b5aaf028fc414efcc485316df8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27718f0bd6875862b233a669cd47f9610b9608fbed4d6ef37ef89f9830abcedfd87e4df4480f33742500e57512e14fcb7a015db1d98c3b84746217eb5222907412a48922d8f5fa0be6c7bc782845c5b52878dae29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1089173364f5cead73a30c4dab0009fe70236167fa4140957c930642d7f093480ee69d7f3066a592ed12c36e046a5e7df216e1178a40d136f7d4b73c3f9aba7113376b2adb0e1bbb3f74c07bede6eded802970f83;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h620067cc6cfb094523942f2a476bc6c8a19c2ef17c95a926ea06eb5687ea94fb7b90bf43a6f3a52a83e229bfe091ea1689f6c07c16d6cd98920bab5bec5bdcb660a9dd087e8df94688dc6d72d7a995541496b4940;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d43642df2720c9d377775166dffee8daf8005d7a33013e72adc1cde3bd0de76cf16f9b7b65642c6d390ba5323b1a3b2865ab7fa6d90d7464c55c1c00ee011cbac9ce0b1a7bc758b13d5370b918ce1e67f1233342;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9901c84f23133af9b45bd1410338bc050d0a9be70faa64c9d75009bf49d0d8debf93fafe5643a17f9b14c6c25877c1ee5a7862a26885a8d1176e4974e7f98ab84a8f0a282fa8b8a22171704ee5683002e161c0581;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6ce5087526f892d33ef981996847a555b8ece170af32e795c45a22743149907166764cf5e28532c3ef3326f13db58386cbcebbfcce7a2064b28858eeac6c6ebdc4a6b3965bd055b532fdbeb3ec8bd0be00e10a93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96c3a143815d82d6a938f696dac49c8869d3f3f13269ab8d232dd78bb764ce83fe35dedb0697937136f7a386b48b4f905a27aa4a65316ce1e189d7a2d5fb6380b650a155dd2e5e5a8530ebbc2ab7567746536fae4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5290983f1acf1f7d383050f6ececb8bf4fca6114abd205098607796c96b93403d6a419ce8378351914a9443329f55706ce0e738fd55ea9f3d0eae2e83970d8b51096dd51427d48d702f7826218ad4b1098fdf6e56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4be9eed4ae5f8580039130bf6d72cc616ff8a7ee982819e1d694e54bc757f74af51b2f588a5102533e6777f469afd82d342c9e51be0da8c55f6fa0f5c01b085b5e777204b64ce58d496d9015bb4b8c097c9960a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4528d4fc8303eabbaaedd279331786ef24311690a431955aa2b48ab9aad2667fdb263f67d017ceeb016c4af59e34d7d7a4ea024936dcc680e6cfa87b8650f007200ad58dd002d78cc788111234205f6b903a3a130;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9a821c499f1dc1b9af43da1f299af83e6df8ac0db0108899661072b693a1516a441d2b040975e565718dc31b0ec7b8df17150c6077d18ed7996e911aca1cf550847ef78065703587bd5704dd1a79013e8d8b8617;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a8cd2141ca463ab36838f84b090fa4dd2f3696c1c35f94d3e9b148958b4e386da21186354250cedc359f9ef6771494ecb7ebdc484e2deeaef49cf9f0c6d4859ce9bdd796d139ac40270fb7b9d6047923e162ad8f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83127fd5e925bd4ba88e9f4714cf8e5994615fee4255455e6b74fcebe035c671ad225357e6bce09766803b890ac6d70bc39376332dfeea5d0645ed7ffb9d0e5840d4f48160385aecffef1c0e55819b35058400495;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb790b02f152db1b91818dc2d9b9d45faefacffb7b19af9ab05ee870c33d47d559bb63cc0f5d32d1431996a444949fa5a1855535065a11d10b445ef461e75b23d092bfc7db0e98c2aebccb5a0a1c9127ce0a6594d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f77a1a6dca13da84618b94945059c01fba6f15015361c7381ca83ef43aaf9439ace601b5f19bb3755ed366cdd3c63ea8e4414e218108eebb515d498560b89a3126ee1bce613ddbebf004709be2f364d58ed3181b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43f8bd7a6a2bd4c88b7ae8edbab7a1f18aaa2b91999ea18032a59b2d6c01326e617e80c6efdbcf6ef76ee8583e5da0d4c052f2ed75c8be9707d19efd67f8663c0391135310427255c36951a4fff2030b163d3d3b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb156ef2e2ca2042e6a595a2e6358c26f96c0ceaffc1ae9b871921e7592a5bef47afd9728460ad1f4b7425dd27f4966827fef0e4bcf2b08bd5f4487fe6913395d7a7999e248dc75191b3950c3108ee93f67a5cd57d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75320d28fdc824e267f0181fbe95da0c4d186f1d524ecf8b917acb0f979ad400d233c76e82f762d5528347f8642f85f7fc92a4ba2042f5354476850d5603f1530253b1452d673de5c484710cfe7e8413b674a651e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h984ad83f82d9e5e208280816730a5edfffe6f3ea4a8296398ff0ba20581db2a14dc15ea7e7b10f669ff0ee4bda2c3058b9faaf91f8bf75172e3258f26b6f93535f59a6c0782239e8d44bc00f368a92635ea8165c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8f5b619fbabf716c8bb484118c58a7b8cb8ee0041dcfb7261b28b302adc2edee45dc45e13765e41e401bc89ebf37190fff37dc2c331517bad90517a1d07eda5c4de30e03fe90d0324dc9fb5aeb1a07490240a500;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb98251adcf05c33866227a5d202c56e5e031be10f751464f2ab520699330ad9ff114fa0c966b2bccb2e02527bd3c7e1964e5f81618ca0e39d09cd7b1b959980f4ea9f7b0434189b005d71ed2b31fd30d4fc68e6f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc774dac36a2eb9313b278e966c4487d7098a0576de3f410df1611f9937fb35d953fbcaca5b75fa26d46f491f0546ef115109e9e68d0f1a940186f43d8a86537ab160d24da3dff3411cc0aacb4bd5629f0f0f7fdd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h878089cc700a34257daa25c14d55d545c3b784b07a2f5345cba8f2831226246778452b475c5d01aa5a77a123185499eb60bba22b85a260f070ab2b4b7c9e363c823bb0da35e6a7073e08e7fc6462869b84659e3cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4476aba2ad1ad441d006459b58577d95eda485587ae13c635dd12f2c9307b3aba1f6d78b00c6461f0c01bc30824b11d06ce8045b001a9b6c47a2ec4de68bdd06b634923cca41a44f8af464b12801aee8bbf9c729c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3bc54ed6e8fd570e0afd50dc51b5e8e891d3cdb4a0cf0560757ff99307fd9e83de6f5a8519135b7503463af24ce947d3a80cdf96c3f0cb8971958d44a5e63ad0320354a55ef03957062c7d3fdcfdca44c27e01d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb06eabef12ce1a3c7162b2fbb21dbcf51156283c694d0a9188a9c7cf632a491715148f3cb58f7a16071b4ed8c339b7af1a7d642aad71c61c6a54e1f2bd143831275ecc68bb1c9665427a925888ad15fd4a1184bb0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93afb8176038403ee75ac6c5bc06d6c1ee5033313b85d18ccb408750094b45b4c15ffb81527dbf648d7e9e592b909dd1c07b4f6ac5f99b6b33eae6a076f8d7885ef3737a00d9037adcc424a9f881bb18fa9fcd894;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8052e875928e9b058e1ca1ade7eedce761da4191490a5e7ae2de2395850c45c33b5eddfc8e2091e96af4498afc8a9d2a7ddd6d658a5981eb722af145a7d99cbc407ed97dc06be6d4b45bf15ca9e6d70268be61987;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6dc661d0afae7ae6ec7d71bdf967b22d6fd1f594a335879c59bf5ed5fb0096655ca27bb8ee0357a0d7757974c15334622904644ebb22eb79540127bfadaae7999946ca5aa1d83f81a3b3ada291fe9053b731838b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4d4ee09655eaaa5e881d0094af6c900012eca53f8bf06ba41dc259f934985291ce412d4174b782df0a4f234b10cd398e5eb88cdb400310cfea03a90a38007fc61f8d0f511ea6b36b6901af3af94cae47bb899b9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fe33943638b48707d32b20aa6622f6b9c0f6d1cc856b96e659f49fb52331ade00816db2854c35323dc596d9020e43043b06c0c300396bedf1811f5d9203584b5cd563958f0108c3abf4e8142be1bd67bb032651e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cb9a3f66eb4d7780fa8d1aad3b8a371db092b57b9bfefc3efb626d389ea75e7f9ed8d8dd363c7fcadad3830d782217a41e7258fad30f0e14cbc1e7ab3692506438998431aeef9d1aadb8abae72e9f27965de8f68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h952785f40df7477483eef9ecbad629d0d003891425993819184167783a508f9c3d0a19afc3f18c4c9060639c44dc98cd34f475ac43489c8628ac3c466f0d2f884490fc1eb984420bd3e72e0a0cd942aa6367450cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbfd8fd72680fe23d1b8068fdf48ae80648f1b30b3994e38236ca8ad9fa213d796283d3193fec24df242d9cfa085498a9acdccbacc2c4e040ab59ea39f35ba32295647916cd20349e290a16e84077c507fe5ef7c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cba50d408eaf01a094c989ebd0f935bfc862dc125ceee9c13feecf36dd861211d5f7b0f0ee418524ba7c3947e0bf95a82a8f0bd0d144db93ac04c8ec215a188808a83702ff8744816abfcf467d077d8ae0c9c7b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h226a65d02439f0a8a17c6fe3815b56bd76238e7d0d4e5d2363949c98cdef3bc207c865ce7fcdcc6dd72880ecf5285c257cc56d9ab68c1398cc764157941c1be9b37618a41d8fccbf5df1337f60fc4c2e8c9964738;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f2bd858b71c5db61cbcdf6492bc986b11aaf03a2d83b8e80147da5e0d8e73b4540ca71c742282f4fa0b57bef54b9c122537d6ef4c883e0c2fa2febfd37da94b664a6fe33f7834deac9a476eafd6cdc037db40ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b4bb36633c1143bbc3f3a703d1a4d3a56d670218051e4fb4ceaaf51b1f5d97d291df4772b181fbed9a85fc93f64f465ebe7005ce9799615cb746203b4e27ab8c62df75ed4bca776f0a15419b89663f8b9446d308;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fdc220ecbad849fe768f0df9e7be0e871d28e14f60348c58155d359c10b035b4818c6ed5b4c7dca82638de7dc2b6bebc1d758326ecb75d950db755e15f05c33c5b351c1278384d6a9b9b5430a85b93504f50ff9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7563f8e0c389f6887f3ebfee2b1fcec2efe9137272b53587ca7937e936619511e8262d313dad6179325d74fa0dc9d633370f87289838f4c379b6c4e7086bde42a1898ed929042319120fd83ed4106988440a5a1c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e64b8ff366695cbc15e94635faed8df2bb3f171eec5226367a5cd31f21f067da7295139e3df3f4f0e329cd510c381e1b7774c7d471ba6b979ca8d71914f0a227ff50b1ed6bedc2cda45f9698dbaad859d736d8d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h791c37f2e5dfaaeb6454b2be051a5cd43db0b3db632761e58e1372d94f5d9438b42c89a613bede21ddd950390aae47f349d08ce6c71334a42c5c32b1e6bfd408d364e24d7ad424c034353d1f6606d43c8b6124694;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45b572a1b5280cc4ebc5965851713f34537cc089b8a35f8c91529b7513b2a56660537338caad905f6bee86dd848f794321ed05eeeb576debc1f53099fc0da0a4940ffd6cf6afe2778efff53d163eafaacf6940581;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd75c73d038ba4b458ee9cf638291d9ec0ad5594f9387d217de48e835aa9fd6fb4faf576ede0539ca3d492fb81b8e266c7d8916233c8e8e14e380833c5726fc345d20846abc88b6909b2d655428f0b31fe1430d5f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee5e432eae47f5fccdd2c670f9b5da56fb57b562efa1e2c00a72beba41a53a7d0cb2b6093af78b78bfcaf0f299d3c37598c634a3dc11e731e760251f6c4cfffde8a65be847ef5b3986ba0db504e381b20deb6d8fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb444f16947e65f6aac5a01c2acf83fec6df9c81b8d579a3e61a82589c20f3871fcc79ead2c823845feb02b26c0b34907f5ee07ba01a149236fcc592b8040dd53dbe8577a44e440a6a6417db7ca2703653e3e2007;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he57359888c808fdeb0838dd3e314b8aea0055b43c3bd06d2027fa1c78444675c2808510055da492bf75fb5ba903d96e6b018fb8cb676a5973e97703a53a07d0f99bea6f719d075c0297a992aa32361e5fe432bd73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb64b0ee78e70ec23ac3cf20ce6bca8c9a4cb520a6a570f2b56ab9edaa43fab77869e045c4b035263707e44585f7784586fb9c0ae162dce23145a11096dcda44a12363c85f9d7a52d58480667651546263e84c973;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd14716716ff81f75044be075af265d74dbbec202614558d7bd0ec5f53e2109803ab9deffefc1ffd17e58e27b844709f8d78cbd5f5babee795ac408f11d4148c3ec03271a6b5546eee03e532fb8c4a37f91dcd5515;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd12a67754c57b160d36294791b1c9a7e6dc9d5c67de4e38f62d55aee6a7d327411f14fdbd61acdf5eb4cfee674bc6f64981eab78d08485c1c99142596d3a8164538bcfc1224f6068ed9deb7398596e94cb95b9780;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89bd33a0ad59e438c4d5a782c7c464f16e35a6f6fe48ac0f41ec3c51a9a268b6d4650e0bc8f19dc7d8d7ed82fe26a6ba221b88b72b44ca28ef32a0b26e1341879781a65a4c957ad7deb17ea2587d3716c51415e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c4aeea9cf6dc26265cf1e58022baa8128346cfd699970a6388c36696dd8a71003bf3d944d56a8478e99a65c2d2c4a5b7364f5ca678e1f76151285535b6182c6194c7b8b915a3088815002c456f6390af036657ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb07e0bd0c2f96e30f6134513506055d6acefc9bb4e7b67489e6e9e95c3d73632ab398f7ed65442b6385db4f598956aca08a280bcb4214c33a09e71346ec6adeaa81a57e8107061510904c03985ed2b69f148b466a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c606895bb8abb63a210214db8d58c16eee2ddb884d6a1d0ae64366aa90d22e1a61ffcfc649419344aa065d507513fdc2782af6f7dc0e72d596ac1c2fc17f4840ac27c6f8b2825e295344871844b724a665fc6c54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbabf077bac008569795686942cf990e880cd4a59c0b8046b2663554f8e3ab93edcf5c565654d05244c1ac070768fdbb371fc13d8c4be9fe0162e92a9631d1dfd88b26e63ef63f30e3ee82689ab53c5abce69f4fe1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3967e3b7748cc4b903e44a1c3b68e05ec611cc9f8870ae51485c11d67567c76933ea3fcfb5af5ff946e78d026ed93dd66094719144157795cf3ef195641fad13f8c5e30f982ca4e4a552ce4806dfa5fe9b655404;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd06b52c32005aeb57a0e69ee5255e39e15a597d2c89aff8dc9020f0a9c671adca0699be057af1d18da4b9af2874de2cf0ffe06d13bb65becce39fe289891b331ea985ec1bf7404fa4abc9b515c1b87bf42c28eb7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e9d352efb75a140e77626dc5e05d0a45b178a48a16271f61e7d6e63cd619cd509ecfdaaba5d8d184e7d34643b43fe401c0ca1a39adb72bc900da754eea3b2362f2d6ff492eac82a70d22624c8b7eb084575f66a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8945b48faf2006f82c9d3fa1bb3d29d707a5d44bf4d9a30cbd052b3cdfe90b10bae39db13f9df07fd9867e401737a40f1e31d36f03ae2f74dbd6e8b596967089923e9169c8f8ae2826ad878014d7cb48c585f9639;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdccea50444e7c35b35cf4fa30ba24b8cdaef9b307615e8437e86afa4b9d3d75a023f2ca4fbe6ca1da80062d9a0494792fc89a9837dd165eb5002ac1147bd9bdb1966f46847770a4eecb00352977dcbd854aa3f586;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4c69c4089054bd912e38220b2065b76207bebca24c5b9302321ac4844b5c049cb4303386102120b437cfe6d6a3758e6eca7fd0658b65d552301483d44a01fd7cd51d09014f27a45e753abeb41aa555c0eefbb857;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8ee2d93c5029220ebb6b8ca25212ed0ccdcbd17258779842dbdf2758acf16b5030adefdab640747b6676aca5cea72c5b426ea0949db734d1e7944aef6bbe4ecf4bc4a0fe037610079167d75254de04a85eb4fea2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2c65156db7cd96187db3dfc82814b245ccab6557c0d9fddd4d2f42ba77fd60ecbf0d018c853dde8bbd380e677aa1093d249f06660cc1833ab082a183a4e948b606f090f0bf438726305d93812ee6472a08cbe1ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39b2f035c2bc74155033978d2c73077d4c6249f454aa3777adaa44c24a3ebfe84da1ea78e51c9f15aa4778e94dc43c96e1dde9206c098ab335e157c678ce43c992bfd738da9eaf5c53c3605abd6f22f1dba9f345f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed20baa7686ece0c6e04af218a43ba5a79c2388216b661ea19325c1282274065751c473062edad3674b4eca446a510349f475c6ccbac4e3c4984e068e71736a6bad1c53b3682c84c71961b4fefddc93134c41e105;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55f3358c5bc45068579e9accdc6d353b76a9f66d10e3b34a80dc353f09a8747d509a49d6867e27f8a8dae2a728b4470281f5250c31b3a6978e194a7ac443c729eed858a43a0d8f01b472cd5efb4aae191ada923cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b1137bc6b72a23c4b5bb18968db6ad57536de787d61f4c9be4ceff6ad709f0f8cbb146d6a555b5ed26e0334869b4cc2133e213beba9586fe72ec5ed36d47fd6f62be4bde2d7670b87bec0690229b08a3fece35d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e893ec8c12ab27a056442a85c98158d7b28d610c86994a070b9ea6f2c2a45855ac505440cb0034f82564bf87288c13f97e776b5bfd162d3992a2d4e5d6419ec8399d65b35b8345f8de15d01fc7d848455a94e2cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb240b4cd35583589cce53aa23df42900ce11b3841b9ff27e52f5115cac05b30ccb44ca0b3f62be1368db7f04495729841dd763c22638b9f4119e3b92561dbdc0e3c4cfefcea85efbd8f3ed808a30d57d770e7ad3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3320a83b0b3fe3b150decdd525e4c731c478519412c8c5e24be1b5a0145c3219f90bc60f40cd82f7449af39f748adf8276823ff07792b5db0283452f7723ae078dd36d7d0779c24ab239c15e7bee0a1a87dbc0d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50d2772306db8c89dd9b600246437614bdd7da4de6a0d85fb8d3761abe60e3eb480ae46c36af83674c17541473b7973a8dd795062dc5897d52762b1bdb0f952a8bc546d068c738d91107a3001bdcc3adfcbd244d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76f965d3b4524c0c47981d1ca9b1d47675d00eaae1bfc410ce4d78b31c7e46d2a7eecdb73439ce4cc8d9e8549114644d21608bfe57e07b93a2ceb41714fb83b4f9b1b1ec23f191832f6aea1ef65986467cd837cd5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1100e22bcd35e8ee444b3b1248f0371b9c4724b03d6bf63bffef8f4e7902df9fbcc8a6a44832d376b50eee64e688fcd00a9fc1df10ced4a13f3ddca93228674352ae8d8ce052ceab7b5689375dda609d652033665;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h676bfc5f2194442f4f870df41932056893555352231f4202671c880815657473cac87e0a6db5315f827648fc7cf0c5fa0fc89cc0ef09e8e05504c4001ec9468e5c597f497ae99410e92a1ec36308322b46ed13073;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdabe295bfa29f870c790b5e6cfb4ab3f58421e04c485155b8f89b771e3d27eab2fb999a414bc3169755a5af42ddf137c5726fb0d7133c2b6ccf8be06dd1dbed80e33e1d394460feddfd95b10d41af29328b59dc2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h380bef1068b5aff0726720b4b9a61e8d4ec8fdee1cd9196c2a5190c7612442bb85b4dc237e5f7475fb27d843eb59bc14d72d3ba3689ecf87c22c0407a2b42f2a24da55a982d38257227b46d6fcbbf8527275eb109;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67b02cc305057eb94e5b0a02ed9f56995e5fa20d79121e426a17274b866c1348c8bdb8fa4ac26359261c5cf3f7186dd4c18231a3ea3e28ff14851de43fb6f578059d0969eab882222d8833106141afcbd733988ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf0888c27e128bdb697a87eee941cca92d60b804fb2a5762dfb444240ea51aec15ae0d3a3533ed047839c342916403ddd5a467737c0dcc7ba7084b4bb6ca77ad7da55641fc14ccc1a3a1762262e8cac82bc7f4b93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ce9694ed122da0923ff787d108bfb3e4642ab2c55a290109403b9593136f4b9536fe132f001b1ce033137eac91438bf0390a4547ac53a48cb387cbf006252bae701f455c0aa786712f2062d455fe92dc225cefb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25266da0e06b669a64b6de66f018afc752156ef786d01e0fe29d3a6953f733e5cb3fee7f153eba9ffecf30ff43dd74bb572c50f61bfa0c33e0871f670111858816e9eee4116a974f5fa00a452e5d7efe7e078494f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41bb601916952101ce4318591ae2ccc6d3f706fda0640ae6e3ce7fcf64ae3d9ebfed3a7043114e211ca886ec8768d93da980947c313bc453b76a72d59ea054302777ebbc49368258d28c4d48e814abc0d767e4d3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha06b425effcecf8c3cca222af7722a4691abebfef34f19ae9d3ec87cc6c3e4b772669e16da531694cb3d5c9b9675a5cf48a88ab00b4cc2e6c88465475de576f97c7cb43d405d216ba59c1a7b762e5f3d618027f43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd25f80011d354913258ea4dc3061c3583ead816d16cc6ef57b040641f4f9ef6e335465c370cf2d77c9426dbf283ddbe70a231361c8c92bc89a73256acb054e8f836c223343295cf6d8edd118da7580a21c1c0d8c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h349fa75f50e810de4a4a178254297f2d3cfa05ac03582b91f15ca15fde4ae0fca3a5b98fd372e0efa11f04789502e7a24bf39fe653fbc0751d258ec735ccc9ac7e4fb67607b1a35d7f41a9d6ea9d9544011a95a91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2c55bfe7097c45e8a0367f886bcf4d1a70134e3c864310b59c2cd972a65e570502552ac0439d9b22b1de780685a3ab39ebf4a4703965139bbf5c5bee75d171d22d5aba0c75a608d817d78e3769083b25e9ea9142;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h915da6e039f01bbbc4642eb71cedd75b0a484450f3dd0d0c87414e167ef578e3a3bfee77e8ed586982649ec1e502b0105f1c97f3f4f7896684ed42d1e5226ca67861a08826db6d86f759c2631bafa6ec6a8291d16;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87c982c18ff97a52dfe1e98c096c29bc85b86a3e3d71e578b0f9d2be0141b904ee96b2558d97f3578bdc8c85dfd84b84a568d0e399be9704c969491ec1136128473da238770ed5e8b347392108e591f59a0f7c136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fc5e24ce597cf56df296668db62f64af11685d592ee1a3dac78b5db462631f60628ab4d6d5f6d7939bd94cbcacb67403da7457c2a6d56b865327088e5a26216b57f02220cc7123bfad6092c95f034411b9e43301;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ad320f69aa66b324cd8e7ebcc89d44ad54965ef60ffd3acb07635316dda3bacc3daadbc1325b35809eb4ad3716de75bfe51360610e01bee06a26e96b9b5b3675569c69de76c9c5fed7940d7ed4a0f26eec296ec4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he29d88d5d2f396ab17682b3a1a4567406b47ff71736c76bdba25f210d301c2229ee315719ddc5a81933d8312bbea417807c514416347ae41d44e923bc3eb8d34b804736de6ecbed23e028a093906382920e468720;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc34b67fe333bede0923dba6edb99c4a53f57ab57933d10c82ece969950d32806377721549addedecb29d24915befa7cfd14412ccf6cb7dda5843d6b6c72a0685a61cb639684d458818623eeff5cd66da878b0077f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5550c9698b25c423dc757b904cb87ad2a176907c346ce500c63f314f9d936989cab056b3eda21d74636ef3af7c53df0009d7c34f5060a8ead9f3feda0a7d0a1da5f7864d44dd6e7611013954d0e1ac3f3548ca055;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec01c5a092859539269e73272f251e2b5cad4f1e0126dbf39ea165325d69176135b5fe37a630479c35b229532e31dc2c1b0ae240762d99c57ab5b9b745714c591f1e7b7ba0d8cb5fbb623e04790b064e837a63598;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6c7c35c6bca3e45536c0e29901cb525e0a02ce5af359a6022c2bb0ac2fcf951219094c601207c13b704d00d167f70dc91c18bc128ed36383c6c2c25699cc3907e10326a8d8acd515838fca7e1a0a47ca1ecbe865;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb68cd9a2cf5afc60b2f4a46ff2388e2704b265f5de885b3eb641ef650f60a02d3cc46a950d961f71394cf2d4f7d8e98204565d95f468d6e04f09c71e1688447893354c03d25b284c38c6d691af3f4eb4d7ba83682;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haffeefe52f50029e02c73ac0fccf850d59e18635e2ab9e1d0e5e9ef970cccd0097d48b050849b852f755e7e1f556f4aaaa066b7702243c51992382f05001ac22ce5368066c2abbd77a9c34a53c49d1013d37c91d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14229d2401ed7734258b721ae4e72df9deca0e8b7ee49309d82a1c5bc85ae47c01eb5c51cb5feef95cd501e4a40041caeda4e87f62829d25a70580a989d549072e9b1c1ee8a97f8527de3e7070b31a7b84fb2dd8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87cf875a54dd828885933b66f74873f14e6b97acd56786dbbb30bc1fed370d3b0047f66a2d64a7a18ba89cc18493f4c3dfb2ddad52a7b09afd2c8746384f19bdf205872008500e936073b53ff8e614a25b81bf50b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf3c9b47a6bf5c66b9859c3007d010083611a71b533066b9f154e4e3441dac551d07a89cc5d32b8d862d8c110e31e7143e4b327a2fa63c55a17491c688acf747aa6abd6a6e818137bf616a420cc8de7d9282d0d55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha951fa05ea18298a0dc8189c34b67a0f4a013fca0b4da25e28a109942727524235fc6262d5b8d3fb3a86718a05241688f43df3eacefc64b60a667332507eee8f0ce7c445ac8b05036bd67c83b206dd5e6fab21b57;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a8045891e829ea2bb5f9dbf9cc20b4df1b8793af52600355ed671ba6331a7838f2b3be32f7ce0a5d1a17603d810c2d54048bfe9c53c9fe8a9ab82e09c2cb6d9b390f008c46c151e87dcc76643b9a0c066cbd50cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b013b560001601e1dc9e92d0d6af8c8ed00ffa09c9405d9cfaf892e9e50678386d92413a8f4b0e542375590b59b925d3c28e475c28a6ac8e1f71dbcbbeb3285d3f9550275339ecd3bbe09b94f7548a5dfc7332ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b379f61e90006fa6312907005192538cb8015038e46c8b5f736deb2f62adb1791afee043ef576f65ba689634a1134ecef71811aaade56f35dbc2b07f917084c546a7d2d71476aabe537e7eab495907301d7c94b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10ee73a8539d3d57995e8faefcc0a0290347c6d5147f0d72d7d90ebdf6c3cb2e4fc7814fd729276898a55a1ed7b43e51bb2633c4971683b7c4f1656e2ba955dd181d1bdc13a8e5357f8450322d8efe3589c4f3b72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha004da40575e9664b2afe750604902b9719b3a51f147ab9d11f9b78913d55da2439f0127bb2460b5f37cb03936ab12e97f0d2babd01239ef1b079037bb20345c63465c904cbe7b663bf9c223d6b5d67ce2afd0df9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a88e2fcedfdce7eb3c12e457c84c843a60570a07b12055ccd7a5c3a0426792cc5b70bac7a4d7732e0db47cedbbcab1e9d645ee7cce4f9996d454b24b5f146679cadf7a683e24339335c3fff8d440f2b3da440c7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e16c5dfd9c21c062bbe0fea2eaec88d46c95e83cb59c7accd800f492d31655f19c67febe8626a7e3ea2a7770671ea990ad72177889d300f98d9d4d4e60ed00180b4612d2c8d816035576594d853d303c5b258fde;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he40fbb474f2164f57f5a47a262a4b4c7fea758bdb1ace91715fa0c549edf0af7f7e7585397beb5664973e17e6c7256d56735b4276ef1fe632a4dbc65efd01f5f191aa53198aa1e055eb3ba5a85a91c3270e60c814;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ae5fc3cb38686f0a99c684cacabdb59e108e56e996b6ccd638b7e3b51e2dff5632d4828d900f2dc893ce97dd2e9cf84cebce9fe53d0fafc5e1a7f8125086b49b93e82d393d4dabeb1c9cbe9d8abeadd3eb92b725;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d4270ecdd5a7626368e7276b389535342f93df4e01506f97c6ca6f2e9c1dbae35227e647ee82be50aca0267535eeeb89196a25a3e9a1188b05ee99d668849751f2a5b3774689c06c111b663418e1fe00186a2e17;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he173dbe3de78a3a27c5bdf6d75799e2ad965adb63644d7f6baa8b6fd785d2844be2a3139cae474e0f36af19d95b9ee4b5dd4749f466f22469731a8e33d3d0dd5e74d19bb03b7b50cc76f9d7126093f2e2c4ce2fcc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2dd6bb3f145129e727418d1381d886b59611526e4122d91121439fde4843f2b264adb876799d7e402ac73685455f10c68436fe73bedcb4376c0c6e4fc2f6b263150833d61acee811d22433974508cefa155539cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h968164bb5ed7748ac7991a1a749dbedc25cb4e0efddd027c445cf0a40df8ccedc1d19b6b1e8b999da03e5479fa4e07c77b1515abc9caec99232fd24b5c2be7ae08b9e08faa98d92c9d778273aaedcd8ceab824a29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85112762369133cc35728a16a169a9846b03ad99b49d0809739bf74ca9cd87c0b07a577a79a375d411ec34a7b206194d3d5a027af237e47e7cf87469efb5d784a2430f0a0a127573f702b15d904c5e91e7032ced0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h404da0460fd595a1c4e48f0549f5f933bbc689bc4985f82cd828e7b19a5a52c522ef36353ab7710661f8a46e19dd1c5e284e9cd8624612711362ada5a5f1a6cf95082ef91f56d0f32fd79b19daaf1ccdaeb4cc6bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64139e4ab06bd465146499e6bf92d32f92878524985250e33a09a28dcd05df52738222a912c7d8a4df8f6b58cadf7fd60e7c44b310d4029d400d6fdb06d1ca89c08e94dac09fcc5abee67426fead3a2143dcdf460;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2db5488072fc38afd9df909f2cba748b8dad120a85e8fb49ab5f8ba16f1b98aab24048519f1c196186017555f329f6a0e14e79bf8a6214769cf67fc7e9ee8982edc644796ecb859830fc38dfd2c235cbcaa3022a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h562a98669de02a7394f46aa9e87e2efdf4bf23ee91ba91f7f8211f58377c8f4adb40e0136d73b65a20db26ff8119ab2c740f6dd9547118629d61679539b272a7cae73c88ccd67d4d7378cd2bbed78b6659004d8d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfbdbaa3ba549d6924f793d84d3dd4703e2b7af0cab50b7fe51d24e3c3f7096b154fc88561cac27b7af3c2efd0a26ab635f09eb791aad7c7ee2da506300634fff11e2a31791ac82f83e61acfabb674475ef6b23de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaec0c945fb2e5c1a533f186bf7e0a86a69a08d6d9bf10104cab24b87a53e6f063c207498ceada0a91b572dd23d61606c997f61861f7ae90f3020d35d7b8ab508e9a4b2427b1bee37c541f744cf0b31c401e94dc1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc296314832cc35c61c19004af9aaea1ec71ffcf3dfcbbe1c24d5a3708309e6f4bb6ab3b4ade2b6cd5ba2b54dfa1801513a6c8d6c1218f579b18b5774477e5acd373730803d9784cb268aff5336ed5f99eb5de602a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1453cc17bda22e6e5434b99ee86d3f01b2a1d53181238d44d3d1560e61dbbefb9a096d6c6a5ef1165f386d738dbc9cb4e6b267717e99b129e59688f5a257081eeb2fa597b1d19d2aa9ab067f74e9c2b4428e3bb2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76dd99344aa3532df207a5131bf08058a3317fe48d6814a6fa5f3fdfc24e6f569fef764bdddb2a04dde3865c81bec95eb4c2d7c5bff1a07e6ed568e5db1bcc3c6c9664dac0b480901e5f9f8d6c22e6c3e855546f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49fab42a59d31d81fee3435a78c1846bc9b3c73d5d2d06ce2386352c898e4e62504bc7efa24ef96f302877976d7ece965450066d524420bee123f2f3d7691a3816eb9cad9a8a04783d1e57a180d4ac196c4312b6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c3192c0c9311c1d0baf65e3892cb607b144b5e1c5b70bff3e16d65dba32deb7caffc2280e8a336f7c72c9c3660fa23e9bd266772e4310d75c2e3e5270f2f77e642fe4114c84d0ba4119c63ade16ee025b127ae17;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34fa14110111e9638975f88a3af6cee7732001b5ce598590bbbfa94221aee9834d7e6639a1e633c755606af9aa35e9bc80c2d00feac07c0825edce9dd3d14bc27f522217d62ccaeca9269cc8ac829990870bc19af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e83eab09e72bd125742264766f73f99d499f21958bec46459c9feed4e3989e6465ba9cf1797e7c9824eaca3ce1f36d1580f029c6a6f4d4afc4b23ac5b4d7388e46dd78442bb64c3e9eeb3169771a7744f3ee685d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h669b4ad7bde08735f7617d9a0ac3f0d2a5029a8789416fac61879804469bc79a1fab95a31b12d52b18c326ffdd88f6e90dc850a36e471b07966cee2f163b92be8cd86e83a4a6100182c33707a4ff986c30b73cc6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f9a7583ecc876aab4d0340d69a372e52562325bf97ca1a33b8afb2089c5126ac2243fe6c7c041c291ed6a1122434ef84b71c33ebbb28dd9779724a935270bdfbe48da037fff52f18b774996d3b14d9c9f9422a01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h517791c79be57fddacdd71c2679c005a854eace05c6766ea77b4f1d9f0cf494477d35b85d48e44ff29c80a419d439c68cec231ca466459bb8e267ca292ab9759ce07f7473f255199808932b77afa237b8053f70a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd6cbdac851b0b0726c519b2a4e4b8a46478de652ced00334be4228d2763a529e565ac682d4270499da7ee6f54c3a54f487f853aa887d6bf414c4f4ae3bf2ea8009fc242a9281bf5195bac27ccb125c73e2750522;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fde9155c7008a68a98d830b5bf9f64ea82c2bb3c02d7c4681aa90d2e01ae2fbb9768b6ec7aab1526de12de8bbc5ecc35f055a7d0d0d80a64c052bcab6b908eaf3221330fe83ad215ec74d9e726bc50bff0edb05d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11413e9ae992330c89e75752fef1f5cdd275acbf3f6e41579a5c98acff4abf218ba6b2b6ae2841a469c7ab25906df235058d029b378078321cc57dc3b2ff2b3ee6b45b72c5d71b0480c01c5cd71a004b78bea86d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dce92eb820070b4769d06bb0403a2218d839d3d0d29ba693c60084fd68ce34ff35b96fdc18cb72f33c7d2c077bd0f11d6117bfa07208fc462a82d09201303e9b109e693d57a9beb5c3ed3a902eb44aa9e465aa8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he242af6c6024fc1badd36b2e956121ed763a7891224bef8b35f2c461e60aaff2713b43e836eb41d27f25dc8a5bfe5606f56a0d02d48c0e578930dac410045df35f0ac4089302ff0cfc59b17f0ba5de12bff0eeffe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64bb527ccede687f42d698d124071ed5630575d2d4d41242b9b99c89a532dbfd85c3faa98c327e517aca3dde74790ccdbe63acc50e6dd2f2f96500d063cb95715a50a2e3cf247f050e0dd2674a8960c4d34f87620;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2a8ee89d8d510b70c70c82e4ecea11107eecd063510d4b11405b9d6fe5317fcae482d92270e7c42c60b9be8ed3ecb5a6371fcef0ff0ecb358dcc61449a1c9f0b5124790c0932234535c1469ae02106a94f2c7f04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fd34ef076614152c5165e3014fe393190ea9035b7e7316f02ca5f009b700d9b5c6b9aa0647052149fcd29a9a1cdc3bc6bd34fdd593ae814e73c902877f1dc95176e9237e08ba64e84e44d72a9946cd3eae45e56f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c276c14f1bf90ccb32feef1acf8960619a15ac94664e293cef4963bc1747b76d22d0b6909c767508c6cd6c6aeb718482f52caed2a62c55f953190d47b1feeaca1c942d91b2909bd64824b0342de2c0ec5f542839;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17d95281eb9e9f1a3d6211c44c8bb98cbbf11ee8749966844df9494cfcd1a0918d9001db9e31146368807314d543d2b49d64f14e4c0ad3e78e38bbbbcca1a6b7f8906de9dc087ec8ed01506f0a9fd762a59cc15d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e5a1a32b22cc377b782a7e434865743e45fb9ea9a4632468cce58b640d19ec0e9be813e10780009fe997d026fe7d74be7d913376d99321dbd603969ac333f23df9f2f5de15307f6c3a1f914482d5f8f76762d1dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3aa9a04186555734b93af6e7408e4ff9607f276b4d41c2a4ae0e27e9b454aa7d1db72e4c2932182969fdbfde338d98c0e0980f788102b7733a48366b67b443028a699a867a0082c36a296e2a68783ac6d7c64e9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee495df76d7ff339170fb7afc7faacedb6365d7d933063d37e64d4f0eed3b8ae3adc56bce76892c958180141a7f24079c74ea4f40971db303180920907998a4ac142373c3be4be8cb221ea4d20213211d6328cf25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17fb9a66af5826f09b65ae7ad88c775fc6cbbfb8c58b27d91fc7b0a728c15a7e1f5507fec28146c2247aa61d9fa069c9febb778d7ceeedc861805785161599cc8e5219f42d9df25e690b15c72cf4c4484558cf868;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5403c9a2a7538781e212e30704e168d4824cd6838ba37a2167190ea18be118fe63502835fa24c9de9e6b01ca9055d37ca836e07523200b82af77c239075235761fbb5ad1aeccc3f6442fa5ae779e9ae2ef4ea83ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef59a51ec23bf62c03c7b4398f02555f89ab9eefe1a665a3c8d9877a83610216163c1528d339ef86e97a3cc4dab3a295d6cd4af72f2f279cff8b2f0a714a8070fc74c3f5523e817e1365aeb0d5cc909e0bff30a90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h992209c1d14ece282406bf9cdc8e8310f81fc7f21d6806e22d0c5e7065c94c801f9d2a9995a90869979a709a1859653433056812d474454ca5f384234a64847ed925c5149ffab6894265bbfb34837703f63fe524e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h940e6cc4a5f772d3c47b0a929600d07c5b461734bc256b88520d5f120c87b2487d5174cad3b8ba5532f9735f250db976e21c7d1ed946e7a1be5281e50c6ab0e2a5805dadb2e8f2f5409169ff46e6b6da3f886818f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7941d0d319fb3aaa940e264ca1f3ecffb9efdf32941c3d5903fdba7727bf6dbb14b1ebde495d3a9e4259150656224c4a088add2db029f7e5cf93b9dd62d717bd7e500f95e260691b459638cd6bcbbf04a332da41d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6af25e2336746b0fa565037a7caadd2be4d6c497163b913b618eaa92ad58c1920869122ade06b117581e930d06b46e55e9428d8c48577ec080ff93afc81510b337326070286967b4a05a12b6ab813d775fab8ace5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2968359bf0cb950693f7c9fcdae8af5748c4399edb28bcebf350a2d1cdf07209c4561d6d040e83c9d8a952de923656885bbc16658c6f4868389ccd2f73328949425a9df6837a8d6718548f3c0b24cbba85343d77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h980f65be71f9f72568169bb034fed1ae55c77d8112c77c478e800de9a6ddb93be447316c382841002efa0f9025943ea7c0aa1871a1cde0388fbf0e7be4466d41ddbd038e5b232a6d7dca6dc8bb7216054d257ff7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h414badd330ad257afefd51ed09db1cd6ace910684dcbac76c78a0248d6dc83bb9f4a4ad1de1531bc5b9b273ba531997d327fa250c8ab6035932a8d484b0f77cae0104565936fb03a9c8d8f77b078d494d8471394a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e09970d9af5553b5290c83b40cb397d216ade1368e8e3e001bdce3769dc3d2be20fdc5e9e96b7531cabdf8f45f1b33cf6561da1ed38757232fae800cbfd2ea678732f5f40829cde249111b5086589af420e0c7be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2997b032cebe493fe912916ebe9da860e48695c674f0c9a8cef451d6ea5736bf73167a649c3da2edc2653c57a6ca1991b89ca7745e4628ef87237d544893897d559855e07b28e07bbf341d43d209c9d50b6f98b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf93bbf7f6038475e0b454ed70e5d460d905f066e8c4c19a6c998de2cee0d3030db1408a6f9eba44283853673dd329eec91a2db26836559390bccabb1f2d1be0df96dc5aa0c3dcd9e7467e32e59f66eb0a0b95533f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33a3f0295b75b24107e0d77c23ffbe6ea669e73ba38e48eaefd103fb82c29f423bd9ae05586ef20879425b94752a50950f68fc73b8fcd0565834c794063f5fd374d2301672b34a5bff1a56f28bfa5f620151dec64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3794b65cf76d50f43d65e2a23ee6c834971c481520d01b017fbc7dc7f5fa0065c0be7d0e5b06abe1b9ade91a0533a463c97b6149bed846e55c697e80aa8e9111714d0696b0fb7d2ad3236e5b494422b441ce67808;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73e01ea450b57d66f61a3a5a73f5411c87217c23f5bd09a2981b161528a149a524dcdae6cd116cd355aa7756fe1055a1005ec21e7d8eaf8b88d55a3456959a58df80386e081eeabaceae1f777983c36bcd88f3c28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd42ffe5d477b61a566136eca409275fc953b5eeb44580724f1a5a5887aa1a91379d8ef75185d823e14c5aa1d3f287092d25ab06045b2019bdbac70e8921bf250926b2de69166e8484431e90a452cfb33db0e40d5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d908fcabb9de694c775d8d20101f53da6f14046ead4418378dbc76f11d7ef783dc020ddede6a515ce3776e94dcdf28349ba0fe9b200a9859f15f2b7aec81f2d4924dbf41d59de6737bb4a90d3579daf7979cb31e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7a5298f353dce13540a4604c7938b081e945a556f0646c75cccf0884aa15a2ffacfb154153fa37e606e154b11857fe044fe161352e12dad304de718a66c9d75c21817adbc0a4275f27a6ada34c5d0cb64b5fb831;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h481e4546f480027c58be0226d8990de35a0acbb2523acd68e522f70842aa13c715baa1345218350e938be63c2de3a0d60fdd563ce8ca17dc90bcc953f6d67503cb542b14d4320ed7463304163601c5a06e7849658;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef5a23d0bc4314fe045a36359713d8949165789f524eba41c4123aab7f4e1aa6cb1fe3479f367cd7a2ca1e817704c24ab415ef2ea226ed730eff0a1fccd50708311f872bc9986e5bed1b9622bec5ee85a1aff66c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9410a60bcc6d0413ba5ca0fda12bca15e24f69cecb245ed30721a308c7ecc9c1596cee691c0f3fcd9f4ac974aabbbb4731ecdefe4031b2c6dcb091c04e47d8a8e45f66704fc2966c086d1423bf1e2fbfe067de281;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2916a8f026b18da57782fc04979be3097ac8f9529b45bf501444068c552f92b53fde793f4a6980dc93c768b13352bd4cd07378825fc3be88fcf7cf06aa25a5d37e1a9a7db21fa78d21096f98fb59841aed88469b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479a9bda540506741f6a13db1a60f5c0df18ca07c6ba39b612cfb493808a8add63993d2509d09af0fc0f9894fec2b4b30098a4713073cd5b50f90e4089d9d4974dd10e0c3874c03c5593c2d8641dd9a1546bebb0d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c967af999d00b0f94ea8e41042c54334045d13265e55a40e4f5f561246d9a16a0fec2f17adbe5b1b93cae74ec8a443100b16bb18abd7ea335427e2ba3679dd861197e91c2bdd9a55b1712638c7ca30f4fe9a93b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc84f4d3c57562387854140d8be294ebb06e686b6c65c1c3c52cba6b47440fae2fa9bb6c2ff3bf92e93e5edd2b0174d7e8d3e0af01954745efe663f8d1b85b763c4b0ed564f1f0d1422d605122dda04c1008137ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha71d74dc6dfa3a3aa22dce6eed0b28cd07eed05dbedaf9d9e6e15416c7c5694fc278488933909d386ef70568558dbb27759f20aac8f0b413d07db1b84855e62e442e1c9611cdb1128d9b98ab5b69009549a2eb1d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc38c8855b3c4eadf8c62a3ccdcccd83df50d5a9ce13d4833570b2f35d824ca429d9113c9286ae792e0e9c1139f6509e29d0b0cce7118fa7e5ecd55f360222cfcf658846142004f63b6b86862c928a80de0c3a5c8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ecb7828e65f491703aa94f8566ddcdf4e935d555443fef16f2d1e10a812a97cc6948f6cfba555e44589f8a8701bb8b4ff7f63ee90023244076c92aba43c01eb38005d8dd27a250839f51c2c5cd51f981bbec2fdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h784480bf1c377b4bce12bbd129906d0b61c9a3eeb43f0cdade31405c350c5db6476fbff0441e4ab824458b25a1ff2ef6eee6554bfde7fc69136bb94d0cf7d5691ed171807fbaf7ec2493afc6b7252fdbd463fdb36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb67e07df8e713d0fcb4d2fe3250219396ae0477a6279f50cffa7b2622babe04563bb6207c3b8051de8d489086a0c47669381942b269528c6a9fc3cc95735ec05a8031d083fdc404978e03bdb6fc237bda61b366e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41ea581b45bb1e02897ef78fa8b08855f62c9b1f2d3ac5554de709d41a396d2c0d4ee7d365d5d7b1317c445d44a82ecde3294efc5c5cd9f94c589768f273f6b64b5a7b1ba8ff1f13aa4997dc499180bfccb5fa027;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf815e18fd317cabd592b92d321fec21a4fc5590c35e6ab61375d65b449b3e2b21e16f3fa3f4847bfaa83d60ba3025594650c80aee4fbfdc1dd7a69e2bedc29fbc41ce8208f87627cff032c0578cdbb886faed50f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c8a1b459a0879d786b6654f8a8ff12d322b26e0f7ebdfb9c9db61598cf1fe856d0bffb7b69713ad1775eaf615056d33f8c9c5b379ea3084eb265f7975b8f458233ddcf58c7e3a094b733b3e71902e15f8bca8a99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h954ffa590cc638c2bc53636f2cde9a7efbdbd3db15890659e9d3f1d75efe99b1df70aefd226ac63168b6461ae248bbdfcf29aa55cc20334fa682f628bc05287fceba64b5271831742a3e83fd66fc0ec8cfc10c856;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d5255db4b65e3ffb133840db3d4ceb736a39ee693154610982dce207388e82182b3c252a25b595ac51c92c9c202ce005c7b2cb8567e91c7f1c69ed11662e3eeb4332a593dddec17e9da6ae7fb0dc5f50149e6ed6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35bda062f794420d414f3b991e4bc87188919268483b8d919803b803baa3c314b7e8a5482890a53f546f4c369cc9c421df251d633d56a23832f6195eaa79c24711a7d32bd1ac49bf07185a8f5ca0ed6155f64595b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h535e9e135c8c6cba65302b540fd051a5b611d3e554018e04637df304971ff0ec9225c73c3ff7c9981b2900614af8aa38164c55b875758d5923b5644edcb1b7ca6c4c46c9ffdce9eee4ef08d6f8ba0ee814eb91f93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8aa1b523e3de17102766bf9f037eff1694b0e9c546b6cc85b960e614bc159bc1f12a3c325c6fc72483750681d92a40a95d3d998cf7670cd4e122ec4e9bf34350128b89926ea0e2467f48b3300f3e5524c4ca7498;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee285687f31bb0580a206c17067556aaf3df69c35fb76bb5742f423e9e82f53e1bf779343312436b45d2bd0e4bc7a58381d6556967711a231cf004036970292539ff6e3ced177b014397bbdac4065553f3635b15a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3e6d55e77ea5384ad20a7a50c93259dd1fb1f85ca6ee8db6664e31b1c6ffc4c23e62f1d6751f29ca8906732612b4016de571c9ef7823f0919724ded532dbceb33fe5366b084b4ab7efc97c19843ffab3abf0c1ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ffe7c19a010629b1cce1c5fcd3a64d900eebb0d46fd0c039b439dc23c721299663870cb465561ce5c6dd09f0c9a90f4f407bcd42ddf733ba781427d6872c8baebf112ae7b5f7ee1d3b1170cbed95278e906749e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aafcac5f93cceb6303a5437527f628031d1dddb16f84dbed3688307373fb61c5152f50705af31be1ba6cfea71cff2205fdda8a7a1a9ad322742b92a267812548a86d71f34ee1b59209ad01122a06e8ec7efa02cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83a2dbc555edb342572a32918e694bd2df814be453c1801a6057a83899a0199ea4da3e703ecaec3989f8b325a12f71d04d2bef7c735e6da3f453c3d181e50bf9f74fe5c8db356e4bf2a12d98db9e38f0b63c7bd1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4f2c46e283076eb6a9d7b5f6be5cd129b7175df39c4a032b7edb6b46eaf1aaeb11f2329e0b4b0912b1ab00d4c1a01edabe68ad299d614215ea90ac8736029929dba1d7542755b07aea7927bf7fb6318e579a9801;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h657201a587f76777f7e1c95b5c6788f538a20b449a42663b1eb8bc7b7c2a959b5e5c878bcc042e0b275a0e56767562a959d78ee0f9faf9cf14ae49f493c98f535a915b3ac2ce95ad351269ad215f57bf4f12acb55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb72690d7703540d26a758bb68417cbb25b264286914a781437f5a7f68422b7e7335aa5c0c0b302f7ceac746f03e7de32423c8a0df97b9691f7c2188fba24121088d4e5e4d4d9057c1a9f30045caa961a6e084eb6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1079f03ab4f24b90eeac5004196d288db803b0b1a211e526cd3837a1d6f22b10194f17af210762a0824bb0224215a41c273628a24be516049ee762cdc05f38cee56fa9dc5e355af516bb3e4614d3b14cfd6cb92e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7172ba65a649280470e501670f374751e29f02963932dd7dedd2b7eb1fd898f755be18d076bd92f5992c2f48236784948d3a1666ca9bba0aa8796a83367ac075fe1e5e8daab2df96bab7b419a5032bde1d41d5e68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1016517b7a89aabf569e1a155ace49aa3228faade752c636c823d087c2a3b0c1cbc15bd68b578111dc90bbe69e04fd4a9d6a98e9fde613b3dba2b796d3faa8b2f58e6d162f25435cc07dbc7ad77c22414256c0de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7312d5b7f12d95944ea902fd95c88bc4a093312bdd733fe755a8d547fac8ccd504ac03375fd69f9627ff24b62d54f007098926b18e6af84e1c33c1cf572496094ef86617e05b9b12021204b2b9d99d66cde59917b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4e3c244ca523a6246289272be965dd24b2b23c17ed6790395b57483bf97855476f8e5c4770eedb93500478318cf8c1537aa6b8c2b84ee48b077d340461309cd96e7a3d0fc4d924ee365d9cfeb0fd11838c589a73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d1a9c88468fd51064fd1cb858176641665109023adf1a8007bc465c4dbd62d19dc0ea6d3add55bb392149bda0315726b96910861a06efe37a06fd8eff1d1653f677ae95a285a65592a1d9189a8a8e2378dc4855e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14f8b5a92d44efb8d0a5ad02b31dbe7c7f330d7fa772688a73af59be24f9c7365cfc29068bb3e8d65fdfd86e4436e8192bf9b5a0c01a6d1cadc0943b018ba17f10a5a9b498cfdf0d07888375d6cdc4314afa23b2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37f06069d537a891f205fc0ab233022603af6ce4d23691f95cf502a512c0ac179c73465294b6c20fe99d3af81829bef4fde2be28d48507a6b689963d2dc7f589905d91cf41c5b957c4344d1ab4b8341b53083b7c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he72c47c6e80c4a27a19f04fd2dc7f6c3a83569a440fbbd0869658f9a46bc7937269e4594192677c6238ce66538355266ef32979dad67514b845ceb4119f4ead165d0d74d1c25f5744b0395693259b065f67211a00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e8ff3bea95c020f5ae283eeada0f3015dfb6b3f90a8ea13a421503a2bf29862c1b4575d170f74e86797c28ea076f72074dbcdb29dce2bfb79e2dcbb8fbbf9aead341d88b3a1afb41662c849c1e3b0b0cec459342;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12867fd91d4c55ecdd5e2ec6211d85e268f60d83483a37d9b388487b93f73585ba29e6073db08a8744ddf1e98b71a6a7d0c44fdb20f28f67118ca1d6a9d2433d8302d3d228f22b54a7ea32795de8589bc2e2793f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d60f649354d6007fa77cd15f1e3a683c2fb66a4fd1b994585c8889ba37f950b6874fc463de4e42210a5b8372cc71025209c17b702a7e69df8cc5c82ee3d68e97669318992b05bfc1e862bfddc0ce15e8001d9ee5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c64af19e67f4cbc6820ca48a826a03ab6cddb709ca3148987606d4459754c48c9e3c6ddfa67de9d792b23f72b3d8bc89a68807082770f59e45db156067a0637cc8b4667427a05d84840f458961ee83abf4dc2324;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9441a38aef17dd9d3ea791ff1deaca61d2d4652a7dafc1a929ffc27ae0e371153365358aae018f8c4e9071ce997edc3d4ce478f2cacb496563c34f8ae7c70bb0b7ed68ae268dbeb3dbffc8a7fe67598e8155c8948;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4929ce40f58536dbeb598b803f396e95e74c7ee3e5821e774876d4a8e8de154af040e4e924c18c02e423372196a1c7d1ffada8dd8bd6d5d7df70343323c27c77288224c15f0e64f6077ed60d95ec87390f360cbb0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e79bd083ca0c7dd17f2b96721a7fa00a7e2b05b322d73418a575ad7aabfd1b9ef959c61a21d21a51e885f915ab2d95355ad3ef4be09383531676acd1f0970cf1329d37150bc7a156d3c9aed884c081846f5c666e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea3875894cdf42bde7e74cacdb949d957b6b6b40f6eb271b5efe8ab160cf1f51cd288dde6fb4effddc037f14e6ef0b4420d0d48d76bd6dcf2f8ffe5cc94add80626d6fdef16befe3ea54a61188aa1cc40ddbd715d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e0d734c0668bbb0691d9425ce19c803fd7f19013dc0a6584254e22dedea1bafc916198b6b7469f0ab309ccfbbb1d8f3012c2314bcbb94ed9d177378960d13e1b5c3828433ac59d686e4ceaa4565cf3afed45495f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3fa55b5e8df5794b7f4ac27ae34ad55a28112ec213be5b79cf035424472be9f09b96355831ae64f6dd2bb77cecebcb4edbae942b544f165a1b506fb6d434be206551809071fd92bbd6fd98702668a1394a28e52e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dc44eb28398cc8b510b46220eab6483b3a529fec8d784b14e6389e273b7520ec54ca118d6dacaa2b2c2ec50c68bbc7d7d96a31056419837c13468ea5e16061b6d66cc2ae8838bf8b2de02be82368f9d5bfd9a473;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce1742604e7b6380066ddf62582a4122e6239daeeae3d87ab387d444cbfda38973a978c3a579437675f2c7f22a05e4293730371d321a9b5cc944758af736813585dfe9f4b9750f495250cda024e66a20ef5d49064;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1789df74b51cef81bd829a00532d2f54af1ac81ea010ec3965e29c631d09535fc8e86f7eb267f05c2e9622bc556d351026749a02af12722ba17c19cdf9111b3dd885f6f8459989d97b0650178d28a09a346393d20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h848735ea106c6d2f5c08028652f31ad077aa8c489fa1ae9bd1554c69433f09d84807fe5ecc6fc243dfd1fe4ef43f9255dd9f24c03b337d9991f82cf753beeb9d7a092a2f3a0aa715fbbc77488c832dbf6fcc3b45a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dbd884a908737841d7c00ac4138bfe7a731b43bafc689b48186e542cebfc079d0b9f97b327c87ec0b2563ab2e9fe2e22d47b80a4fa59d15f422ccdb0fa1c816febf010de7c1f0d89c9578a497522f410122a2746;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38bb7b99eef44be9a9f77017836058b31de40b93ae7b06223af7f3ca5f05009fad9be9fe379591ce5f10bde61e52d58c3d2491876c681797e3062cd4f73e2cdbbe951ed2d7a7d19ce4b060cdc20f829a5568f0b60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he69ec4f32c3bb0f9a61b60024522f57ee19f93ae4dd9c354d7ef559730e20b0331cc5aa17f400b3600821a7ef43949661fa8730c3d0e3f63c683580fda8f9bf046adfbe99aa8e79212e12ee903da08e699bd90754;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b4f96d98fb0cb807c3eee2b16df55e22a0939529c881005b6adc1819a83bdbc8127d5b0faa58ce1255969abf9957a20f68472423a372c26c91b1e35d61cc351f7b5c9f5bdd6b7adf10d45f2091a04e9c781da984;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6034a3e411366c1f99eac492d226ec631aea20003bd31e125dfe71f17a122e8cb4aaf8b3a04ce693d764628e845a38d5770ffdb70641231ddca56f0c58bfad45a28f66aaff5598f1879e0c8bea49e5a31d2dddf26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f41d2fd3c22ba9b3b7a7ebe5fb1487955fb1f7a4f30382f65358cd6c0ff7e357b6d56d531b4efd781e9a52db63a733edeb40cabb5746163e2a4926b3c34b6e05e247cda0a2e39e85b3788d1fb5bfff0b5ed16e7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9036124d01830fba11c58b15537fb4f2e04a0361c7aa6f81b2583cebd9cd54ffbfbedf5ed02c1f17998c43b593aea2f1d565308a62f2c8de4832c80065d1f5b291178861aca59d346db2f80d48ff0e3735ccbd042;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha88fac89357a5d61e940da9c78ed871a9f6e4da8b6626d534237720b1f27cade44d7f00158bf8544fb54f399f00f004f324ef7aa167577e0079016ee2e238b7a062b825504eb3a81bcaab420e473ec836ad8aba1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc660e28fa8504627077de0d33f4bd0593a368dee7b5f6baaa26ce03669e09fdb4967ce5f2678273a355235eb80320c8967efbe95943a64d9cb92f569d5b4f4ad627008323e1c816e7b32eb5db96691f6f56e191c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7002d482294b55349ecb9423546c6a562b48560b4bac878aac8e8880ba2ba18b82c37cdef87e550ef84d30a26990baa5ac966d91b3653d6c1c07bd787813e87894d727e52743907b1e00686e5b14c34b62fed362;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d30f0add2811bf011fa4de4d9eab709a21e363d40e402080b6a4fd932314d25480f3c5af2604e4469aee5c92c4c2bc43d3d938134ca105ed308352ba43f0aaf4722a3c18e5c17ba0daa9222540d79fba0e9de25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h523bdd69c9b2cc88b321e863f9b3192b35e06d71e0ff359d1d27d764f5516836d854f2bd8952425cf4693e2fcceae36e8f6f52cd9b5894e5281313c5a3093afaa7d32da7014c68d0cb979c6e9fe288c6622146352;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16561a73c0068d9e1e27ade6565d9d450c2c8b1736d9fa191f87ca8e1f09c668b3fd3ba4446f1f71f98c8ed4c2f9a73188caaa12f350d0a5d36beb1ed1c9a00306eaaf945478b371d3b2814aad8b10e4773f18d9b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5311faa0e04a97372babe4de022ad54c34d6cb564bf524ccbafd5bbc12d4fd398a872ce1cec40a0c7ed1ac59ee9338ed62e3a73bf1cbd13282c4cf5eea4c3bac5d52c3a565d9addec6b6f2fcce9991604d25e6ce1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4947ed3b5a60df04dc06491035b35f63e2a45b93b5872894e7aa5acba80d029bd07c3b0fe0ab130ec1335130d26f70773bebce44916531a60ee91c399bc6a562dc956a132fe06e26464b90cfbe466e0f519eb89e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6540633a55f200598ef79d2eb85e1c1e5cd89445cd75cab5c18c86c8b2afc6d98972500817b141084c643f9ed820ae3493ff8b664b2e20e4c2791cdde9f695a62b8b96e7b7ac9557988f1b9a12ef62d7a62c0f0a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a260666c43bf27f1ba702fcc254882379c9b80bf38379d0f9b4398cf6ace1489a5da18d525c68e434a91daf5b6fa0665dbc3eb03e6756f7535f259d151ec5dfda8590713e42c1641a58cc5e9dd230abcd8ec9546;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31850bf92665b86a334fdc5f6554c424c62e2e323adc24247ff4a535c778326aea233edce99895fe5a3d5f2c74a6556f66bd80b2a4d26a84bb5e6f53c08c53bf7b06ac4c7190929752bca847c17e295739da4903;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h226648377d3cc6b2d0f64aae6a3bc8fd2a9a98457e7df50d357f3dd85e20003791bc0977f08ec21e5c8ae6d1312770ae6ee1804f46e4232c443a6f4065507e33c819b5c6be27943b17cf47bc7fcec672169b41c43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d58aec83e03fc7a479e97eec347a44d65d5691665890c0c2ff160a65c88807290a5c15c8449fe2d655a2bb38b357e0734d08872e3dd56d7393e0eced93d1752ea3c49c13f302a640daa10a293fb49f81697d36b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h582478abba2254d98152b7d2a291fc0af10f058ba34954edb98853272eab0799413479bde2444bd09d694108c9ada9faced8b2cee1fe350bf8327295c5d7268bba46b6ea16772c77debdeae7caa84cfab80d8e8d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a0bf132212aa3f63b039710dd356cfc56edadb99511d3e444042bef525fa97d59a8414afe30e5950a3c784b8de0b319ca309067fe38e4bfaabe888621cfa69f5a7a1a3d213ba2d521be5976277f9947cdcfcfa58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb438d81587ecef623c7b80e60cb15efa6983d84a4f99f5a9d87db5bc24a7fbb3cecccb6a81402052abb428b528fc24fd825a3da4a2ace9d5155513ee74224059a5b5b53c756800f07c4c2789bab80e539976c79fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h148470bee7009f1da847d7b69388a9a31e0119ae02420407f3f8428addc36d28d2dfb26dbf62fd924cfd1deaa9b8aab3458f5df42cd795e2b35dc24d2ebdaf8442c8cde161085e9910d26dc9220703f7c29d51db2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc239af80c3c2f94b8d0768f69a43d0ea2f335646bb4546b6ef028722da9852c753c598f4cb90d540a7564d3b8fc8c26b47445494ef6cbb95246920c13055b678689f7e44587633acc4d0d4fdef357b59dc67e9662;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2d718869ba0a831b71b97406b96b19b2d2a028df7b4898cd292028fd485d5aa2f302bc0ad61e9bd26d0c9237182701c3ac80d7a75995eaf2335b3d10c071848fe02392814abbcab2b7d0e37d48af8dea67090424;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48a4f1b720223300ec44747b15a5ea93d2cdd34401de3b1fabeaa7124a242ede25664586cc81322876bb4210d1f13074d84b3df464e084cf37f20ec4f40073b2942494b66b77fcc8f52dfd4e47b374ececd181335;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62454e3a26d89137c3176f8fdedbf3341b9dae5769947f1884e1679ffea194ff7992b5657d47f5f90b7c38b404329a0fa59122c225a8effe7c2336918217790edff5ca77e18e1ce515723ad29834e4278b34edfd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h628a52a38f56fe0acb899b859eaadd2784db9e9ddcf60106aa70aa872b5b50788971e84037f6f36bc8862c2260b91ada962f73a8ad8a17e68687c05294e3551cf9bfd7d06c921649aff67d00c71e3db5c847214f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c4e92001a2df461ce3f92e579574f69e1c09bc95c64241a0701bf8e9efa1b3a0cab3323d479f9a572b287ca640db494e5776c9ea49cbd939935b691c492ca63aced139e96d48cd34ce6170c90e58374278f7286f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha781f85d0204a55859fbaf301b8fc80cf88bc25f30cf267f1745f57335cc8e8fdf38fcd8eef859827d8679d6103ea2386ad3db8c89492825b04c2a1836613b135de807ec4d936ec8ae93f839f6cffaeb7a5ed14fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35a449ebc447da69ef8311bf2ac942fc79c3baf698a8ba9cc41c420acdc6178c9cbc62046a3d661eec2f6e01d28383330cd1cbc0a63df7f5546383ca7385df12bbd98cd9f242e71f10623289852027bf2cba4c55d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf87ff0a9f1c1eb605ca4fea9213328e068e67ff74f0d53e0ee590aa01398f1a3091d6ece94a17ac4c7a0febb0b93c3e6b40b112ae939e3e899cf65e3da5cd18fd5886144d909fbdc7540500917205ef7eaa66d1de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7b2a3c5bca0f7aead5b5f73d1b570259ac942e9c35a118aac7b3a11d5363ae57853263423293a34dff1ed09d669a311a828dea16003f12d3e46ccb1d66623ee36c78309d3afa599739cdfb17477d2d5047a9f411;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h889836cde1a7ec557fb2aff1acbba71807266bc3255305b8aaab0321b991c349e87ec7b73f139bba20bcdd5ea064b49453d859bfed690773ab7d8582e05d36665e722fcb276e40717b9e9b9027e3851852e26da85;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98652423d0116f92b90f67aa90b8d3ca8ab1efdb3bdcf3ec94dafa6e270be284de4fd765a907412f7455d098d3f0fb3530d9d5d313178cc52d42be9e72b65b4050c50e646d4dbed8d7d054f1df39e65d922b3156a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e2cf25cd76c2226ec8662e3b8201779c32841694708e24375f128965caba270e04e269982facefdd454a4215bc9f73dcc121a9bc4708973281a6b2ebc58b013908682ecb6c17dfdf21b92a912b823dae5be90bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f3b48247a13f1ff94faa107459402e87c60e6e36e4052ddc1fc76117fbdc320fe2d9c408d6113fcac8b7d2e26e7164329961e0db11490a4a030aa22e6c9492430f97e4936f1efa0199d659c8ad01f5654670de1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bfc0ef53424bacf0602862ee88c0306994d3f381232262227bf9bf64d8b430b664738c3680d95777296548e4d1d145daec15f37f775eaa4b66b2efc4e61c88ec50559b10ee201acfea2bd3bd99b0669d18dcc3e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h968c36b15334e2c075182a304464beab7dd74f0824d828de8adac26f413e127c6ef344608f8620788762acc6fce737a86b99c16e80c292bf048ab6e23d1be370e0a1e1b512a619016603d4e18ea581237d8397196;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44a86e238e53feccb1b999ee403e7492ce22f87c5137c592d54b55fabe0dc677bf9240d614faad29d5d4939cf578f54272a13e60def4a734e0b0341863cca03080eec4210724394e1cfbfe6152f18c09c5dd2216;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e899fd3a70c07c8f00a75785ee63cc5215c52cfc826388ee5ad04cf38d89af1aae9dad90d870edf8fe3fd02932726e2ea9df41744fd6857bf44f311390c7d128437c0c9b139bfc979da1e4aab918417108751577;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h811a4f499e7778a86dfeb0a4a0076e1cbfd45535a3481c469d5e322c0c0c571bc20d9bb35e7e69ed443a35f975ce46238d5df3a426eddb6ee214604a165ced94b9079bda65cc8eee3854c2737eec5c7baf3f2d869;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4db2e65f78e25ac0486bf05f59961488931dd13fe1a8c6f6bb59421b2dbc83d3d70d36360985e0587dd13ece7c23f3fefbf8c07f289c0c65acaf13835bb686d9bc42768db0e1c33222ba171b1417506e2979eeef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf47c39733ba1ecd0b71dccb5bccbdacb3788e1b58094923ab9cce1da13f9cdab086f4db4e84e4f7c4e18a19fcfb6249b661551177523d2b7bc836dbbf5fb6ab78d4a90dff8a908cc953089a02c3dc001e25b43a38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd60e7a5d2ee1653854ab339e22b7a0fdd9e8557b49899533517ed822c96dd78f1dcef56292bb81324ef25d050da9b185627f47ffd927ec4067dabfc318d65ab89a5568f9d827f1a190c7a2f22f1dd44cc406af890;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35873a0300c04eaab80b1e8468ad7c9e7e8ee6acac0255965808d62b76acbfe650c7b7d51027e12bdec497b346046a219040065c9fbb56c80e50367cd56162dedfab322a4bf0149478e10e98d7f2abb0e21dd6d5d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4aa4f52cc7cc719ea142fafb9437a0870085480f80d3c97b22b22a760c2eac5692436af72e236268df47f94754501d3b7e7b5873ce3dfcdbde167078b78f7bf02ef363d3be2458a225bc306b4755c42b805e6915c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1504b017992d34048cdb9066c7153261206b47d393c8ef0b65419e6edae1cabece5ca86783a002f6729489a2820f642c8d462eaf0d15baf83eea6be3ff118aeb0f974cff3e809c8e286b8da56f60c2c2c0aa76610;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8f8e5d0b8eb85a8856314af93ec27edfde802c8c173ff5829ce84e54dcb4a9eff19393422075d11382c2fa83f9ce2c36f6a97bc0a648ee7659472df841d95bca2381f589af142c2fa45b90595616af408f15daec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha69d30cdf804dc0f581e51b23fc746303f9204a2bd9ab0569b1dc22672fc54a8a4f4833e23f3789cbc956a6f76c92cd4bfe6c20b188f674d14e29e9f348a3d6910ec1422641d127c4434a6b0fa8c4b5c348dd82e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h715e9859daf8c0d977251500d3e1036d67baaabecc6adca47977e4a02259b9c831d76951781525c1c9368f2f8531e25c7dc6ae36817293f2dbbbf1b37e985c6055c0d357ae6adb2d7de16dec0f1ff7c71669cba32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb50d56ab1f154d41468efe7a0208a1dd95877fd9c8f804127e0d0c5ceca3506b9d2810c6e3e90f2d2623a7f1aee8bb781ed3bfda9e712cf20988f6482f6e9c4707d11258f86680e59a5a4f01671e576b024663ebc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6248c6746b50867c2289b5e938c2f3cb07b0a38bf6c5586fa92661bbbea5db6f926cd267f0acc2570e5178c6529fee148f13d3a7b5b3bb27cf15083984c76b7ad4ba264b7bf994389a12a5f48c567caf78cc1baf9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f22700f98ef7517b4328807f924d959b3d5308135c725203a8d8f2e2d3c38841a9b8450505d057c00eca1e833e82b8870baea07c0890bd5722998d752d818dd4b2e5f529afa82f64628c74130cd065a03ed7f6dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf85fd6ef534a594ac56b781d022570a4635e72dbe8c5add84f3ce2b10489317ce2e822d6c19d917af635991c0bf6d72c170c523a89db31d95f89011e7f705e5813b436d017209bc1d98c80ed727e790aad22727ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7b83f5d917fd61ba03800a255563cb22474bcc8ff8a3d941317342895e3ba9e711d5a7eeffbd2b49fbd78cadaa57d4879dd34482b9483ea1418b13c4e5810588ec59b23c68115e028479cc3dbe5dee32d453ffca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd96bf8c51cb818bb5fd2e7c1f273280435ddfe46c352dea4edfefbd32cd877c88146b528f49824ea58412445086b01e267d24e17514035d6b85542ecdc2af64f9114e805466b9bda73b2567a1f81e2230162cd07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c36b47d40ebc97d507c2fc7a2eca32a7c72b26466c7e034a30b3d7f21f8a860e4cf00ad3df5baa3bbb684265ecd5005c80baadb7db83ce7bbaab4dd89450d158c1b787fcae0dff53d54b21c91fba9c2acc26ba28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71d58ea37e8077d082b6628b9b2eda1046bd16eede306ef9d5491f50ca05e7cee7f58dcd015c019eec946d7113811c9ea9d8c648f8508a3d713c2574eb68169b9a975a18084b50fe5d9ac7427c6766e3c8ca7a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2ee0368b9c09676b84916f8db668d0b0135c4055746a9ce2168e81922265ce715c45bac8ac705e361232ffad823c848140a90eec1b221fa157f8204032ed177e2c8443d0321c1ad2a444e0009aa5f0ae05aed112;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf70946a2ebb35d93d0f8874a60eab5441525fe1a0f7dbe16c4863f4983033586b1f563e9a4424ef028401e47a65e8072f280e9e4b8e2b5ccfa0d81600430660bb8c241729d7d51a85d06a4c7836f78bee49df160d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38ea13a5dbe8c3df722c98a5cc334b4c280310919da6a2c6fd3effd15a7aca796b3cd7f101d64d4e912ffbd1b9a2fc055fe39e23313e01cc814b8486e7ad29f3cb0409a20edc0e96088740a1bb33ba092e197521b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74c4cf14afa5504892794300ef08d37cf54782d52b6ddb930de19fe21774e0f3bc97faa429203e11f44347b90abdadaf7adf6130b290796c27b475758316aa5488c1810701a5f96faa35e3c4dc9c43044567e0b10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ddf41de4fef31297cb7014be2e9ee976c21959b2b0164041a4039f1f49008c4b5007814e6bae2b2ac37268088974ad1b8d77687b4e84c421b3ff7fd084c1ae05e6a68579f295abc693c87b2cb6450f11f637e922;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8da01fac8ff6e63e9999c799882493366789e8884fafcf2e759f9af2b76bbdd5527d738b1cbc3c38bf91fce05156947d4bee03d78148be947c8addeb3462eeaf161c30d19e970cdaa42526e08c79b5b2c200a865;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7937cf8071d89abf5a2cb00cb8bf26eec071e33a88b4e3a00a8dba2528bd820e2f9685cd44418dbfb05d8dfb13f8ece0e99995c716b72450c776c095073565b7e8857784a1bc21e017472faf2295f67ed3e4315de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9c5528f5c9ab188b4981a19710cd13ec425baa6c0bf660bd1b80ae2691de1dd00e028f71321708a4f1651b15214a1fb44c758ff5a208357d235872209f89f2e5246b3cd19eedf49ed93a6d54e42cd16aa4ba555;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d1154f1ee331f6ac9973d1b284ca65431d00f318bd4a6096acc300009765898758294f191dae03aab79cd7181d2d721be365d3aa77823ca012c60f6bea8893deb5dff7215d8b629248e9a7d86bd3eb9c2b427bb3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h745adc156063da1ef5ae423c82b4ea8b5667112de0f344f9bb8b5c1cbf23af049545e2f8bef365c28cde478549ebb733f7d28426e08ba582c5cf075bbc208055ee12c5f4a2b226b361b7776323405c23224c62304;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b851f89543acadb62225bbf0195c927517d40db1e80b1893b9a5a7291da65505500005f378a247aa920186a6ee57352eff3d2791c05f06636067e49b72fc61effb11995d79b2727a32753bc06c0fe6de2edfc156;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff57863f22427bef17553070d5784536fc743090ff777ac43f5d23277dd9deab1d16b56641154db7f7de0aa6d0d0041edadd62a89b7bd00b1881aed97275cc3d2f5e11e9b1445f67fb975f01a1ce79b02261aad68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bba8525a9866143a1d92abc57c5af78de8b98abb85a2e7811ac0b5b217032a3087ec7c234b43b80e3c022f5e33f358d13a37a4c306a9b59f56e2e52a71dd0ea37bc4e14e47c1578bda61ab6b6eacc7d0c68cf386;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hceac228d900dc22dd291755d9dc2be27e3f9b52b8fdf265221af0c77459f6e73e6d5c001400479235f3402b974eb13fd9fcf192ce59ba7d08acdab0df3b5b1d5c84ccb24dde251d7ada492b2ecb3afc2b9d901782;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e39a35c53d3b5526254d2aaf8ae0e805857beea7ff65918dc33f168513834f5799283d2c677c8d383582edff1b5b3802c9329bccef6152030c9d4d309285fc5f94a2972c3c7eeb6fbfc0cd6eeeaffdc8fa97f7f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf37e26fdc44a1ead5df01af2be7146053e24e27011d2691cc55ad5f01dfa5ea67845db9e06b1d55aa4b09702b2364277e5a11a3b8a4d376c24e305e33a01862e9f5082ffa73be8a6ded661751b76f086552e6ae29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h549a7baa4715fd2a3ebd5efe89319c4810078387845d6af9562b68099cf83a8b3ba6fa2db2c62a2fcbf37e990f6af96c1d8065d7ce4ebf42b8aff3060712009a31aa2a24b46219e685e06854196660ea8902ab357;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28d9def0afdfd5feaece1dbfba6816faf0b8516e80c4e98bf5998798018c005ff38c52d9051ecbb7d2a90e14128b40b65da3de99a48c49174321dfe431e5a60dca8ee5499aecdc8ce6c1be6571d34368caba69af6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98494b96f0623a934ce7078b02a0afbe3065abbe8e6081b5b99d614b3400dcfc1eca6805ab84b958c759ce8a890b4a7cde546abe8fcdc52eafa9b525d88cd8fd04f1154b56f10430fb2f9eafeb4bbaa3c4b4ca761;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h423b9bf176fbbb883bd37e2ac483cbb75d9c5f527a056dfc36f24be4da5f1a00e480c25340bde839981c1c13b31ae35664bb52be11d247c5b1e475b5fb0ca0ec4c76e72ab44f84823c9125a41f727b9509874f2e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc330cd6161fde9e6c32bd338a4d272718b01bfc56ca852336031568e1717cafb57f0e17214a77a6bd7415d88761c30614ffe5ade108b929b73726124b25ff072c0d5406edeca028c748e3b627f51d5d1ae466e4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe1bc5ef982d486767c4727ae00172a138b2c30d692f6501e45b1602ebf40993492cc581c59a8ddaf185176ea1cff4ba3e5481d6078baf50a912dbb0e5e8fcc80493682d4f6f89e015b14c9514c392c74e4025859;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaf37e8e0fddd09e4504298d5f0a2e0a440ad19ceb6b756368733a62370ca794ae1fb4f1437716cb311ce05b1a230bd34e85120d3752fe50c130ed5a115e02230648c7ad0833e29586669bcfa187914aa799e9628;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffa3a528400a84da55593f2c26c193cc0146d1270fe5d0c91b619704acd2301db979a3d3f4f2b07000068855f65076b36cb26b248906477912109c09cc791d862801e29ad76830fa69e1b5472ddd2dae6ca7cbc0c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47b276734cd8a519b6c1171de830bd03c2ba2f8d6c6618f7aedea7ff92badf5ab881ce7122174ed055ed8cfab762590649de38ffc0eb234692d2acb81f9e441b4e770debcf6343193b87aa30a872e1426c8622520;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf331918c80dcb92da4d82b217233fe1aed51ed7d31258927f13a21704d9bb4ce176297c0e7c3f091fbc1b148f7cc1b45ae6558db654699950cc5044cbb6e5c8b40f25a98df99f6004dbe2365c4eab90faad5ed82a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33981857c2a52d1638c952f1701053157f71794af4470b0c6c15cac185c3637e89adb44cf48494110f6e15f97cf6d7cd1fc07047142837f6d2f6ba485a9d85cf740ea7ec9662947cd7ecea85f4156d769f1acae2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3443f303780400bd9aa960d0530b2aca2789b44cd20f53ba3521e369880205a3fef289ff828b5f29d3f24815ca2f9c41bf6b0afac5d50784603848c39e15f5368b23add64c788bc939e21e0e29c068b5b68c0c2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heda6e00a9d38b640f54bdbfc1a883c56d5bdc8e98d80350fc4d5a5e00317bf330d08bafeaf20dc00e3fce72cabc2126f10d93bae7077ccf07af45e0be39371e7f63cd5cd508e2e2d8e5963267e3e3b8b269d1cca0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1d2f4fb42324c1e1e369c5bc70025690da6672fa1b6870f926459182e0754b0e5f9a76ed4074698b4f22b20eb62c9c9585394b69b2b9d8729ec964aa5d6e62e867f9951ed21867eb64f026d9f28c68a8ca4894b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba4bede0e787773208a61d29bdd2995349462038fb852f9a0ad2ba5f591cdf10cc1b1a6e4e7e41fefb3df7c19cffe887c11b79afbec44d8937d8165c2993a1ad9cc69b6ab98b30ac55525d9d8959f2ea3df13e08d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf58af39d0a3b78baaa0f3d4dc7cdb834dd68d68dad67874df0b8ca9255b0004af506b8cd986f14f4653806a6822d6ee28aecdba66a7f9354483ac6be9f646a6e236e5d97d595a95aae07f1da32060a4c1989e35c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56c39f77c8f3763bfcc11279455b59f8c7ff1425bcf89c990f9e0a90a9fe51b15f94ac5d082e2a6e9d1758edccd232ac4cc3de00dc6baa1d6cd8e822e8b9ef587bf828a2665e65e549c1289e04dde5c4a5dec8502;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7db80e173ee7f913c9fc7492757880a347eec10ead08b579a1f0ed3a6df65ff3546aaaa1adb2ec8d75023f0296e394d5743bd05d5980c640cf8ecec0806e5086508c04a104ff9ac564c6663ba96a6daf19b4dfb2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75cc266e457dc58be7b413a4945ad6a3390e0a2ba259a089b3a57fb6b6bf144adfe16b5263725c8d1297f3aaa5d6acda51cea59040b933ffe62c346624c97a48ea1c23c23ccbd8ec55324964a8cf40e6a4815264c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c4919ff7deaeb205bf281319379b3f8edfbba2eaee7b179960cfddc357333eba68ce82d3c2e286fdbe9b03db4ba7b9e9bd7d206f1b85e40909436d1f292ced44309bdb045938c1b8227c177ed5e29893e60f89ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9d2906fab79b62ca70a43844fdf7834569906ec44edaaa85a9a7615872b3c9ca443416849f7a5cb9e84bd37f49ada884425e2ddbc7f0c71fccf9258e2b319170ab7280c4e09a1ca00170664ea1427711f57bdeee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52dab016ec16d2e5e7352b09bdd98154754ded691d016cca7df1cf345265f86ce9de018e6337fc89e2aac8653255b38149c38eac666d6471415cdd64997618df9182911af824052dfce9e917bb9b9cab9c58c0ded;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3e97d9c779d5b771dfa92a47e186043b1b6220cc7567c69f62800f1da6680cc77d26afee270c475c73a3c145be38822a50eec0e3979d498d091b546a6fa50bb0902a676fdfe0079f96166464bbbbbb125075026c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef777416b468f70beb5c61734a366517601eb3c6b7654693ed3be3e15e28708283a6acdf23dc3668bda4a4c02828c0a7a451c9e4b4f59eff4d7ad1534e20a61016d73cb748742214e71d084f9762df548887d2dea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he89fd796d5f6f7a7e7accb61aa0471f6d47ae18ba2818f13dd2538d1ccf93eedd4b63eead4d51c9b6a3baa4f63a02d23093774d39cf8785ffb0f5eec3bf9bb8285cc2f8fded7fcdbaa4808294d4e0c40e2701ef6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85c6260d2b40029593501ae6ab27b3e637f9407d329f3fd6ba72fd2b6d6bd37c80ce3599463d891f7585f6bebc1131d154633f3add3009df98668871f98d32f6fb93f24e0485dde261fe50f9ba8b2bc02b8be989a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a5291590281ab9d2899ab0b8a82ca6e16de12282c84410801dc1d13fb19663d6d6f375361873865ff42f89e09f0c99c5db232ca9055480f5993147045658465aeaa70a3ff18a6eea86a4fa32c5c66e761e3bfa15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hded7e7ecb4e621a2dd771b3d8c75025b10a317640ee1eb3e7db3cc360a779ee4972b473b77de9873f1097db4a36d936d81d7bea278d3730aab555e7fc496831d6541927f0888edb8f958ae4e40d23cd954e93bf8f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ebb7a031e8dc134c7a2920992d8acce9d546432af81dcd9d3eff36eeae36e8ee30458931fb80fc6ef57e380d2cce1e62c3bd062f710e65036cdf358bcb193b09be84f37aee3f7bd1b950d610f151c9f514e15729;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd06bb08e97db829964bb5476104eef5685482177a214f0043d656c3e9ed580b0516e6add886c30a1ed749c2a50f5b1c30ef28bbabf27d057168d3aa2f7f941916814d15eb9fdb36c0ba67c688eb52beda7678aaa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h508f1f37d1244fc8cf875e64ab5a1ed8c18c8d5c55eb20b9e3c77ed3f7676b4e9bf42e5ac54ab7526675d051cf56f83261d38352b74f3205de8693903b095ed78017eb1d51cf86106a6ed5cd092c89182050206fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93c69b7a51eca620089dda92e5de662df8be34dc0de639717c1ff99630eb71c48a16cdde30e4a6a83509ce80cdf3e5996af71423fa34343469ecd30d2a9335293d05bed946e119d9fb3378fd6d8cf061f8d745ab0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d702a147d4a76bd51d6c8dafe7c63687db3c88b7b34502bf709670e3d80d755f857c9a4a3ef70d854967a0a5d24d278fe9bcc1a22e9a7d61146080aa18fd9f45e9aa4690f9902ad6a9af23966ac5778410a6c7c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1fd6a1758ebddb49f8a487c75a6671b439ff61d2d504e7f7bc127d64eff6a55da5416ba08f2fd7b6b1c37524d3d03b785c7c33b30b59a416e27e87f796bf159c8d36e61b104f21da04d22e9dc050a647bd7b66c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb33c17867cb23d60f991d3f2a34f80da14242c5529fc2fce8267125786d45daa8745846e2925e01950ac69c5cfa658fb91e380a25a82e8715a50706baf5a76ed44e292544291c5b3ad15f8c77e782210959eadf9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ee1481f21104dbfebba45631b4a62120e31bddf1a2426b0eca7ad13d4c703f336791a28546a979e007b35fcd74ba341f868627d4e806adcc0d970b87aa95c02212792d95ba620e69f32132a9912b77bab98d84c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1ccee2023d2e852f67980620243c57792a5eecdd2326e2b881055b418d91d5ff39f292d391d5490e876fbb4adcb73549e36fd8d483884ba1c4062b899ffab58a76c244c196d6b70d08036871ce3cb8283065b612;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9986ace047c87164603542f8320d34b1beda894700bd9cd155fa4fcb18838b1f25d0e31dc565a92c7468e74ee6df4e06db743280d4804a6d4c549b2abe7aac7c77b977bd07b3a6cbcb5a62dd82a170abc07a646ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd30706ad918eb1e4f56309424224a406870abed39821736339231972357367f28fe74e163c5cef91c5928bc03ef0e6132828dd6b8bd1c3a82eef9b649f3c2ba216ba04eb592b0602d72a2c1297e67f60049d13d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfa77f6721b433cf497e732ccc9d20562dbc419a103bf665d66dfda77ad65932f3606a5231274525af4dc96b1407f353215864de197e669d05359dbaf899817d02782ffe14bce5ff50f440953c2164e37776879f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d0efb1e285611bb38c8d667336cf0155f190fa3771e3a3c2f8f2854ccdb6c4f15077f6af3624254ab912a92a9a9898ddf8a592e9d9d672abb587fde97559af55722f47dbbf87625ae1a3c7027dc2d56fcbba7b00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3731a423016c69bff5fd36ea553a9345e642f89fe556d6ab6d5ef2fc52b5ada386f3a19503e06cdfa30df7310a1a05a4a8b4455bcae29f3dad207b77d09d0d7ef8c04e7ccccf952cf006fe5ca30b6e2b1cbcb0450;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h909825e3bb561c4e8ffbd674d3055bd05360938cdceb35cb49e1751c02da0b1a64ac99ccba071f29aca96a1713a0d1c12d1bc6ee00ce92e5cd56402b252d2d503658af3267a4bec0538063dacafad8e225f4e52f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf016dce670b044f6a01540bca59850b2cb285bdbcf69b3464d35813c7c2de969fa09e6a016f822d3b04c6c59cb4d6409f25709e9ed27b9cb784c0f0ec3ba7dbcfef9a0416053712b2d63f50ab51bfa22cf1a6d04b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4508a76e10af42dd93ba7b926296c15b0e2fae81df13d33cf1f681784b6d4f66410ae126963d39b8d3a03e6b0633caa0b9145e09340fcf09c927f16dedc917f88743a70056c092c5a7f55a0eca3b138a639f7c5c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdff491b926d24f454cb6ea8f556f98ee704146ae0a41ea785bd95dd96386ba3bf38c84b94b837e83ddcdaa5579180cd46174ce5dc938fdefcf9fe469de5dcc2616b661f8499a0bd561140022b9e01ca8df2abffa2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb47b7504ee6e89a524775559b67cec13317878c1260f45be8589f3eccceeeb4613c588f98e3f18ab816f1bb352bb74b61a3282f620ca30bdc5e9d76d14d0696ea3711bdc6835f9baece78572e852bb740ca01c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha49424bf578a41b983cb126c305f70cd8950cd0db9e2e618e20f5e5757571e1c4166851cf45eaab3b48c8649147b0fdb0b87d41064c79d7b04adf23b8b25594021466542aa0e2e50f999c94fcc7283d08587ec0b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcea4658c25180d11a074be7534395c050d2978f74230acd6520467755f0cb3cb8c6c48a61ff65a947d1d815713ea4cee139e9ca5c82b67bc3aa08a29e24aed9cfa3afec3b8fe35604a95bd0e99fcd0002f7ae7d51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dcfe1d2bca7dd8e350af249b09daa29ccef41af97f84fa6c152f91c1b298ce110a6e55d60531d2994c8f96f107f8297817fd1eaae011380c4339a2c6c978b8edf959f187e7ad965d70bde5935c3879110d4d5672;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h510531e7768163946df6cc54b88c7772906b47d55cb95dcbc6fd620a429d7fa289d0e9659445a6a96977b3c8de456462722c02b4f820f6b817597b7e181db3e10772cf22a92201fc10d9dff23b0e18efa4e1c8c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cfc70207421466837a4d561891c4c9bdaae02f031dae13c2549ce9d7499c99ccdae694a468d4ea65aadf0bcc7e809a960c846aa1094dec57de8aa98f267f70ce2e4afb6a5589719a353cfbbfeebd64922f2cb5ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d983cfc7fa989b44021797924b6e30488036360d7fc0c536da20d3fb4b6052e442f8a1869a3637417e134a5c24fab5841e0000d029688fa8881f9b61bf4d870653e7986b283732e3f20e1e2bd3f12971e3eeb601;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he69afe18f024e485f25a488dcfa3f1abc5f7db77136c05c8e82c5d337d074387aee3d219ad74e6bc581cea8a9ae4b73072734ff9bc1c04630ebb36cefe607317fd1b7649a60778c03437f0ff26ea90254bebd6498;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf31af75c847679a8ea05fd4dadd04155840a4431897a74c5b0725df4729d515b285e2414d76c74bd582465ba0b8c9457286df02eb0305731371642eae86d122dc3836a12f55b45857be9d84be534bda38bc18432;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5ec80004e73fb11d37eb6087facd1c052bdda55c075ed40acded68655b62d9665bcb185948ca3d9b129447a5089e9d193b1ea7f39296b6af9562dcbce77bee0ca86cf9124a714e156b2df9c268ab88540448a65e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb16967f853f5bc3e6efb9049e59b1e0bc7ce76da628318b3b43f7502678b3cc7b7986754701272edb1a35bfb294f9a2907f95f53104a101179e8814c5a9d1b2cd1a414d8dbf9488dac7a769b22a4e6c2f83549ff3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b4b82afa27b42e7d65b3c7dd4b91e5cc7582ba3abcbb821c37b1554a4c452763e4d2590591a64638bd9db5be45b517fe6f57096cfc90d5bcde61ea23ec9fe25d5725a0839fb7917a0bccfe6853884f7168bf4677;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h954d07ceda7b529274610dbb5a309138e16ad089e07f11bc846f51ae4da09242c7d8339bd86af0fc25115256db6980e76bff950d2e95be3d3b97e509949a0adf214d0f4ebaacae8c84bbcd50cf4f71c4c16ccee38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7838299a3c87abb32684cd71e3575e9e244d763bd19a1db8bea609b5bf231c196317c69484c3ae27769740e5268875bac16a0beaf979ff428e4b2206ed486a0856ede254581b3e6b96182799cf6e1b80fb22c108;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50c73b039727548d0a247bb92b3900cc4fe8e4017b460a98fa7963beb3dd62f95c089ae6929de6ad683f0c62ebe7c5d485ef8970fe5ee5ce7db25cde884f3f907d8375cb5e60ad7b2fcf83c4391a68d53c19aa636;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4b46c5d27141b5295f030db6c8c7b9dfa4335e851b228c653df3b25a19ed13be36ac83faf9ce550b9a4a379aa04473013172febac272de13b6e6bef70acd3d3df34a531921129f103264058fcb1acad808cd23c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6057fc88fa4dd8227d86a467eb51d6e1ef62465e238275b95ba6aba998602193922ca918124e46a9d88924163ca2f66dbd56dea9c75660398207afbacf3fe23dfe6ddb8059bc7343c08c4ab58dfec4f40915d64fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h328923c1bc97cdf71e17378cc0b33b47f330f5dc2e11d1ae700852184ec4cea5abb61f5f454ed46378ff9169fe6ea650bbe14050dd943ee80d5c70bc22314b9c56d98f9a0ec3331cf6abfcb0c11962a7ecea9db27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d0a785246b56160c8e2d184010bf91050f3443efd456195f98cc45c7dd9a862008f54f2ded864ae58d5fcd9374c5150f19103ead2facb067a32168624befe64f7a51774b2122d629c164272307f9af47030890d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82ac76c267403c9b2e077d74b5819e4e342a4916a081e7062d7e64d60108d89dcf496eac2314b04ab42c281afe190d67ff388aa78ba6c367796383dad38815891b02917f19f715ffbfd9075ef83a7c4107a8e45fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd6382664860003175121c045f5343ab73d5d3397fa41c8c264d87261d1e9e17b3e72c74fd27d3d8dbb9cf769f66ab0decf610ca97fcbeb408c817b9e9f3f51ed1425fab688d8463182cfe8b5a38fc2f289162a56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3a7b60cee1f2faf9a1410640750592056bfac59614a7f113200ffa0a268499b0869e4a7a0a4f6288162875eff4456ee67e496594889a65daab232dae75d12a06d9f8fa4a86ef2684e84e44b9f151e64508c3da54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2305b050a02a0e91bd730ec95a3a71d32947f2ccdc7d0acd44a0b1e25c048b633acd42d8fd81b7d63e86f49880667ab2b2909fea4d32416ba62d0811d5bb6c1bb001ffc370dc0260c26ac205a3790d2d353fbd253;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79558cd7ef6ccc4dc068ce836cf393a7f7231d481a4ea20c5b93ddff39b12720cc23dcad93a8efcd4a05de8458fe448aa4e27dc6b517e575e8acb69ca8bcc455fe7b57f606ad968e4f7beac94b8eded53a13fdd3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd03e15cfec12020f28aad0c7e5649a6b686a813b6e99348f573c7da652bbff34f3365d6e067a5058819a960f24fdb5c4f766e80cd1cd041763b9d2b6c55a299d41f7a08ef7de7f7e5352a4203c734b7b04c15c340;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e22edd92434f7a760931424bf163e63d4c0b9180f5df886ca7d0b70003a4b1f97d833c0a6805043a300358daa8e90e19971adecac13d9c9c9786c6fee8efc264c7f1afc60fafab8fc6f88c073e630fe507d4f7dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77a318b6565d63d64d4df55f0d45da5f20c684582bf9c0c53bebe6c66eb1498ba14f1024f6d95d76ff1c45ecea4cb58ba5dd7f8f6e6c677841fdcf6cc0c64cef3a820a5ef0c9dd0e02e7ed3115f97c89d559966b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cb52c9864c3d70bcacb71c2b5d987ea4beeb314e27bb097d64ea2465cdd16fa3c89ea11e6998241da8492729488d9d02d937221a066841c512119b6db036184dffc1f1867b986aa912dba8014ebad45e389c88a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5afdc49eb8d110736c09b11d6563e85e78ff87db4a8cdc400c856a940001425bba6084543bcb60f22269766a62a8de3fa72ec96c8534ec0da7a00d6fb40fbcebc12c95d51c392b7b5e2c5afe5781293b6b64d4b6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h811b5d1e23629f4a6852d9c4247bd85057ce0899cc8aefab77c3d3f61d83a0413c8d22f5b533710aad35f211fed3993d52cad3a796ad70b46d3a7b202a99527dc4619ca2c4d4ff3418e9ca263d0c8bb62f94a375b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c13c41583f42ca4f5998f71d73de6744b02aafb46da802075c8d043ed7bd9b0601b35338a61f4a3ea7d823bfc74951cee00fd5f0575eb50b72995b2c8e384f26f0ca59ca1239f96518eded62b28d84323ce895e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35da2be9c440096fc1cf524c945efa7510e2a05b1112aca028e858253b38b5c64124de44c89eb29ea1ec3ef3cd07f29b77d762cedd40ce364b5038d4964a405dfe52e6418dea6784980dd1f697a2a6dec6b2f6b9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1388312f695d85e8e68631bdb7747490fe6fbeefbe20006880b50f133b3a04b741e07b7a37f461741ae94dc0e1f597d526510fd68fed06bcd0c0687c72d37444e824612eb2cfe846e3e1673de93a8af66fec0bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf08982e344b264fce468eee453efcc82efb3707f4b55c7f7e5f3df8db471461763e48c74cf0c78327759d4f21decd85970920736b5b68b1cb4473923ec64cc8f59fd311c9d83c4ea4feea2d4a98aa4823c075150c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c7d10aaeef3f533b9d4fd6a82541d7d44a47d607713f9a16a6834294f34f150c95bf8b7574e742486af718ca5af906a6307ef37422d20b7a6d1b32d0437129d3dd087f3ac0f149ddfe4504206e5013e5aff73dc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ea56ab8e9f4ef760aaf347b63c4476cda0e5602258102865376d5555537c53787d4db7b0693e38a0e779e057a8028f4c371df23daf9bc2bae97867f21fd5062b4b4b2530525f974cb8235e5253e25a9305dc3a7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35c6f5096a501272afdfe0c69895949fe38b46f0aab4179a465728ea5228d1a41308b5914cb2137783a09dbdcdca1dc9b5f69e87dabb6ea7bbce56390549e196e6ca018e5c9cc9539a16bd640c18ad74c1338db6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f367f6572267d8015ec3fa269490f671d6fb11bda182e4be246d5551c0249140138d52393724fcddd2cc1a82c034f6117fef53b906e018ffae9e07d9d5f54be46db6f859bb9a3e38cb01bc35c6dcc7a70e555b1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92a2d75ae70438ff39aeda9b28a694acf9ac4b96d264d188e40c14bf514486616a1e0aa07f69c00e2cae893ba8ac20e356514d711ee682bde79c33f8827f791b41d950aa3db45ba41890a770a69aee54a6453dee0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cd38ab290b2bb0aebb74c7c4e102d66b6a18fc0a54f887b979d9d6053e7515ddc6fb458737079db00a7ba0b4e1f93338f081a9aacebd7619b151aa4fc147771f49adaaa1088117180f64c08c6774180d49a5cd0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bf11fe1e8f05d8faaa1c2d7dc9b68416b24dadc616763edcf451e4138066df3cd9524d1e213922a378859a34954a35443581070ee8c9c5c52915df4b9f845d107a4ced8c69ffb0cabeccd8b3176de9dbb3d2784c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fb710b4537864f2e0cec445fedab575e116f29db3a3759e47a47e13e8d30dd372bb31f2b2f02566564790dc7ef1ee2d697e478de0de957d83880f1808aa29e6119ed7be96eebe4dca95272288a63d9a84c6f7441;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb8be51a378e9557005c89fea659af3c206e697ed68b53db6a02f2faf3272ec62aef8af51680bd459a2a6bc42c678764aaf02699f951644ec61b99ff835cc687eeb141bc93125b6bc7f0a894c9ea21fa51df776ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he99f880abd8898788560429e9973ff39d99166f3849682bb1339ad7f3c9f2bf47c5ae830a21a6c605a28598912542fc36714b8a16b54aabe4bab6debe1909bae2cd5f1ca6b4abf6a945e47817948e8e77665eb6c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac55fef32928798ad0de41a2ce60c9ea4a07a7354306a75f215d83be0e8c208a9d2192e01018868e9db0e8f6137e84c97ca716a8f672c705d0aa0b1157d01e567938d4a257f0c3db4fde46e0ebde3329efb99a000;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ff31ca5fc07d3b2f7e0143edd888cc8e46e3960c3bb139b73b93fbdbada1696873b981a658981bb3aad3a6ae8d5e9362df59b498ee9db2b779235154d7dc46c5c3972f727d97d64403290b52a89defd888f9ec63;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8708aef942fbf17acafe245c277a818b3330f14eb4f3b99e1dbbc2f1e01da4280dc7de5365d8894d16e46dd5628e08ad7ad42db87c079fcad3deec4a566cff0af2c702db0e543627d4ad0bf0d2ddd8ef71a605119;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca3bbb7af387c375dffedd0cbf92f8cfa23c8de2cfef460a3d8ba6c6f90e89ec137fb0235edcfb1b8325b16a7e8bbbcb13db564c0fe090b0f0918c0e1b39a44a20be025252ec00e8b1c53822f3ae7f91e44998136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8da274030cf5b926ddbf1eac7b9a2317ae5a7050a4a11258100d2e29bfda3eafa8a93f43a0c6d08f4bd643db7b39f3d8f77d2e2b8ae3ec5cd766f981c83aaabb71cdc564b6b840e64cfed0370b7b26b57fc8e96b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb28d19750518daf6e8129e7efbc301721c242b5472c42f143e972fe8e22ac538507f9c73dffdd9de6877a5666003dee486bc0f30e1384783d82cc5877a3f8df4201236b96004ba5b63ed60a12138680c7e9e355f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha42567a1ad192c06cce46fd61929902e181c44a0c1970908173fa2ec91cd88e5ab8ba3504515109cd9c794a2cacf9da8a017ad8a0f9c885da5bc19e4dffbf6f1b19a5651d48b23af16b0e9aaa9b8ce33b6f424562;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc09e73b6b3721826640fc19555c5a2a6b1be2110d8992d6cad88e76dd3c4e8a883c09304303021b0f177b30320bd8ad91f90881e5cdaef48eea91c6f73a2fea39f4cbd9295449d511b8370da95675798bc6b27969;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha19e0b203984ff1ade8d60e56182dec7627437b3c0e2e032786be3476cf6c36164142923563bcc1daa4c842e71a7b4af4e12fbed5ce82f8d71ab0777213a34016e8bb21d715105cf4dd44227f8d5bd48cf380d6c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h776d4a3fa7b4f4d9c5358482c2ff8ffe0252ac766d392886175a4e0756d6eff0713730cca281d3bba308a084b79d357100fbfd235c2ea282646033c118b822d7af1f0a84bbf213d308e123ba63e6aab33ba527750;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1292209c5a2cad773712424d9b88a65eea0701734a5940e9bf959ce32563af12ac51a44dc5af40be7f95e8016610eca607dba20f668ccf876fa9366b01c863932962ace9d79ea15fbac1e7ad6c0be3ffb69c02f68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he25e625c206a99c2fe7f4de4d9e711bb1136c684232e39d0d7f2fc420118c62f1694cf1b508df7f889a617c1adf0db2d642113508a0af29f8d7fae7f6b030d5e07c198e125ad10b3946fac850f4c00eb31fa6d501;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd987f923c22c2a1d6698c6bc51f1eca3713af64a7965f15abcb7b162ce4fe1c4f6723ab381827984acdc6c19384b0c68b4a56402a670382c83531832706816dc598b3441b2555060d0f6bcdcb40167198869eb2a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb122b7aa86472476addababec656d7c23833f5666a37b9904de4c363946da90b9c002c33d2eab6bd406efe44e6be4f35536f954c9274371feab4895ef887845a6d6e3166f941e57585875606bc627618ce214ac2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3707fbacfb49e239f8d592388cf4e94fa5865bba4a9cbed39bd03cf3da8aea054ae6e64980116028e09434d0bfc27046e5003d2f394c9a4079df8010f7be2f642d52c2a1fe44348a3ba4cc5a5673dcdfab0053d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe1ab722832e7c15b98a124b462d21075db9325141b89fbb739834c2b2ee74e72ae07b4799f7dca11921d22927380e13a2ef880542bd06ac085b03c3d9dcc92988a10191e56067a84cbed4beae2c96549786dd6b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8e00c3943bc61f4e81ebab108ef6d295be51d58f122553e5d9365df25493a67a63a3e9c498bbc930a74355712dbaf7bd283254bc5c9f86f412da1fb414ca2e16aa0a913a1db23f8f85c82f7be8d832d9db4ed781;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef43d4574f644f66f31f3f2cf5fc3d1c72301fb79ea6c909512b8f866a6b9d198bbf2055986ec822bc408aa73e777bca21a5da82e387e37649d0ad68b9d01e40018fc0099ec6f523705cdfac6d6d39626c57d3d2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h918a644436de83751c2feccdafd58037473ba205ebe81180aeb6ed830a1bffe115caa5a36b2347ede5b6c7e1e0fbbd46cd8cabd68b19930da6a90db16c45096c3e6e034fc0d0e4d0abd0674bbba52d5fc745ddc80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38ef11295f183df01d5c23991c8199f85ba328ff676d603b2dc1d067c8dd486e75406da38e75ec3f9b76dc2d6a711934628ba0d4dbe9dcf63bd36a93ef980b015a38a9ec4ee0df92f5b500893cf308ef53d814f88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2b8000811c1a42386698775a635f5addcb35f2db7eee7c812c9ae3d4bc01346ebe6f62c8607e3800704d9a25bed2ba29d46efa90eee6f53cf7ce534730edc48cf6e36d74819a0452d7fe8d417c412a5c65f7e480;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9076c3e164f13052df67041573f675bcad318b6f502cdb7f64cde37afde40e8524976070c4f9d5d289984c69e059cc3f07f0cab066c8f1bd1b9288cd326079a9f9c729f6b6ab6791b3494287f33d0dde7139c0a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d6b0a8b6fff11c293d349ac412b87c4a5e528eadae7e062f9f6128cdfd0ac9b6c777d33d71104656dc70525a40797cf08c468d08cf6086c64241d0ceeb7d4ac30270e2bba002ad270a965d7f07d7f474d5845325;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h153f0df341caada6a7aba8671fe06ad5da5ca6b2a7a2711651df0fb5d43771871ccb5d4c91f2fe635c56fab757aa6e86e250f318e2e851ca6d53ab3d90e9d6f6675859430557c47ad23220c6b0285725c0e15299f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62f1edf6e0568a0045df4d65b175e43824e26fa9ca37d469691fbd65b1b16c6a048b127f03d91258f7f755e8879221d5280adcad67d15c23bb66b11ace0764ef01e99518983c452a5c8da79be4cc8f2b541a3aca5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff5356403d68c61606c4f11b8bf2105aba1e1e0e7b928ab1e91b825fd3f16e76dacde5d5a8945eb9334eac06577f94465b8e4fe41ed0453d7aa89a28f60cc4c2bc59c45a5dd9dc6ce37d0d67747a8d59bea16194;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha63172e4e3303ba9cd25f33affab44c06bd50ec4c338343062224e7f46233ab8737a03ef9196f0f10a84a225562acee46fb7e3c17a81f096f66c29c9b04966c8cd46200ea8b32cb074ea5115ce95ba4d0a2ed0c0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5beba3b0aa6c3e2f81fe8e172b46b372de65ee3908d9b7c1a39d6cf9baca7211e67225752da70d3baf611f43cb338c9892dfe3679a5cffec39f6620af7934456fee15a7b61f9ace3dc321c85dd464c9dfdcd18b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88620695a9fdc5f3136ad940717b931ffcc5922dc76539aac85d3d8e001d06693e226625fcad26965aa6da8ad4668d6af776a903509dfe94d439baa3a72b1437b877d48f961ae2afeea629d53173114ea6e624be0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12bc6f59c0cabd7d9a0b78b7607066257c9d217e3cf8981a18ab018dd233b5927adb7663f9694174a1d3338484de78cabbc10aea3f1fcb3c02afce1cd1df755abb4c0d56a0970cbb3c5e632ab2340f6e4493260f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdadfe6e1681b5c63241051fc9744fcc7a3db315e21b364373b85aac9890014aa152b50f523902ef454c0c6714e62a52eb5acc1354ea1e17ae496824d897515c7e98cbd859e3462982ba3c1bbb68ec4c25d9656b49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h964c77ddb21c8c2e93610a4f5c49ea354241a52103d986e0ceeea0f93cf308b82f13ba25dea9cd9ca379378d919064118c5b80b32361a57f3a820cc39bf2616a03762d96a3c83e8602b870c257ef15174faf49e88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bfd5a73ddc932c07ce47293d6629d3961dec97c065f9f5cf21181a402cc2b7d79839c7f1eabe3a836f599b815bc1b1786bb4b1728f8a7a90c33325b89ece3d1a8751d5a98ea5011a7c0fbf5011144cf28449322f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde29addd45e27df76e6eabd22e7038ee48495a184152299587c3ae204a5166f3d0a33b15d5a611bfd2e65de21acbad7b094c8beb3654d6cd29dd5d5f9d9bcb566337c5d85339fca88a47016773f04cc02f1fd1b95;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h720230aed76cbf1548401f8f45bb80f33490663d8e203f4f290ae2d7c62b198d75c656402c2b0eb094c8faef1abf3a14ae65f5458b86f16eb6e3218cb935f1d6a2c6a305a05af2e0e6c74c89df1b7d91b1d597379;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12895cb5e055fe200ea7db1e2c46dd03f3b7eb55512cfac62f56c271faa4a51e5664f6fa0525ab648b07d34a9dbf915477eccfa7a5807503e5b2ed7953003c2344da0e8fd1302da3e7aea3af01eaedcb2a616171f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he689fc7e125d7f5b198a97383d328bddea67309aeafafa91424771a8b565bb3e56a1914c29953efd228dc1220af8fda3cdf47d452bff6ac25cc6a17cf97b80dd486fa12405357fc7e6f723bed21b339178cb02ffe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6031a4e37916e0c8f94550ed8081e52184484087055333e3d7ae1e79383b31fcd45dcfb7cf919bd56258ef947deea6003436a7ba6cf18e3b14ce0bb0886a6e43d7d4f343a422aec9b5f4b0860832f8fd931631d61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf85860ef0f23dfc89cb09846cbdee296e18eece84a911db63177f518e17760d0ec1514ef08e76820f22945fb8b33f0078f41162b5d16c1b49c97f64f13ac10b1c4332d9a6dfb093ef9e2786daa17b456906c24533;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac164e46907f17fdcd4ddc4e36711ee508cc9531f3f9b1907a87e1202be219e361180e18d640903502476337e118ddd753a5238f0e4d012ac7e501965ba04c2d50fda71a36d51dca36273ecd44922472a09759f0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2b7c13e39bc39c752c22b070da6541a93e2a84075399278b894199567a3af1159952f0084e341ae1f08f9e0cc7c48f89c55defa5c9ed370f069b5b5d3c90d10a2ad0bc21c78c7ca09b76f419a84a287d6ea37ddd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b2c61f5fa188b36eed4e09314d23187e4680400bad91da5859cce1ab6b8c315394db8ae2dbb90ef75f0f4949c32322fc0583b3a03b055118cdcf3409ca64d5d4bc0d660c31632db5951f274179d7b5bf982cebc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5467e226004cb5b466a40e4825382fea6ab36243965645e45d4540d63a1ab48dfac51813417637341513bd6674d200727a2d3a5b0a9f277654d1229c0287f84435c16d438cd58947d511fed7f2162f16c539bc161;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9692cb1717fd492c9fcbffe49b202a68c631bcc0231d6a54f130fb819d9e09106af265816af3aea57c85d4d9d14945af7f99360c4a454a30949142906d3537751b3daada1eda9531572b9e2176d6e250646c60716;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71a6feb64aa93b767e79a930676eaf00a59cff876e9a8b6a508e38021a141c45d4f1bdd676d42c014da90ec0a76e7d2ff35b43484158efa971af3c6301321695883685c311b21405a455b75b68c1e4ce52b1c876c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce15e4f22a239151bb5ccf9a02e54ab2d0b5c3e0adf1134514b6f07d53438dde40291ba7ee3adc8a7e975d4be2d9bbe8931874c230aec19940f7fb59cbb1ba002ebd1577201651649f79e5a8780e3fcd2ec7ab7e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ebfc48187e008d0a29937624a6a7d507c62d2194df131f22c8b4e67add4b494eda0bdf1399185a380a06d9f232f8e1493a5486c86e20b9dbe9154f704ff780349b71fdd4d61ca607cb49e552a1671e967c054459;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffcafeeac48d029614507a07b54c67a0504a84fc6eb3e3c6372b16698183f0e3e2cdf95ce46bd7c5b7ca7128901a45675a14f67ce610c03ea46227a21ec0ec6e86eb5d72548d1c2dafd15a6d4cd21d8aae358c22e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39ba29dc8a9eba896d2be437e8a73fc60167b830f8236cb62bc023f4e9b632e826b2665aef7c6e359817b5e79b30353d60610eb87bc65d33f3703d57f91b6084acc57b89685c24efceafa1f73c79113d018575652;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c25d4e2d036e15bc2f5fb2e046f7bbf50345064705ded19d18840403aa0761289d42d42993c056e11fdfa9d80bdb4270c12f33e668ae73ccd42337b5d8da452a02c3800631d9226ad62ffe94bfb4f89081c3b6b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7d1c4bb8199f45558b4b25c4d6a8b80dfdc4042a46c61409ffa12318878c16a55a72cce3dcd8787c8a20942de7924817269763a721a1967fa18a1057feaae5fbe76885f080000eeb12f275d9299b496d0b3d96b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h535e1b6dbc3d3393925242ffceac8e60e96532d11115b2e99487781de5d91f0144d490f197ed01d710b216a34b22e6b4be4c952a6e849af1161cc1b209fedbc93621e19d875fb2369cc97facc79fc2bbc15c8cf1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dc731026d5820f36fb0d4b07a40bb6f34dc5144bf2a51455cb9aa97b7029f251615244139a7373a7bfd663ad875270a4d70daf69075769fe464a17bdef9879f867dc239ad0844497cac0b966fd461171b1eee7d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1112a01fd29e74741d17ba2d792ab090fd0732057e6cfb41b75be45754d5b033d47090c2d39d0243fd37b6a7b35a5a018670cca2bd5479032d83d3b3e95fabc7a54a6dc9f5ecd07c6c60949bc01084477541eff6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5286705dcf99b3ba59e8ad0b6fd51bb6b953b955b147a3f1b4e7085eb611022b21cb0df4302c3ebdecaa78b307073e149f587d8057f3b28cfb70bcd49204424cf0e5141d00b805c1cbfb7736c1d4d9f5b5b7d483;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89d0dadade05eace5d76dd61439684fc3cab47e2115ff71e11b8039aef76f0a22b6976dbe350ea4f11e70cffc68960da422e474d35e0a88a6177a650133901baf7e1ff58168f2029d7797a25fe468f634d8afd4ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92d32d2a5787697bdb2cda7882b7c2647c8705abdbddd10e3c5d3cb2dc8c7be33ca4ed8c2b667647c95be8082925a6c8b995de0d00068bc8b5e2476796523d2dd1a1d0421b8c88e7f4c2ae443399510a7e24a6e00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd566bfce587f8498d39baca2c72e0a1a7c8028216ba5a26d094aee458ddb8d10cea80ab65a82a2c6d9bf9aa6b3be25129250dfa029fc470bb99eaeabf036a68db81044bebf8f3479e9cffc21612272771c687dcd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8d0fb3661f969666a56dd2040098b39d756071a26e86508c0cda4d714ae59ea0a066b0e849a164fdd8c4fe980c00937206f73e79676ead7e72a0f336e7c8b1bc2c3ac60e9bbc9e798efb5402e5857e09ea5cfe8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1513f19dd6a55c00462507b38f796a4be52b5df6a633f48ad2f6d3c3fda0d001b58b7e6451fd0930e023b418402e7396de63213f69aa345e258c4b389b9aa391c7c3c134e835c6731e1e2f9f964b0a2c7387051d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41bd6a0eb200dc607ce477d0afe423f778b7c28f8e2f497b63281e0e32198ed889a65c3419acc052c3c9e04807cddf86ad653df30f1b054a0f88b52d8ca2280f5aba7d7cbc98f0134df0c07b4bf9de05c5ef6c6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3c670aadfe891f129d8fc2a5c92c84a6d9eef5d23a0ea15e79b69b0e0be4ff2aeb7835322d3ae935f55eb572217cf75fb3ecfbcc53f97240f3b8a7396287531b148bbdeb2cbcf4a555ecbb38f687977e5aca201f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdff65e6a4db10b6a6e575e7123f6c98e025cca343e574f2005ac468e5316dd14328626cfeb4dfb3edc292996c52b0ec67cc7c6cd5675faa2dcd7f938d6e79182ef9027dfcc94bb382330c1a2262a061903f744349;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bc91fe6316198c2d1c2db86b51f9f5aca31991ff2998a0055782cd2fa3e5e7feee49621e307f3eabe5e216127fb53b5b860094fa4f070f23a2416d037df288847155638e15736909db3fd1a815df3c967f4db7eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h643c0eb7c102a685bd549828d7b2b8423c208ba03dab7685d8b06e198caa0f1cf594354258c297966cd7d1dec59dc74e1afcf4bd58f107007027717dfd2b4bcc45a0164dd76f85e7095023ac054437a32043959b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde7fe98299bb443ef83b6acb4666a5f29da98570e237ac59c95ed350f6f0fb2ae017d513c4f70526e912e795597ce5b24192420d84c67a4baa306ae1193a4578b90712d2d3ddbfe7445aa58f9bdc9281b2facb689;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd49efd5ad0e7cfd2d99a877a1ad0841c52f8aef21c6b71785ebcfbe856da9223ac5979597764209ed46530d0e000aaf55263cc6f72d26290f9105f030c59a7fd4e11403b4ce90501b9da4a4ab4d0d45f64602bd4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d518672deb195e86a0ec0f2bf4e13c63695463fc8630f33897ade914fa0ad03c9253fa9a37ce151c73098cca22a2cf16918e11d4e6938734f0306ed37346510f491b0fbff713466f8b6cf08fc99c52e149f81652;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69d1f39b22d9fa72b1e225f0f16ef9e5f8512787e74a0a73795a9df0cff83b5e50ce824052768bb59d4fb747cc7a4c22a4289768ad7595453223b845f0bdd925277c3e8e69638de5296d8054c576c537030482768;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81a987954c93169bec25af28e9becaf838159ae18e5114883125cb2046849b55946ac8bd17fc169702308d1ed5efb940fb9c1cd8200e9e474831651af160fd6aa0a815f20c74df137ea70eb5649fda21bc9195065;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b60cd1d6989fe7c4f5dce9cb23bd8362a9bd13f92beba742a66fc959aaf6177d7bba59738865d493f9aae95579181ecae57f9579d50af973fefc291a9d9cbf3d96c5b19d6482eaf70f803dc4713fbb51aecb2e43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc32ccbcbfc28c1e26a0a2a05f16b671ea81604aa81cee8355ff57e5c2ec433dfabc8eac6e21deaea4de24a3d47258fe1b31faaa8e7d416347d64052379c76ffb5b7b37b05e922a65c9557eaf2f0f095872dec3960;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaea04754ba3edc8ea82ea1f1f3c925fea7ac1b148d64ee19d4137c051b2160b37a76d33418717a8295a48ad60d51d2152aa3c078bb18d86af50862755a8f7690a10dba99248e8aa9bfe91328c5760afd1351a7db;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30da1b15d582228e2f8c40d702cd2eae24bc47a1d3a52699222bb0b569b95ce7585cdb046f09f3458ffb4fd095e6c8375385e63da28c5a871f347fd4a96bff0a541e5b63475b92bb8a6a02d8ccddb491ff0b9aa15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa4a9e5ddfca6f873b75f7fed8477aa4658c47e9c4b685226ec6b68cb126bbf44cf8fbe0842b61be0e8bf0d4db94f01b1b4afb35e24537c188947e9db72fdf73338b0f0543b2199cd7a46bb21866435ba06540cad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64ff4ef7f38f8923f0089aeba69b4fb7eb6cc15d1ffc1e69f2a71d4e23068aca5de2e1d3f1129be17caa08561706c4b7bb8e2e5b9c11310143f81b3efc47aae7ebaba78468701df77fd166826160860c641d7f3d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b19c98d9cd6b284d845b241f60d38ffddfb93ff95aec1d66dd62a6f1e25b5f847129691718c05d7a98389e5dbe55bc72236646810f5396e47a624537d336f45e5b99e94d99173d394aacd4cccd1044df3ea99e0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff8dabe55e5e82403e9d2593cc981dc797f855022d6496bdecf6ac95eda9cc5596639f0a78f643d47ba7f8174e0446424437bc465c9fdccd9c90e3abd50372b24c7e1e5ab36310e43597d11ca4d30e9f69612b3fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h797961deaf9c9274a9613e1309c3c9a8b32787bdf18825e90655c5f651fb07c71c0ca4a2de46cbd816e78ace20277f5cbb68902d8484d0a912ad37fb747d5f052cf9a5ecc5599bd4891180336e9de2ada89abcf87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff18eb55e54ac7fa6af283c65426ae6eb1d4173a62ca170e1405b55604b2e19973aa4ee94d70ec4ff48eb8a588e96b83840d046216c458c2e7f105c70b0b75394cf9e6d4f19053a675babb8e9f60722b53b18d703;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b624e5539e76fe01debd8578312ddb2d472c41cf7c812425ec674d9be9acd640e3308592b09eccd2c244021a450d6073de287d878691aff6fd3fd68394f63112fc7d9c8edb4bacac010a4818836311cb8af7a826;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18df51eb0feec985ac8e47fe42ad06811f894e601019847a50fea35c9a6926d41d6d140e6d7b3e0a0f07af763e8df32e08a97a600bf656ab33582d7276e4871209946eb5bc8fd43ec469d82eee8ad1e3957f95116;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdedf78d63cf521639b487ebb748902c62a59d37c80d3fc991238bb1e92386e95d2d4281872fe1ecbce1fd957cdc48ceb757b2c4494adf096fc2a2bc6c9c0a40dde8a0ba7757d22fe4d1e0770b3758efa0ca08e2d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfec98a942758ed4209d8abf10ad5903825340b3388fa88ebc0bee66dadc1b4468d5a0b6bd28dfc830ee5f7b5754abf5702a20913f46a40e468de3aab6b1620ba5529b2d3e57e5ce935e8b43fe8995fbf4d154840d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1851cd8dd0b41b46ceefb5be848ea26bdda85e13f79b9625955f9afd2cb48c7e58930bd094183390cde6a03f0c0dad019711e0baaf295db90cd7cfc5146368337f89b35fa0fdfc5b1213788153375c81e49cc4e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72a6036fb14e31dbcc70668cb4800adb0e0623adf71bc31c43d4c95680cd79bbd6b51a4fe8cb662da4d7df283d053775cdd93564ac9488a5de2d5285b3d1a809bac132f4e17e86235f82367815a1f36f67b5ee18e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4efdf1f6a4a5ec438290b10d74b76973659df22f9d92033e1157b088085ac14efc1187b916f0610efcfc2a7f5b1343b38e5f6c37a88995c1133f25d053a6046ec7df386cc10e09eb60a7bc00aacd60e093d40a17;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf78a86f0e5338290ee0abe1c44a70a4be1067b76d46e54e540fcfda0d66799ab9df75a08c37fc37f2a8f784d0600a990486ae5e5935e676ffd28edfd342a655a7457f4af0b09ed228c0194992d81694f075b067f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2723c82f4d2ac44e2b93ee3daa40cffcf731e1faa02b5363a0e67781bc25cd5b5640b5290ca085c6ec27d48cd3abc23b58bdd9a1c02281333008434b97b6edbfbb5d8d8e8b7fa0e63cf36eb08c9330120520c11db;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h665ae65a25c316a59f71b3f2c14920e3f3b74e546107149cb48e6557432f653304d97280700231cb1cc83540116ae14b4f11b20291e58ed153627a56e4c7055d5539aa3afe39b086f88cb6d83a40fa3951d834abe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h141521fd1e93b1fe05eb3e9549fb6bf0f25bc01943efaef400924f012996c156c49fc68e453e37e7896bdd619abc7d0ccaa2a0164bfb64a794d9c2bb226f93a01cf624bfb0da90f6666588ff1d7772635f50f5551;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc802651157b48476efb6b0422d3243b747b0a0283e760d603a2dcbc05ed925c6cea11b7c41f949bd04c5ccdd71721587f4486e6179eb33a71cbaa62319453b297b28ffa69d7fc21beb13260089ae406a1c72a5789;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3c1481efc4e07a31b8728c3596c5d7db2f1879ca6d269034f18f4b33c165a2aa60b0e0f43cd6afa97299bf020fb3094f4f99dbd58e4d61c08a9ef7948211220601358efffac9b6afce73a53d88a0122ba7b4ce0c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d5225bd76c246e32a09a2a59c472f7ab85420e454dc242a43642cbfba896d17bb18250bde25f9a50993e1739ca2fd91a221c968b8905765c952cb15d13fdb2cb4ab3979380f32ee24de896a191872b335387ebe6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h750f612fd24951663a0c627a253606e84285156d5e2cb490a35b1d0b533bc7e0ccbd4512ea11a74bd0ac8be67623e96da7f0daae5fbb0ac9cdbd5f1be8ae5fd37e84f3fe5338b875806ba4a321ca9a782127d209d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f177270eea15428024dbd7d36fbef198af9444e720137dfe3dc15080b3235af7b05ab44809481b2c666e7bce03c4073ce5863d7c05fdb0d50d5624cb67d8410c0cc2dfbf405e8beeabe1dba24ca227a788104504;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb987b95ed3fdf4048ff99dcf4edf269b2b2becfea20a4918798fb5a1ce6df844715137f43ddb222d8c2e99d794101c9c68d6233cdba7ede8b28ff1b7ca7cccfcabc1fea8900c1a43bed157ce6cd96a632633bd3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ef470818ace4074faf09feeea92578371f18d9c5ed5484cb794b66eaa9e6c90dbc05ff1a4f09365bf2942b73095cdaf576c9ab1228fe8893db2eb31f65d7ce267fca344d6b03e004c7f5496454ad8629fbc9db64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdaa34835248e0ce52ff1384864a39c21ff39918a7ed9e94ffbadad93ece86eb807647a616c2eafd2642f36646e4643675df9d040fc3e6ec262f2a63ec5a35431d6bbde6a8383311d59ee0b267e786355429a919d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ec605b374bcdc25a9f7367c99ad019175e3310dd5087a441a82b19caf5fbc696eadc93ac4a1249007dc7f22860d7fc1d445f2dfc930e9d377215c2527a64c8ad471234df0d68eaddcf1a7a496958ef207fee05f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21eb74effe99792479ac3a36ccea458d55dcc6bdb3d3969efe537946efa5690b0efe186e36924a8d87cb76c77cb1a2f1a5efadaa2aa1a77cb3164005e6de0ea72b0347c6c16e25a6ccac3e3ce241dd3431569f2a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c2280b8e3bf2653cc40ed28fc271116a7d5bffa6eba74a2028482e5e11bda217c43cb23ba4513c7debe6b3006e35ed4838a09228a6bc7bfbc20d4d569b2f66ffef25ca92a99e098849bdcf3e30997f9a75633c4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74a11e60fd73ce607079c7a698cb2156d0611a823cc9b4839129c21bec38fcfcc714a316b50c02ce963191a3f86cfb5b4cab6b567ab5b5d1884872581175980263f91c1c8b31373cccc3cd74b59dd893e499e17b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h739a7619b9035296fd174fcc659782c29ee093df727da57c03b55a29f78c8e11a6f5cd8fc0fed7ca016589d7084569f5be0667612c511d0fd7ba094adc41405b9dbeea09a4b999f1cc9fc16117d6e06856d8a3a16;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14bbdc891d061b08ee7e8cb62e4330b44efc1233bff149eae60fbc7f03f1adfa2ad66db0524d898cfa8aa27b12396ab68671e32774daf8150d80097162cf5d43e8878ad605906e2eb089cac1388e6c79c56116d40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8073fa5736178191561c5a13c9b659bdf4837733afaaa6b3cd384890aaa7759b6b938b04b915eb852da3922af37fd7fd5c83c2f465d9725da6d8120cdbb5393d9e64a1a533144a659dad38e6aaeb9be6b589063c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4e02da9002c008e391420e38ac7d4b88d6e937c4fa463d549a69cdefb8536b70dad9933391f5a47944c3360f211f7337ee036c5211ee857d6a42f288ff4b4c6e064ab457a81011372af52fc2f39bda1120acd53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8917907010cc722ade7167efa3fe0db8adf51d1aa608443ed7c3953c986b43087fe7d95e55f69635cda24ab51eb3e6f0d7f0effba383ce4c7eac8a77fc6c69629d7e6fc39311a8bd8c12fb6535d9eb60659ba6762;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba69cc658cc17d50eba89cc81d8b5780088044c690b1093847628ba4bdefecf2ac6bd956c305f5b37a276af7faa668ddff60b701e6ad300e2575c38d77ab0021159d82221c3b44e681f70109999050f22df245d4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8de1c5241d32208dc5877929d1fab574a4057341d57ee65eb0241776ba0d2bf3e1832a2803fd5be1ad007ecb693ea617604f085649fcf047bb8f4c6c8de8dc46ca219f6a54d046bfd4793816c21e2d4e3265e08c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0e435b241531d45f6d9f95feba31cc176936d1f6ed37c87f0ade2944369c9700391bfb23619a5171b4b7f9628caef67050c6220c85979ff7c24d6d68e740a4def8dd62941dd9fa38c4c084e2607ebd689a760a08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41fbbbddf4b6cd7a536ff243110ab74dff404132d34cccec411bab14058b6796a65d953a26c6b17e3f9533669b124ca27293482475ccd144bd6f588d9b03ed7ac082623e8a4424cd812055d48daf03b6f00237768;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h675ec1205a107a6ce2894891f2f7d8412d45e89962966435f47c583de2949021831001c4445b7885f6290d7c2fd74e8ce8e4046002ac3419b0a67c6c71a6300a708712a58c5eac1ab933a4d4bd00a1161b628cd56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88af7004c3485bc393de46bf4719b06c5366519a3bb8425c7828da4b0ec233f319ad1dc9ade42737e71b4d950dcd0b5e653ee88fb4e7f084e886b711a067f563835bf358787f40cfbf84bc8caab649fa115895222;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84a70580135d25a834dcfc75fc96467940bbf9497e8d4e3bf8e37160c598cad3183dc508cdee5ddc3b6ab86a40afb1d0181ec926f3a284312f3dd4ce6e1593048331c2f7d55b2cca606708d36056cad5cc7ab7a0e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11b692930e9e9966a4306bba17561cd016e688a23844f62d5f32fc38615678b48dcfa5ee44c7356aa0569b72b99695a0fa57124acf1453b8422bc97e65b2808467e3e225c4e994f807b508ea84160def0697e35c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5b409898c35053251fd720ddecd756c3d92bd02a288c187eff885b3166a752143addd830baa319a0342657f13b5cf85153f3cd66e6df158ec150a017f78034cd934ec02fc92cc7a6c24c96377fa94803f744bb3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdd8229158d40d1e3ad94e669237797a45c6ee1f3200df9d1407923f25098bc49feb99e05367536437a9efcf3a2fbfe249b85c5e96800e002f0d030380c330c37a5792760b520a4b1b9081a8c2c30ab799a389909;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26fc66e0b81d0d9edc6b2d1b884159a56a45116807d4b9744b4d3b026cd9b5a68526690be214261a1836f2b6bbf41bf3ab45d14f480a760aa6171c6805a806b802349841a3bde91fa908e46779d1233c920d5f69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4fa15cef66bf7cd7b551a11a866f49d34ee9f497b5d3a6797b295e4e70c08702573ca57706dca8379ad906862afc8bf008163e14177eec497d8d9f8ee777198a3fdb5281ce6654dd26996310698d67c54893b53c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2173aad93e0367a3d50d300b9c00a6d53438b661d2ce2fab41dbbf5c7bbd29f4fc7ebbf93bda35782fc77f5a479ee2da1797176fef97c91bd3984504fa8187a8f63b12f031c4e9014a1b3500f14698650e1fb6a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h874a6a5692a5f2ed78d4da9c4e8eb669a2ad4ae80109b87d6512eeb3ad0bcabf80aff9b8ef9a2f6d10cf96ec6f3f1c4b39121f270f0d32e8146c3f40168d0084fa45d047b056cd63eb82ba1c708b5e518e6940e7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h278948fabc653733fd61f6c982e96f5a378cb6fc8ea20d25b01fdaf9805e5806bc5d57cad56be3db138860181f39cd6eb3af5eaf485ad863883cd5b9894680156192ea260614533b82e78e6c172d86c461ddecc70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb541b1b1c1984e78eb8c041bb2792f5d1bf5be782caf5e2e89ccdb695d65c62a6cbae590381d778b3b5fd5cdee6c4bc79b5e0c53813f3d3171bb6b40ee56a3785aa82802630508a1275761e411ba85f24b284c4a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e170e939caa751a3f75d30d0c07de93a78b61fddc02710cfc0a65280a17472d15dd3ce189bc80727a45e4ba54ca15d0442e05cbc43064e0df34bf8e7db2b4c4d7614eb40970032ad9510b5c8765c88843ea4c45d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67de8a188f6ce51400b5059c8d42f71c69bfecbd0e1f3fc9a2661547723bfc4b4f7469088774b91167988d6ec7d0c20166bb423893a2b3642730e75fa930cc5c0493ce6709627e41d582e072475e911efcfa5da9b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb835a2a3e0787e7e203dee83ca4f407a3acd0615ffee835f54963000765d56ba562bc37ff91cfdf95e0f1f05fa0ad6cf4aa47784c0f07b7d3ca6c788d17dd3381c54902f6d96bdecaa8ef7f30568c05cf2ad4bab0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a85318ce10ae2f9c80915b8b553769ba6c5daf20865fde03d6ec2e2cfecb87de6b1ff752e10688055692dfc6e05cea989fa5c1f07d016a85d3f3593287d10fdcdd2e661a78bdc49609c07c5948ccc2aa6260ed89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb56f9bd42813571c78c49568af6b950e1f42612a6cb0b77ea24c0f3840b8433a5636a82de6fdf54a97d86458a23c8ed91da78c4f92f6d30dda6d86ea72e5c0606e4aba0cb5e9b95b7e87736de127608d30f12c036;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7286e2b8258c83bc9af0011e25636ada8689d21e2bfbd2deb0a9785c1e979c2a2157a4883fb716c6d28b94a40fab9614eef5d7d31c878024ae7cc985655a2414d625beab78ce641afdb2f5c58d9f6a029fa9d8bf1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bd176e69e3de7424b7b1bbf7c78f41cca80ceeab43478a3c53db945a692184ff76ae3e908b998b9b41ecdd57d8a4e51c129b9c50e15c4caf36ce25454ae78c45ac45e490519979253033e62e168d3fb0584c0bf9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb34908d3833b32cc05983a422b3b03413ac45f1dd1b65d9a48371fe39020a851fe4ecfd369197ccd05f26971446b0d0a95e0a457e699f240a42a4f009909f7e77474f8f542ba8040bc81033f72202ad0b8a96d09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56b454781becbd4a225425f5105cabb435b2ba22e088c5b5ee6f3179774e19e5f1f801a711beac17b1dfbcf8f00c33a770225364be205b6968e2b5e8d08415ec76147c4f1659655f8e344e2c041db75c3cdd0a3c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h367ff156c55cab0bc9906b29bac3b6099e72f866b3dd0a01739035a53d80809f237876da6bf89f97d1c14a6a204487783469aee5c002e4c8686f293f5761fb1758c73a892c083645937aa4129aeb07181b63d1e7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf745178fd1c98080d71318ea1b36c61911f2058f32978e623ffcb84c366f45b2e403bda2f7d84719eafdf52620429838c65afe6beab3cc985962fb8d8d39fc11cb5d93495d57112623a61389f14aafe9a5a39e0a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9803494bec148689a841021777068b6eab9513cf6b537c937eecd5efd47fdac312712def54f00c33716d893049150e97c4d14a305f4e3b242b9073fc50513d73cf32f7bd3db84843f72043165d2c3532cde3df627;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h278a65d12351888976fc9c02c0f3f7477c16f34e50e4c65a062ca8207c1483d89f235d8d553513e8a2f2d89d7e48056d0f1c841b9ff8733efd9f74a321fb84389e71de9c5733f5870738a79675063f4c75daec40a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf93d6a2a4e6f63a99b2443e63e4920fa6ed2b6d27d39b11c498f22c133a96599b58aa14f98ac94a04341b0d6e7da06abc20f81887d402df419e2efe24e0e5f37effee9618e732387df69348d00e5fe81a18e1c4af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haeecdabcd32b9312af325701d555029061cb8ef428ae94d94e693768a9026e1869fe6170a73bd879ac37047618a38a0972f79736437028698aa0d1d668eca9575dfe92814be18e79d28952d354a423e77ace375f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f324640c9a3f55606fe7258934e64d61ac9babfda01b497f065fc5d133279bd17c6a61656846bd2fb1b7aa66a2dbbf69f78d42297d56f9d872863c2316cdf02f50918d05086ee4253caea9e85abb44fc348075c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0a2448171499bf38b0c784bf76b148b791cd82faa6f3c5acc0b3c0b584e70ba944fcf472f07734b8e1947f4f999ea49d91d6d73a7c063847eeaff70035aae21b905c3e9baa4aa62e60073f42e04b5b3a5aa351a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4dd52b6242883b0ef1c68f573931cbcd708288e9019457d3515ac317a291bf1a2a5f412c954b60766c354416790d794c0ccc955352f31a57e2df8a6f396a120f1a46c1801187dd669c5954306e6948f2449664dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2886c2cc51b296f7607b7b62a10902a6be60fda61ea97864e33edf637a7a70ff0652dae788917b87f4e04dd205f7a6e598867fbb00bacd87befe6bf0125c6201147f002203b6cad99c51038b963e585997212c86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae19da7fbb890cf8fec76b38e0714d83f8c279ab82b50de177bbc982c6cee09faaf880b58c7494d5bd53e082461bf6fb9826991b2cc5ef26f954512a6b305ff12bc95820e50629a7bd53c2a2e7abbd0fe832a03ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35c2f0db15922f815a406289e6fd5be3508ba8e486b3b537f7914992badc2303341f4225c5c74dae5f50025b6a1187d90ae3bfbaa6d0faecbdfeb0c1c0635f115c0d10349d9db923ca50b9b194d36a842a1431af6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc35f8ce093ab4af18474cd93a5ee787f5d2176f0528578060795f6fcff5adb5ee5ce6753d005d54f3b33d9439cd748df310e35d84526cf39c69310415b202dc26b7f4da04c2b1fb806520cc93c642bb7bbf72a07f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38e72493ffcda34c53577dad0bad645434fcd631d4fea11fd335740c1e42787b3e117cc2b173187decf080fc06eb6cd1944b33dc0be8bbb10461c67f6fac65f5bff4beacdfd02bd68d716bd779f9e34e797e43b04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb02c9584ec0fc681b4f83a8c01179837bac2523fb285fd00f6601a2b5e36ac7f4df3f792c1c6e1763ae5903947418898a98574a118c2078198fa85f49a728a5d064b2ecbbe6cd70d0d0d730ae34582e0632295aab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26902669aa2efef194b996c3b9568976d4202bada031c0c4a186c4419c014a9b2035aff3c0f0e4341e6c28dbd742daf74eae6a109aadc2827ab0934f0998fab815c436eee79f10b22b504f81bc86c87e10485470;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ae1b358a02e35e7ee9be47a19770a2cd8796ac1a274777f2fe8d12392caf79ac69ad309e0398274bff7076783583e28c642f69b04405f863ef10247d1061c6a7725b8eb2a1e7901f5cf576adb1118eb6bcdd297f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb8df3a7457ae8c3d4ac7a10a52684219f09e358749484f5b6a2031244a9756816772ddee634870af555fa3923996da18782900e402c973080fe99b54d5a61660e698692b7fd2f03ea098401de7a65566b863c2e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a649e777eebaa54ed9585f3a38b6616f4f7ae534d7f8aeaa91ffd3cd6090ff39d8dc6f2cdd381ff0173c72fddf7e9aa822a972fa6bf666f163eb613a528409b471acdea746b6329ace69df2245221f29385d20ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9815e291bea509567aece912c4386ad58424d92965197d8abc14208ad3b17e16e3f3ae2a32403e037a02250e182fe14bc95af798e6657af92f5d9b752fae7fe1eec26bc09f43d968e5964b79a4f19f1ff0a61cfe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b766ec8880ffc1175987f4dbeb7dfb3147598293a7059f62eb909baf8cc4a3052079f73873c699245985f03273a77002051c7132278e8e4678f57b31ce9b6861ba8122613d875d3e9d35899a8ef1bb4be35e3ccf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed2c096387dae983ea0b67f9b50ab18e11cd5bfa89ba0c9ab5cd71262c285e08e8bd2d452628b50059a0159e82c6f33276ab203241a5390cb2253271a931d7f1ace4d57d85a8ad27da4f2167a7302e3aa28978ba8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc84e6c60410ec8b900e51167bf166c037f98991c511fa9b9c8c12d5348be8a58aa72dd15579da8f36ff3d1c67f681f58b47ce0c23814a8e3bf30d3710b4bf46b0b7e7f4c4a972886f07b1d07f0153d6c052620dd3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h825795e863f764d496465c2c3ff82e378bbf2a7c60ff3c2fd73207c5f5db2da3d1b096cecfab6de5e5d0386eeaba0aa47ea7d4847941d12cc41f5d5a394f8894efb61311c6b3a8ef3900ed9a363f212aa49cdaa44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63f43e515fd40e44c02a76728696745c9b82e08cb9b75300b7ae480e8ccc1f0346d44b8514c649ce593cacc8298e3a534817db1fce91679abbda9ffa22659b7651df99db15e023c025fe6175d577c608269a3d818;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b57ae1081f274ff5983fb11393e7f29062bc6d059f4495a2ac66908b460dd853ef937232a78d02e2ce207127169562dfd692182fc6dbe1fcac88534c0ed91ab9f823c6d382ee58e2677857d84df4ff2f45299602;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91efae9962582b39f960a725988fdf8e7bd34cea9f6f3b6c5f4fabe7b47914494c74c6ec609dbfdc92ce6625f6a0dea34ac9447adda43db9a770cbe85644cf3e2dee7004b594362fc1e4a4a632345a5168702bc58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75ef943f8341f9bec80d9796ee6f6204b55f046384b43e70192c17bf6d74b3884ccc612b8c24094925cf26505d97a8e611c155fe7d589401e9b6f5e278ad3da727277493efb56bf89db92c510189181bd544755e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecc36ed6f6284fa2e16f62b5eb7d262c6411a5b6441aea02613d5ca8f8526b22b68cedde5eb08bc4979334a4f8317586a1636061b7320ddddd8bfa4694650543b6ba807a2eb4641e64d0106a33d30026ccd284d59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd3d5bfcd848206f31e308a1dc058d5f629505c3b78ba54a9e49682047451241ae6e6bad0b6346792232fcd933847d26129ece8d5e52d6ddd1d8eee913a8f08b4cb5c0d7c96ca742746c2753efac49b31ba4d5b4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78db9fe20b6b336a9edac68b009ad72391d2df12fd571741392070a246fc5409196ff11579d4d5d6da67e266982c220957e1801a825eb0fb477ce4ae984f8d1b7f394f6b6ac31035ef72bea5c27b5ffb751486bd3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f28a2fcae3e735bd304c4cb92aa6369457c6e9c58f1e45bb42ad6df3f80cee45485dad7d8318387a91db6e9981dbf1fae56e04d785873aabd776482c1502b85276d2b62bd116304b1fc79274e1d194d0e3fe8ded;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha86e75ec7c0e5511b0c9dbf450e681e795dcc84b33584f702f37960f0c61875cb410f94c9b18a48ec6e79a4c5129583fddc301ec8d6b714ffe7d142ee2b748c7fd79c12d3d98d779d49b0ffa6f36344e9e03ba722;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45cfb7a310324fc3a205b057672161641e85877d7f1b6a3309055d061dff99309a5396616a6cbc7923e20bd6641e96d6f91883693fa243739b6eb886c50c266255cbae68df86ae0e5bd9e309c839cd3c01c65469c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d5deaac6298143fe35666e4528912acfe7f060df3df9171bcb337fc383500e0a4c143d5a7a287fe603fcf16958f9b7fa0c2a04480dfd4155e24b3184f439239636adbd17e6c15ba02db512cc4d20750d9c4cbecf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bae2e19e2ee0c014886b5cc912ec22e0521be03ed8be70ad4d17e74c69dfc8fa8e5dc264f56784e66edfad09e6e502883f0cae1b7993f5d2d6ae8f4a37e36643c188b3427877291193ced2dccc3fbd7f24a47ea0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e33819601c01291c7790de514a649594a87939affa19e82c9a81c0a291ea140841fe31b96414469dcc3caf4ec1a55a31fd6f498bea308b386a760156ff76402f733d6f16b30be2832f43adb84fe5770d2f7c88fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79002e89070b1e87511cba3159c40d01d3127864b46cd90bf42c5efb6b022cdd52a507ec86c9dd6c1513661ab9f84913131157d310a8455d263f185d7ac3cfd8a25336378d9e480fce08c25706a1a6b2415ee6606;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h182a4e31543ffe76793a3ded2be11c6b294027eef7d7d0f85c8b9091bf3105e861d2dd2ae62c9107f1984b47f0d262757cb3227659d764b1daf45c4c44e398e877d209cee928594ba1094c96e1c8e6a92bb3828c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34b5cae981c98a1553de6310a756b0111b80174ae8dde932807c9a28650f887f5eab46edda1a58b11d8178ed76e1bbb4f99da891129c845b89dc424c97a94737b17fbbed505fa701ce8db777479d352944647eb3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda907ec086c8dfd885e5fdd3f97be516c48e074e84eab3425ddc01a9fac344778f9a78cc7725b55abf921721be950f8532dcfa689db083d86b7e639cc7288402de3201082b5d40822ea852aab47bff3ed7b4606fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0a1ac744cc39b0bca3e5c7fe4b6b21a9525d579dfebf9aa173341f9e4dd2b2fb5a85c41ed499171618ca9d93cc8cce49084b894bfaeac21ffb7d3c9198a024521083d9b6b44de7e7b225b670008f2486aeaabe78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66361293a2d7b4ef5dfa35f6c1b20219ab8aa31e0168c7ddb5ce3abbcb074e1bb670d667c941f1a925963f608fdf9ee14a4c10e84aeb111b58312c325f0a612868504f8402b70be43b4168c3936d1be564865d6e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe43641bd0930f14cbc16d8d8a9522df4f84a148f9fd22765105a008e90e56c472ed58af6f9ad8ddc3267ce3dcd2a7875dcbe9f84baac1c66e27b6572481b6eaf85b9b1df47d51086074549ef3c28e3b2eb655743;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2db86f038be95465ada0e1a6e2a49d30a07e2934f107c00791f91768192ec4f896b6e33fea2fa1b7061910a530bc50b4b5d5b6be59e90070ea5b340ff885ff93beac6fc3ba040a0b5fa9cabe5b1c3b88ac110130;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ba549faad5e40af233ba44bc71ea91cdbc515ee08f0b5b7a29d3deca5e3d00fac6da24c3804bee92f0f5303dcd12b6d8e27e1cbdffdb316361771ddb30567d8b3ba054d5c134d9e2f4da4c390082617dce6ce567;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10f1854a17646c37cc5dc96598b286f94057fd6e30cbddf46115d7fc59fa169dd3d41cb43f15b9384bd59d220c864cb99211bff04773f91bb0073fb4406c0f1c8de2bc9f790c0ef25d9bb62c52b766321b56d6310;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12f2c08ae5476f80e566eb33a60a26490169dedf53020e231d4397acd86e2a520e022a36e05ebced7cfa5fb1349db25bf428c369db978b69ffff7509f2fc75cf8f0f962e7ca9d31e952141535156eaa598e555fe0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5e460dd7583d461973d0f835918ce8e467f3df619ef8c7fd8d3c2104b432c51d6bb6f7e3f7ee1de8725d5bfc461840e9773a67bbc7225f87f8825e3f7bef3e629bfb19477c8be9533c92ed54685f3d48b831835a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cc60a20cfba042ebfd238f4f18bc9086e95731f0533104e97cfe95a0b904a911fdb137453ed81cbf4ee43e2da04b3c75ec4bf38b590c47f0304a6e0f77d8b89ab98c1fae41814fa73e5e0b1a6bfbd52ae1a12614;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b54c58ac3f9ea8fefdbc520c393dac9db230bb107db260198fa685a33a754a278b3ea4f602c08384fe613c89d04c1660dde348d83ab2997f78b049d25ae09809d506d971819d6e9f7cc7d12587d3f872ec3eb972;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h402daaa294a31bd23bcffa81c06a8d77544c21a95ec0bb4f6469a2012308281f373251e7b464db598139f2d7495cb14a30af5362919fda4a85d6238e5e656f76bfe1b7d0ed994b4a529c0c663d99bdfb46163c009;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebb11a2ee2724247e5fe51867ad3a9433508a408667edae56a11cf81f78245b4e347052beb2c9cc936c3e23a3c95cbe5f57d42ba0f746d3332aa395164ca9211e267748247fca3c58b049215572923a678b44dd01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54c4fa93cd1b8b24e99ef63c9ad489ca87f11b3a905d1e393c1d50c93bdab7ccfd019a88f85aa468b7319950a4eeb89429f8c50251c167ab611d3363b7adc898e45b696fb3919a65cda9b9a8e5b031a0d4b85d0c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ea33234f48aa26c88a3af0d998ab992bfdcbe34803a3e2af0e372d48890b4946cad0a70da7f2d0ae2542e8b1aa9d0e3d0a1319f6371fd327d46495864025c04372e614f1af61a98148c054def32007ebcdbee5e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde730602d167f1ea119ebcffd3be136414f2a146e6d497fb7baeb568196d8470bf554ac283a0738609c965cab58cd149ce3bc53133afdf3e43e88afc702e3a09a0cd7778a3d50cd44c2a3e25190d93a94c414e4f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a8ad4a992417d10b98cb89b6139c24468dc106ba0e80f7d5c68d5967c252c5151af7df53a80649dda2d14e5d28f640e0455de8e9a2e51c11ccce6b7a8627b3c49a86f9db690909039c7118a3b967d3cb0791bd6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf254942db1d78fbef4ca396174ef7383948d45b82a985cb315fa4f3da951c6614657bd190974a904043641c31580c26b3c4de1d1af0180662cae89bbb24428cb2f44174719ff0e4d041437ee251d0853ee8bf9a47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h404b867da2f8023b81ff9f5d684469fbda2d7563a05b4f0e0890c4eabfbe94207286765626da05a8f4e9cd853a7e57df9fbc188947077b5b317de568f16cdd4ba7fbc8f1c2839a5a000446f9c429ae50e84d38195;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72d9a87a5083c72d3a3d221414fbb64d16930c36a916cab302f82d56f99daa7bd13eb46ca1b5b0d23cbdeab7b8eea1797838499d8d9bb0614b258c4c50c4d27a2c6d5527f18468896159beed62762489fc5387136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a88c96e47edfad9be6f4734700e5fa7a74f5c0653a417c015e75ae803994b5c58ebf71be41f3e9adba87f08db78305a7bfe7d6f87f8078a050e695ceaaec6bd2a5ed248152bf13b1765783f79431308e7066d5c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74c3744d353147bd897989890a004a0d973aee1b8f463904efc6cf2a230662a2804fbc23042bbbc6cfe647dfed510efac9c85503f42f35af57a20d25609b2593647f22fba1f20d25468394599f8c48782dccff58d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h607eda432a84011b08e25749cb3b79171ce24fd6aaf47d215d1bf062055d58dba4debc0723bd50213f97f3f2f16845726399d159a8279ca728c72f5ca6320ec92ec35e73305cb46ac451e3ba22a8d38e7a97715e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h462ba4c555db173f67936c21b34b6a746d2f0b7ff626dd4bab9ea7007df488a9d10185f5b5ca617ee2ad4e2f3e6528169a33dfe266cf7fc22ebcff92e19457a409f5452500fac1b06a79ebb8c533a0243c3948471;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b6bfdf8f55dbc018e27aa0aa87b00fd0dc974edc5205a07cd5ea83fdbe7cffd17ebb85bfb31e1365e7d10d26b898a3a1482fbfa906e6082ffc9b4ea970c74537eeb588a99889d4138498a30db0a6ec8d2ae067d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h474f5c33ab5de20e3a499675a655c529704a39cf8dedb14291b99a9df8e2a67c117854ef98c91d9554ff16069b777da9165e3cfe119453df90eaf779ec1a55e6072acb5c8188bf6e59d59c33d2f09ba72de918b67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb8c8077a2299b62ad93c4c85d9c72cd2cf6908702b20421bee2ac19446130541a01dd4b0b5695affd741fa9ac294f0a3bf11d90a97f74eca65019f1953e79ae002f89f1cfbdab550d9971105519553f3fbef4121;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35311d75a1521b360a0371a48cf86447ac4de90e2789526aebbafaca55f07bed7aeabd4a95f9a19d5e47df2b832909fe2223c14a52c73814dc0836418054efc34c4bcab7b71b129bf39c24adbe3a051da385f394e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h121c8846fd0d07d22e78673acf5249090efb9e84bc90cab7f119f2862ec7c70d3ecd4e111b2658f00329f2bcf33173c4fa52248a76e4257b67c0cab3f986fa38e36088fa7d3fa291c22f5296c0b7c41c4348ee183;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h593c6457cf9ad68dbf73dde8bf6b8abefa6e3d63853e512bc642876d55211a1460449eef3ec876b6ffe1b60416f5f7cae1ee3fef85ae4df9b7bda2134c81342266bf8e5c2bf172204e2dddf1673547d10c7d878f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf5c17d316a34d0709339a9cd85d5b6952008c69a70c548e5ecf4ee482161e05be048c8ade6b5c12f93baa17c130fb554d6212e228f8fd6883602d411d215e6a8b1d6ed06209df39e8ac54924d39ff31e0d14e4e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77a717aa1e964efb07ac055deec3fc0d6fcece44b51acb423f0e27bd19c856fe0354b5fbbce7b9210d723157fa323c002e0ebbe01fa60de83b1ad2f37288e6e0677a04d1d3ab87cf7f4a55fcc58eaa9d06bb9015e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5a65ddd79afa214a7e619bae5edb9d635b7aed60595beaf19b7481ad3d172fe2ef4cde66905df396ae6747d07f2af6df5db86e629b677ec2d78a4ad831e5f327fd556810e23d3858025346f35948c6fd5ba14db6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h336d70281764846aa1f7e9b118a2e36fc4e6858bf69ef00ad31192aa0f498085823c8b36628722044b9eb2d9539f9c558f425f57e8c5d321854257d5bda62d6ce6e840781b3b1d0263657739a5b4e56ad4a9402e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h811e0cfd364dcfad5e0da6390a47c3447c0d29bdcc9d4089b547c767be04f816ddccab5c91a565ed1d206e1c89bdfce41ae284b8f54f1492e25f91265f206f00c20dc989980f7e0db4a25e183364f5fb8c11349ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62b85fc4367b3aed3de784ef9aa84a0f1501575b61358f5f56a86b628415d012353c0183a34234de92019492f90e31ac4792a8826db82a38c8bc0fcc3a5f3f705a9f6bc0ab0e1858964bb76fe27d28c8499c9659e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf524ef1545c6a30c2b093942b27b1e358c5226353108571a21e5e8cb376f00cd1547fa62d3e83e094cf1c2a8a2525df66c51bca3b3583391288fa929fc2d06234b64fbbfe2433ec80719e8a4b29ece06a9a2f9dda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4066843e9650cb9bd049c70cd7ee037ca446162de70afa011c2fcc2e8a9bca10648ccd431db87be121d25bb0197c58b86ca707f16c30e9519a69b64e8d25486db5780c6db849c99136e32a594c74fddac808fad8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5dc0085faf45d42f61298c8b025b1b2df1f86a9d85e1661ff37252420e935bd9ee787ef72239657315e868033d7451b5ec7c191144caca3635cbdc660d5c175d5a884fc157030710d99877bd441d8d15768663fed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf7b96f938eb5fdd48c792e8e3d5594cb95504e6f64199506a258b5504192b26094311b0dac964d59b94a7908d03ad02528c78efdbbb6b03762047f655e6163f6801b3955a3d6f3e562ee02c82889dc6d4d55b805;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5240ea3dc3d99cee5f8d821b70bea34b87b1d50114edad0f48a23197efdc143ccc3ffdd9a78cc005e3ba7d4972f7db6bd080b0871439754e5fada205a8f5ac2cb9478839372ac3ac56029145f3f5ed901f3041593;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b56191d7bb3390adcf22f2c40bd5ff3a09e193a5db342ce3e018f97866ccc7b4839b72474170831b4a7fcdcd641a2f0c8b8ee7457fb253446a22809ce99e2e5ed0fbf33259f41c2e021048592694a54fe669a080;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa9a94185c410f63c2a076de4479189d3541d70bd4e2ce155412581ba26959bad5ee38b34903f1f4d314a5fa2644d6849641cb393e0aa53df7f73c9b0761fd79c2c7aeffc563c7d487a6cf9d5b7e124b4d36f4149;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb8893e9c80fa46574bf54758e05761b1ee40546bae70436e39ee4e439f58ef12566c1cf0ecaabaeab2e3cfb8119020617843c737b5f9d5d87cdb5b37e0e5fe24a45b62c9b8380089069b81e0cb410d4778744794;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24aa204674ab4cd328bdbd4854fedf93042b9bae39cb9d3979df01828ce3349231882b86057700dbb57cf6c8943aea0faf44afbe7dcd5c5b1f390d046329e285b825136b66c4801e47b34447a46ea87dcfb3c3607;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h439f7239efd0f9b5a1e8080cce28f24b067cfb78f7344d197b58dc70ab764fd8f7cc379cf3ccd96c6b1713b1f08c32622521d36b93e68529fd6b08c8b53db3f1b4083391e4ab23ccb0e93d436fdaae39ef3a5fe78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5568afa6eb2065b078ea86638c6f81606277ffca6f3f7b994ddfdaf2fdbf2d5c5c7cbd79cbe47bc76fbce24c2051def5994e5e49344560d820cc235d182a2b500fcbfbdeca1a766c8c6f329c31c7762a5cd7e786;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20ad56192ab4e5f373a1f0f01e3dbf82f3bbb840f50c2a3b9462649000d4b556bb23e8d5220714a043ef28724873a62790d8dbf81a5cd0ac5fffc5a135ea490633eb7c75f45c99fe9e2d2545a0771b7b711dc368b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19903c4e55795e3098f8fe738155c7249404ec9dbd89b7c47577956c725c99cf74854bbe04874110055f757eb3be186714be95a40daab0b841b07e0c4525b0de3b72314de815d28cd50829dac82a52645d8617091;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36d5ce11788f78686ca6c2c8653bdb5dc91f8d656a3629f42f7771778c04957654f94788c7be9d8cce9d57731e862335a292e72639661d1dd4a65549d54f73642cc40b75e326bba77e569a471093d9aee0f3cb151;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1356aef77a43b928b2897390e77552f9d1f17658c8bb2002bf12d62efff39659e1c7ead30bd0b3b2cffdedc185dce6ddc5a4bdf7e84c8cc762c6c0b06bce8cd039054601f621441030f5f5646263559ff9cdb6f02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab9bf4157423d7b46d1230b164ce9bad08f123fb5db832c27001dae54de0ed4b485081e7a5b8dc6528dc7b1d357d0467e77b246ea35db505589a542082736a11f0f2663a3920aab0b48090179881cf552ab36572a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he564eebc13b26f9816df921c89bd2738ed18833c13b14b0c44c7e7e9199b6d67fb5c3490b0acf964e98ad44e8ee82c6652b37cccb734a9a588535d58da66cda3f981502d2b2283b8558ddf70a78eb19aa5b3a7f70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd16fe11c00369da83e47653949b3fea788c88d98554b329a45f727ae3671adfb610e7e12f305636f1d7fff3d6ec6c96682c2547647b1168c52dc64a668191ea0c2b35782a4da5393f6850886e4b051ae2693db490;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2569151da3b5d87924e1fe69c765f7c07812e29ad1984473709b5362e125db6b56e0e24f6bfed9badf0b64f3765cfb6c225f060ebd88f236ed80f5862e9c4da75bce36df5971091b00d68a65a1e77c1f84a422ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5197bfa53deb065761bf2c71ed7da0286fcaec86efb8e3e0592b5ee53fbfb1ce9bd5a0755f5693e84619f0a133ae9c6e0716fe4f4819bbc33ecc078eaa357eeab60a13b11375e03069fccf826937e14f7ca245325;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8352f228489597288fb2329978ad49cb69cc4bdb330c27cc818f7e8d05683bbbfe3ca4008b87f60f559bf564021fe38543756cc83f2c865ffccea2ace9571e770a57f1fe62b4e66e0336dcac6ac0f655f6ba94a03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b861ecf854efefb095753ea9f05c6700bd3ce66ea51cdda236c203fc09c18fd72e1b17b8c9a7b749dd17074fef3bad9c6569c81d2ea8280ae5922b19f327abdba875d63fd7b15204d0b5bd9314aaaa044a52e74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h688cbb3fe44bfef3d86bb55e9d29cb6593a7e5a5b7110713186297f42b3b786fc13010d5337e27ff7b3e4de44dda72386bfe0af92b99e73bde1fa36aa253266326a4bc51ba69095ff11dcdcac6814be6bdd4d0adc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8f424d4205ec9f9bc2379bd33517300d085eeca40b66d22b3fb9e3646fed6fbf0cd705ebd92c48fa2f270f6c7542d52af857654c93fb6f297de1a13e6cf6ffc805b40963ecf8c6712f7ebb00b6e7ce7cf8547608;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21f66c718f24be00b200598f24b0172725f1954f1d341b48cf6dec848feb41384a11205f2458bd8dedafaf1331e1444ba3971e08344cc96bbb0bcd42468e7c0778bc5dbad001f703828ae6c55ecc80babc5623af3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h675ee572d878dfe747ab2bf8d9e889b5447c2aceabdd43fe4320f5bdc904890063b4b09bc615ce4346ca7176e8dd50bac98e168efae35a95cb68d13711b248131be081f4abe06512a3bd31c6345956c32e9ecbf27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha01fdde1a393c27d0e44da47496f4ff774c696aa80406a4951fa2fb367bf4eb1521a0998fcf32f0b15373abfa81e21666fc3e2c58b46bcfcb8524a8990ea474a6ab7ef98a2b029df670c4040159e7ce1f2af554dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33789713e39772fe4274e6ec31c89919de71b35987c6aba21789a802d067d454ec97ad0932c6824618c195853871edbd4f68262b789b3358d9e47a22a3d98606cf31c07c9a228daaa3f9f3dd60814ba0f8a729a4e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h370931b7936d0e1614f709286298cf262fa093c224033a95824fcf85820ff09ecb16f7493d2df5fc12ef76e57cd497b094b878915c32341430103dbcd47b353037f7944d4b79dc5bff6e9eaa9619f26b888af6d9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b36f5045828ef26901ea16ad58d7e25db90e5c31062df4375bfbdd123ba9deeacb6131db115718801647bdc0a77346345c58c28f19cbc50470599e1652eb3739b9e54219ead9816638cecd6088496c22bb5d60f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91ade95e967e597f256cc80192a1cf4acc7750a2d43e18c514b1edac339c73a094c8f6999780ee5ca754af8da3eff733f9f5150678c1fed3ed6e4b4aa8c73ac6c3222ecf8145513259e1e3dd431a48e6ff8647566;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78454c624cbe169d4719f2610414a0ac3882fc4bcaed15b95a134e67b9c3aa241d87b35a5446181d84eb2771014787aa962f808487a900e83b1542157737c78e46b35f844a9d2d16e19546330c4fec99aa927101;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1d0512eaa4afca725aa606b21d9cc3d6704ab714fed6a8c39561c1b7e06db252b8c58de601ec4a6f5476a0770a256e57d5ec6400fd5151f5e6081a3449206b46c485922458ed4521d1d44eaaedd899d36fca522;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23412bc47b9abd0700ca523574df01e1851377b075a3074f1d1abe2353e18f0118721fd5f7e2f006e335da3101bf6fb0025619e96214f498b2d2f28167b444908eeb9e8d46f4e7343c1bc8ee0001ae36e4bf367ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37d7d7b0b5e0d63e3677e07adb6e00055f1c7db3ab4072a2d17fc49ad777559f7e38b31b2270e5d467211d8e42ca3adf24e404349aed02bd08d0c703b442dbc78f39562686c04900a55be4db525145424554eb292;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h198efa688776f86e9ebcf3555480063b2eff5b7d0bc35ad29436d2588dbe0e2862fbaaf68d5f1fd99835425cd6fe73b00dc0c705849c0d590bc1d5d0af9f3df8b371614e475a579084539b6fd75a2dee2233b877f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a44a979fad6a20bf4a5890a0dc1d85d2d295f1ea4d2c2812b56e9fa4dca4593bc1987fe4243f1385cfea91fa3237c7bae5a858022afe440ab73bd51733ec50d660ef4f7015602e8ed771319898a828b75e987c9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6296b3fb62ffd4c82f026f86f4837e40c8698f8dc4751453f78fc52b81db57675584bbef4e9ffd7cb16b8aa724ea528a998b6cfb071316bd677175349dca9e409c301870d5c8f48a9e4edb51adafbd07a29612c99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b9253db703e733ab8665bd2702e41db76f8a49cdaf2a6ab3087a1b0ac20bdc2bfffd218bc325f617c4677f24bd87cb717460bd88b101e8a5cdf93c3c72c9615b341f8e8aacd1313978e0ca7e8c0669d9ab2ce095;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cc926b32228d6a221d01b76792c9b0db97f9d9fe7b6ff0326f4ec1dab5cda499165da07b101394c515f7d685e4a1c48ffbcee7274776c88ed4e235740b55562a010b0b608e00d06b2cfb45286ac8e7f4555ecb3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73f7db8c0a609386b8f0455107657d06776866491928229b071b9083ead650200a3f26b47d944a63efa892bd3e9fdfddd84556b53d94b04435895125057e9b1859cbf2010a0f8d7e83388e225fb5e77d8684ac179;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89ebbe54781eeb28e95926de991e5cdf4799ef34bc789ff8955bc48af22ef851f1a3338125d12ff1058d071885545ef59a8e4e91627a407f85fdc195c01040b9c39ef9c9cef6396bf5301a3ed2a28c041b9f49204;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdba85998ba12282bef87c9506a7172e9e242b6033af4df2f249fbf976bbe9bf99fc4c36bff01858e610706f2ce61b895c51f603c46e745564beb98f05545d30e90c2052640b98210b3e5d89323514482dfbc2a7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76e2db9d0c677a751c67df8c7bb031c5b030c373877737ecc117e4a0b850bbf84d98ea339d408627af63b20d7f94920144f7e012eea1375136c8fb214299d72f7c374a2a8a8bb43a90efa8772b00a565a6e7e5fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h534c4a6d52095de3ea034734041476b420f6749c8b8d29a6eb6a383d2712fc705f8528d7db25b53ba8886d46c752c34f8d5b8df183500b3487c1435a789547dcbf22636349f699b7a705c1778e8b9923161d6d6d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde24018869ec44986b589608109530ef159d55818d81a44c9cd2c74024c5ff93010027cfafd9b31f948125d3b7c3f2bac61dbb21e227e2dde13e1b40ad6fe32b0a5671dfb6663fcf0c2fd14e9567c07d87cb53b4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ce32f18744bcdc106ef12ec8e93a9c0a300375eb0901775161d412646ef56f283cc14d44ca4e27528dde2e2dfb382a813603aad4f526da5e7b3ea3a6081320e24d3db9b6c0d1fef64a55c7f345b0fce0362306d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7431cc54c4d51636e69f4ac372aa2550e7f9cdcdf54a65c5357fec34cd262d7575834c4008cb3af8f8aa9ed1a77d7457f1a3b4b8d0954ea13ef7573827899ce14d2957dae5aae04c8bdadee857ddf9e7d19168de3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47e45349137be2241ae902b40d65188c7e54091936b82ebb1c836bcc97b47a8dd70cdd4ac46378009ff5ff24146d831dea11e8d1a5ef236dc080d21baa5a2b471a967335be2ee39915a1d4af2a699c2e493f53a55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2eb2116a021c6bc03d4b225094219548127da6935d0e9c2cab044838d547c9ea595f4d368929657a893feb3f58b1498cb660cb90ac5f6e371ab3388f3f8139e6a94f7572af71f97901dc5b22d60680b0948185f1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bd9324f851052bd134dfc73676e638d3bdcf93c27f19fdbacd9e6d594dd86b60c2f05a1250a6df55bfdf58b2cd79c0ace389b9013a5936393300fd7a05e8b34e6fc44cf30fb763bab5bcd76c1139744061e96432;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fee0ddd6f345025446c50a1bb91ca1c4852eedb732a3dbd5786b026212ca980db6cd05430c393a8827ed7737e26ce9f9a2d1c97748a0123dbe2fdbc0b1077f8264c350e8f3a6df51a276c3750b9dfd61ea4420d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc456900012a4e4ef76a828d74100e6f426a950e90cf9397a9e2ae7e30d0b756888a46743a65a2e7939b2036a75f3c840e63614b7d3631a5d058d31b298d5ea7c58805a286089ee4839445cd898e6c2da30cc97c11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dc4ca057ea7b05570976cec967bcbc4cf000acd933c8c9cf6c2b568e31cc76c63e1b361e3f9257c717cb6e32bf3c1567d1599320113cfec40af032e2b17bb398047a646f2f294e9bd010d2bfea17be6a63cec402;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9abd831bb00a14f9da4a75434aa9d861affcedb17fdbe51b735a2571b05f6bc87046e1c2ab98aaea3dfd8e1d2e0bc2dbe4d8ce5529fdeb809b714c6de74516ed293d6c2a3774d7e7be998b848392180fc0fcf32eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d957d4d37ac34353401fbb2a23890a142e80d3f41ffb6bd47434022126546fc5d953f4cc8f27498655479e338e67344ef07f002f1383cac29c13d0012181295dc6dcc1c71b1388feda6172ca100202387c4ed6b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39fbf75e7a57db6e779e401e367ebd9d22d32146b0746c961cf631ee374b29457cbe56b6c7988b22c6791bb500413fce4c430d41177d5f744b490e1be2620d922bfb02a9eecd40f8a5045a262611486867ccc06f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c2a33225d31ee4a6970f5adcea92133fece135ce55929cd02b9d11005d84e94e00da37e582657261b5623735cb9aaf7a74e0cdda14bace53d0dca9a688fee5c8a7e5ecae4506bc777cc5358903aed5fce93dc5dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8059d8af1481c13fe1e6c679622e7642109156588c14cad32db00140cebf128175613b38692e563845efaa6949408ae4c852258ed7597a66791bd566e1bff6c2ffd60bbd28592fa94a6533e4b6997751d7de5a09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e18e69305bad49aa9f7ff45f611e91829aed8a8829fbc88ce7d8dedfa3748f008b0a05d4b940b8cd20d8d49703993f589a70e37fd340bd5286d47736d6ed4914523ea4557a9f5940c92d391109ae935a21f0cc55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafa05ea15cdff0fbaca3444daf3ad75e01edb9f770eb8486db5eb38c9936cf211bf0bc30285fd1a7ecd7c73eed67a1e8e85025e3b97718e5cc4fd7620e6e151d130735ace09a4a684e62839f2edad65dc3253dd78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f60f524953b4d688db920b6dc181f15def90bea25030e508b52c818953bf0713382f4d71999764c47505ec86d0cd2283226d364041555247b38c9f8be936d8bb7a104bb50bb623169c6787a4446ca1fe0eacf697;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8bb05a0fda627e4f7d7433b695a5c5f77d375332950e568d19e58e36d0b2db389a73bf84500318ff44593ab539537c1d14e3208dc13458ba0c88e2740d65cbdbaf05759f50fcaff009766bb6cc5af1c1a87401e81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66c2fa04b6de106fbea8a9d057105b129c4ef50f2b1f3a3ea5deac24cf6b4e00b5ca8bee87a1c83e60f42f16a9503deb4aab11f1cc5a5b42f52448cd149ec8d29af25f4f5fe791472d9cce6a3d50c6d07076a28d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd19ebb14d7f86b9872298c0f3e977c66186a6988beb931d2e9336dc546e028e38fef7a71bad32275f68518755ced12e1485eb9e62676ed655b5683c3b02a5efb19c557523e0b76c991cef26850180fb8fea03cf4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h122faf65d009f057494ef30639a80d070505d6f77a83de5f3415638337feeb382afa93b96ec774b7012754a50f0f08c373cd5552dad9836d84e33d4b8d05b81900137a974a69e563e4bb038fc2e0e28fc003fb5aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3949763532f0d6dd9827cff4756d118d81245ae854f478a908fea4bbd286a0e345e1d57c944d6c737cc4c163526cbdf90c820f52344bc27bbded864d8a58b42d13b2024ec877abe393f8fb0df739c4f747d916676;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9eccac3c24651e06cfa568790d9355d15de7e33d32a64ed03bd9674d34eb52f36cab385f9f445131448ac2fa4441cbfefad8564e436acfd52ca1d5b14a584902a24ad13973e8a777f764312b9d08049c562bfe2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7875d9dc3e8c0a198f8c61335af77167dfaf89b84ad2c583ef32e0e1621146dfdf5ae986d7364bd12585fd0ff520473606b264459fe7310e30ef62c00af4a8cc751b129b06a474b0fa5380f507adfd90f0b7b31d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6792a1afb4a8fe518504d938bd75b5e658c2b6cedab64702467b8823965ecf9e2063fa582f8d93e677baf3f5188e31f1639a833dce1f58e452bd24c55562eae60750998fc9cddd49baf8fa93fb26ca1cc61641508;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5905eeed024f6affeb45eaced18c282d74eae8f48374ad63c725d6db248524d6a63f0ecdd71d4a685b4994659db5761c46ccef637bf438bfefddbbec2301d475bca533d91d0c3ec977937414817bad01951be9a92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d611d0d24ed22a6a5afd593fec7661275a3040438ef978bdf1ee786ef8b2f2b96efb39627f7269837f47418a40bfebd2dc3bd344585f5258dcc2da4bdfd44e94484f9157c4c0eac0ab5c469040f483c462003fef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bec848aaca1dab5a8ce4a33e0a3f50c42f7c5164e2192d857511dc7951544f509a029b7488fc2c0f7a97b33691778c9e77d2c73f5def2152b582cd8491c27a8662e611d8192c782d384869fc285ff12e2fe50424;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93d9450ae8212a6aac0a5cea24759cda130708bb6fc6fbb4d5889403f9ce3b219ea6e08157ff5aa30d1a9e0bbc39f93e7bfaa0babd939deaadddc812ba3d69095c896d7eb56e4972bbed529eb387c57caa6c48b23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49f066973f19b2b0a7e8ca2dd9c84a68f124d2900508ae72da98b0af50e1c66263aaa4f9b1f6c7d50bd6240fec325227d4d99105827d9bfd5708711e42c66a9cd805cde824da432edb735098b1dae7189a3bc9f11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d30f9ea66af92f043c328a73f9b42434e4d49496d36353eb9a7e3f45f021c3edefea9c449090befef381ac8a1ece07e62f721d3ad9a67d5951fae01891ad8f75fb5d8b5e97ac0767fbd69b4b3ea0554aee04e09d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53e0a3fda65368480fdd3e6cf5c3dc0c485889638d3e6b80ec467196cf9a947b4997f08429ed4c257b628e61fcd8dce76108fa8fea3aa0de3ad5a313308a2555b2198a7bfeb9ecd8d1715e0671b8756c45dcf6469;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72454b19d107e806bd23d2cb73feb1d9a80c936fbc0c683d3c5337676efde56f8f6dbe9abc1b2573f9dbaeafa0ad5c0a656b88fe2f1ec481f63769f68f60b68e3ac4c754b593b6e5dbbfd36dd339a2854e7577a29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cffce1577988511f79bcb3f637709c99c6119f9a9309c83c5081a9b58d5e1b6c2ba6beea55bb27de1d65330115013b9b976d5fd1c4d07531eb0b9f0a81eabc6077680f339779ab93c9623351e09a0617638761e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9f66a1a373280b648056c6878576226d8d79dff5415261bc5c6be91d858b0542e03ef2ff4a6f8957fe69d476de463d835ae9f7b9219e12271f17dad768b355105fa119bad106b48b3d1ad544c21d457540a207ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbce62351478783e1b43799fdab933d99fc9b4bd47da1178784d4f8d5ad2190365ac94e16c0d303b682414fcc50934609ded11bb07a90084de5776114a522f20d4035973547e2f0ff8984957c39655aca428a64eeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h922c7ca1009253e96f4762313bd1d5f1a4f8079dd51d38b57c54fb68765824b4413fac28d2d4cf58507c676b628dbd1cc8fb49549f626aebd0f2b3fb49e4d49fd467ba8dd559cdb4625ab2baef7ec074e05bfcf1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6173613d1307846b54f689abff4a1e7da69b509ff330e6c55acf748245cf2594169716398f52f5ec29840106336a7e647c7f41b4623cd4460b48963d0431f1d92a6802da5dca9fb1f7ad2097244f8cbbd1843156f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f450dfc4c81e0354be37546e126f43df2d1fbcba42fb70c9206bc1866eabc68bcf6b94d37e1609b5c11abaf74851ed56afb8124edb53e2352a077a7cd56d94c8981bff7877e3242169ec913afce96fef10119cd8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38216015a0fdafbda795a996df76e9a29be29c11a94fca168d4fc1ada1fb88d6ac1631b70e942ccdebae40597709501be25de2633f9150df3e586a97133ce4a2b9beebd282a79914a77ffaf5ab03eeb1b5d3164c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdc43ac6645b5182cd12fab6d7b16d09334a84566842aa197a6a0fe3273220453e942199c877ff27e692c90158c7a2d31b8fdc8bbcf3e37faf135fe38c3b5c6823c51f2164dcd5a8dd4410115646cf4c4e3d430f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91027ce2e8ff75a49b67c7662c531f54bc498fc94fdded3ff5beddf96634fc9b784387b1b5fd53a3123fbd9fbe84a7f5add0bbc8e53d105f98b39aa9a39e3f33861f87b19b23e27c1cc9f97a4793b1cca2c767ce2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a573de929d7976d56cb9068728179e206b265d2c02b6c569b5d822f718747ef3c7389c6e54707f6f22b0ca5eb2198626c140c90c56031fa4c055dcc0ba1f3acc665b7b8e7c20be5185c0fd53ebf4eb1f935b548a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53b5671d614c28ceb52daa83bf4e06ee99f81faa5565434ba43bade51b0ef9409ae5ecc664313778101e1a6b55a88c486c722281d4091a5d9a2f45b1d4b560716591c2337cf01f9d5ac84f4061bf8cd9af7dbbd74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6728d240b1dad87d3d31c83b8a76475a7f5a19424cb9e733ea522c1e10e8c7f613204b459b172221b8dcee6424466fed249ff39225221c4decde381d6a29c87ac0c087734ae95ea155bcee8d8b82f8291305a0ada;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h946a7a4b7d4aae377aaba79877ca26c03a931fb5ac1614e4abac44aa8db1b1ef683069f0dea8b7a66345f9fb6045ab3dfab6935b56943ea45018a2a5d39c79329093c8b135b57226acfc76aa6cf2d176280aa8adf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd284ed1b9e62a4f22f27b2f6426b95c593153d25a3c9acc0a85e9578067fc094816e88973c19d1424c199182854ce18d721ef983504f8ce94c588d97b5d4d4d92458d001b437174f087c9c95e9a2f833455b78e03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h177dd1ed235df273385bbff585d4e5fe40553f68724b9af9396c80de5d3049aeb79880339132eb9c9bc673f968b24bbe433de95ddbeb76a3938d135e8becb9682e79801e547b8084a475370ab4d8f8173650503a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h811f675135da90dda167ff0429a32e7cca99be729f422de7c877f7c5f043aff470ed0be9ced163c2d147a442b7b5c8b9ae5ac5204e40bbb304b0c937847d64b3e1f7d5ec60685e44b11cc8e1b8fcacf67b2304b24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6007dc4b707ecd60e0c2108a3f257b0171dadffb0f978aecf3a894d46f56770074e1b3febc4fc34043e82729723218046436b382700764094ac09cc2350b3d55e3098bca19de035774581225a46e6765661e90524;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h380c558a8d6d53b59559915165de6ca1dbc0e156f4d4a0cedafad8ea0d8b212a9feb32427d518082959d23b32a59743a49114a0b3622f864dccbdf0471af6ce910a115019989454639d7b77562e85c7e98dac6b68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdebcb1f23673538347863e4ca8d928a69691fd4708cef141921383b4bf7aeb1b64525d1ba937436211f9443f3790d08243087fa2c255766df933ef5e22151d55ba011e51ab234fb37bda0ecbf1aae43f3f475f438;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a573e4442472e92ca5c343628694cb2dc4b718d8ebcd7d29344b45b2a4ab321c10e5eefd5a362a2571323a09a9711849943fe1a489d46829f1340ecbc93a6926bee0760d086ed0591257dbb494eedf17fbe5b343;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa989617e43938794025189d0c42fb5e07a8bae816504880646d8f0630f81516be7f0723c23da83b19f87015518be941f2f9bb7ae2b29d5d04c66bd6517ae3860eb772e4159b5b8c06d95da5ede4e39366a93b959;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9c3a18cc1342f92b5783be4a3c76f514cdc239821942c59729767a2969aa596d8ac8b4db5e489b479b2d480c3fa24ef848902a08bd9a648d8e64f3a102c6e1398396cb95da114db7fce74387e881566035ae05e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4dfa8ec96f131702c7a0670aaa0944acf22a71743213d857ff9c3f2fbf78610446f90a7158a147cd4520b8401c5710bf2c349c076b698378027d2297a182dd20b94571a42d48eefbcf31d92145a0f4cf8536c83d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b78f94f5ed52f40487cf20eaa64ace6177b57462ca31c5c07b89782c28aa1c4d01c332988d352af2ebb613057eed034f276088739ecd66a4818fed2778bbd8c3c35dfe3a23d4476a5bac5a4afe059fb5c2673fb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47c37496a26f5cd9f1f4d7f505602279c904b8a6a8547c6c4f5d8aa60bb262490a877ebd9edcea621d1b7a4f963e4cbfaeb585aee56a005618247d3393ef946521c5f86bc92fbeebd25fc697751101852392ec9ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79b321b5250cd0bfbf3e6d2d23a43da6a479bc830b1b4b6e60f8ed406fd25004bde87a7919994a37c3bcaf1d54af1ac98baa658e64e013608dccaea23ed7ce5707016b49a3bb48307759ed4ab3dd75fd31211e677;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47b1d12a4b18aac9f4643c6f1b7950ef8ba3d5479cf0d47980d73852e5da6cb4c3ed7d398d5b1c3994584356ee9231bc2f6fb22f4b901a85e3d2d9ecfa37e8b110fff10ad6fe4a56ff877936db261e6db2c5d444e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79f06f123c12b9a3d7dc7e4e31f4273bb937c84671cab5fa6c434472a83e431177f33af0b2668b3aa0332e9e9ef05f2a79c9cd08bf70e5cef9a057e1cb3ba0d03b6d862d6d99d7532b10509cabe3ecf1874df9cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h516e8f3620fea33cdd2225483cc0dbd6b53642ec36d07373143e25b287c7eee2eb628d52d698408a55037cdefaf32e940a6a8b9353c80dc45b1241ccbca868b5720972139dd396cf6c212f0fda7c6c06cb9162669;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h667e00c449a09bfe7adee042612979bd7d35399a10df16d0e73f811688723d0c6843807ca3b3c215191826bf2aad2ff757d596e9e3429c2764d99933603029b0ebf0bef632ea10e9eafcc0d401e528c1c19684292;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49fc2470452fb16dbc1c3767029dc9253ee3ad20ddc377d9e94f833764a0a8c4b6e29ef0549bc83c2a827453d4726132cd9079d255d0d15d82d9ad2c69454ccaf398c5b81b1cc716e1f5b15b14c0f8a7dd6e2c9d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40bf2b5617c00d834f0ae1c1ac3291a695652fb7fa3fc4684e37c974e71fe3db86ecccd2323de742964433c2727d45d180aedd383e9b37d47dae8af1d9373e5c508fdc7efd7ddff6b0f145a4baf65155b817f70d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46acf0a5083544de6c7ea9af7211672200965f0559564cafae5c001d3e19ae49cdc9a46bed364f0d8e726b9750fd731a99ae17b56e731b2bdf544c535233779095660466c03dbc4925b991b381f51fe5e048f9113;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c5a05d439db7e0f029f4778641990de5bf5f65d05d946ea66fd7343cfd9de86042657597a8f1847bd76a38cdf661c537c5b4ef0d8cb06715aac2524f84652e471cae0ec0f2fa4a9d322fe9187e86f25970163876;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb03ca0b75fcc40f1124316abb32d9b9dcf798686d010478e4c342a99cd997a25ae62bfbcc0ebe0541920e1849d12993a016cc8541459a14144c185155c0f6dde2576b205f8f5ac357991091b86d36071831eabdf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd88d712cd31012da3c2480acbcac8291e33184d53a9b07edb326c2c6ac9f7bf5906af9cf8df3b727c8a180c8a84219742b527f897d07b906197d542070bf67d2a46f608dff2ced7fb6834a305c7885c6668a8d27f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc392769d8b8737ba651e1e60da6a2b479b2d022fb91c96b6b0d899732cddd6102c86ffb32f639182e9895ea62ad9f4235afc1bb7892d869bcbc826efc7de3ffc66842ca47ef5d9ae99dcde55f2e1faa8cdcfe5bb2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0a0d4342d0caabe26d184a498ff7932cc0fa8fde467b4ed724be43a76399ac4cacdff9340ecb4b3210945a8288e8d8513526470651d140db3f009a9b0e7cd96a992c2ec5529efbe32fb81611dee6060ba0d0c207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf91793b1c1c3ceb9915fdb7a932b090bdbc15eec075cf1d52479d6e10cb03de3c1f3ba822c987d0f566c4d48860f3a0569a04528ea413579cbfef3a3b44a2b982664427d6c196d75e0ebf800fd5034c7404c786b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38a1d3f9158e33b5a91b5ff10e8f74228c8541882ee37777ebca4012eabc93bf891ac16e7899dda17de15402dfe49d5057a70354863cde56105a4018a4e7a26a3654b9081b9914560348abf16da5b966a6bdeb8ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4443e5c62e54a397c44b28bc3be803b8b7cded36b44d94a781d9e78aedc2c28dac308a0ec733d6ee69572a1c70d796f2e350a1c4487dd8cfe6262185c15e45c6a2c2d98c9e41383214ab70e77d520d8c34dd71e6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14aa9c2028e23dd1b51c181006ab3adad0355efee13ce68d6313a71028ee68754f791934b279d01cf09a3c80252781f149a8a2dfbfa2edb77ecf097fc8a6603ca9178c3a3828d3f8bc0a5e35da1fc1e5a973fce4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8ecdfbab36223f2620ee2c0d8a86c13511ad750b5f76deaee832f28b49c5577df41010ae65734e336a2b25330cb171f3db68d3a7b37427e7da88465b631afafe00ffe40a767a6591ef73b376b3e5fc94fdccadc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42e24b0c22d9aa65eb95bbfea94650658d1e89b8f0acfc94e5216cab31844f6388e2d1a898253f8325b59287ecfa078c9f768cca5c96d8703e204ad17e0ab9567f4ef7e5ef347cefa5a215cff423c70de45fe450e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9450ad69ec8b6872f648db1aea80e8ab60bdc6bb64c8e6e0808215b192b65422709b8d76b7f9b9a0fd1fabfbd9f3b57e7f441c3fd8afae7bccb74fe7da3f35af92c818c324ae4f8ba67377795211904253d19dc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f30082c1644d3f7ae11598917b5d6bf90902e34d918852533eb5c8cd057e71ad4807a600735176693655c4d5df0c470cde7607a5c32473525334f7700b093a98aed2c4fb9831e401bab7d3a47fedf6ec66ddff67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51ef949bea6503d563209c7587ee8de10d92229487a0f972e4e063506823201d07307fbd368691ab50a2c7a5e8049242f0096aa25ac9672ce33da7b2315695fe08b474157762c4ed236b095cfc801de8ac52f0e7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11d2eb34e98bda52622b662c0884684c4757e47b173fd13415ca24a7cace4fb0930b6ce4196640fc673a40901c5c07b6152d031b59b603b5a8d485dad36870e62f0a5b7c53639b4cec7ce52aeafa750f41818f39d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha25997b764a88f8dc10d52f1e39c36a2cf089016c08c755cac59795f3e0aecc892fc5051d64c1b939d912ef8994a9d82eb1a8b54a399bcab6485448f0a4e520a548c4d3e28636937a8f3829cd554d8876920db5ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6544b847f0d1fb8b6b0685f8bf925d65f7e48fabba62a5c79e925d698acd9b89db43db250e3ead563e2bf5ced4279bb02b6aad92c677a5fad1f60334fac3e914c833519d87804394c1258f8193c0676f809f45989;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h529da2532d1944139ee595bb750488c4d6d6474f0c861cbbad663021c7ffb3a4dc2311cad63b0952f56e5d6e38b7f30aab12d141a1d28f779c361f6f513d839b993d4619457f1db41b79b150df7f8e3ccf4e680c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94b45720914cf5242997aa9ce89332c62c827fa6d2558783252a5b67c872ffb89c7d9e5b574008138756ae7fbbf7018809225dca023c1aed8c2417a80b685a7540f54a0be1d871883e6461807cb3f647f0acb95e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3cdabb0163b24e7249baaefe1011939cbef0149cf1f2dc1da47419b0d30beb71f31ff6be5cd00be6996ff2fd47746b243c890282ae6dfcff6e8bb8cce90dc4991d41074bd85a5f5dc0b381df19baf76fb9b8b0f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc5daff874a117ccbe9f32e0148b56278ace385ca471a082c39f1261db3493f0083b50124b59daee8d878a56e31497d25e8b8604c7f399969c6a23355cae5af7b6a213dd5cbcf7913b7905f8a3ce1b130b5ca0200;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5477a6549bec192a96276682ed80c3d6a10b1e2a0c482f49a9f9eca23011bdb974420f1f74bc4abcb844f99c455e2bae87733700c2d0271057a0ebd85568889e26ecb81230dde725a1b62b58964698c335301553;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7926719eb038aba15c076fd1b007e79f8456c5bdc57e817a0313020383210708d0f830a5fe9d3d6765add59ea266f97a904653c5f2df9661ce95b8b0964e72e8f1b02e6bc856d52d8ccb952bb554f57afe6803e9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd301bb27e2d4fb8432a500e1446ea7a097a612c06250104b8268ac1b104b5d7e7feb46c60ab7da44ed1183dab4ec0433573f35ef96c3ad5002fc21d6a30382f0c6fab1ac3f19d6475bc029bfb058a8160c312645;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h186f26fe53441997bd72eca5989f9c8d6f3d553602f3c61475efe92aaa4e71e87f6ea95e71296a6c4645a28904f4f54968cfe1205310a0f0eababceba8cbaba7ce14ea1187082056e6f336db4b10b1dd84f0a4b1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb241a1e2d12990a6694021e916b603d081abe5e7f639083d3bcdfcc9dc72d0fa8f3b8fcc8a334dcbeac6975f51161e8f291e7de7393a0ccf23d4e6b33c7cccb038dcc541788ae5d016b516568df0f6832782f9e2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ac9cc0d585fe278d11978aca55ca43f27b4434e79d52789dba8d32a3cc1c606a72b6e07dc0e53f7bd84efd2668fde48ed1da53093727cc1b88c04e055c11034d86bc249f6765cbbf67b4e90e1487a9807a5b6a12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h235404b214fa130de6d27b05c8455eca000de756f2ecdc15f97dace7a62a0240ed4b9d53a79caac006a894be1d04bef9c99e331d2f321e0bb6fea3d43489e1015dd133f3515235bbadf3933ff744f6c1eb15c8aa9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f318c7576dcd79f386833de6e6589e24af9fdf1e810cccdc832f4e88154a803f6f3d18fefaa33fb455b3225408774649b74d1db48defa556fc8d471c5d4b1862166c8a2fe44ca5d70b363fa064df2e64b887cd2f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33a3d98b7a1f53c3141f3e897fa73592252c235e115f7864bdf7ce3d3b709973358edbaabf6b592d25489fc15283a891734f4a63765e0abce59d7abc5debfb7d5ce26348849d1f76e659d12e7a3f4781493e804d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb8dfe115a7f89cdedf6fb80d272743feab00d2629772e2071bd1bec2041ecd3e7590099384d7e13c2962a66b5f33d7f44069f24b1366d027e2703a94575f7f99ab59b8796d97b2ab7204a73fd0b0fe502b6feeef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe30a6fb0171ca06d47d92713108da208c8f406657510d6cd2f020d2bf2f528a3745abd84e0c12738720e8852722c45854221b1395008eae2fdc01ba0d4647b104c62adb8a463df1b23a95925a3d2dc7c1d585940;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e3b15b237ec4e5c1952d7d9289539c8b0ce1630c05ddf7981840360c6be5bc8adfa75a7b566e6bfce6d1684f12e677e1f18afbb7151e32a69dca3130bff2cbcdeaf99137aeb416b614a92e6286c8070d50241f4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44f4cb8f9f0e4686e56c77f17377fb1379021d814c60999eb5cf02d2db11bbfd2dd475ec5e307edc707360005bdb772a085661aff2c9025ac065de849231a456d237e9edf32a6385cf5ea32327874360089be6353;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63c8307424444450042c21298454c60f62e4f99a64440868c7f8f3d4472de1f2712cba23dc909c847fb27c9721af6802fc410fe9eef97af8eb80c80ef72572630bbdfbfd5fbc2402dc386c5b4570eacd19fbfce1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d6adeb41faffba736feee6e894a33898e676be8c7052dd34e23882ac33b7e84b822c2396304f8996ce5fe8a94a5f87667f0c62c41f0e2fba69546ba001de052418a6b6eea13417821f9d161fe6d3f362b4797125;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb095b519304c58d3de03067164c0ebb37739a3b3ad79d6a22ab7234046ca4659f1942ee3027f733b4eab57e7f35859d07b2539d624dbb2f859e0b1159d0ff67421b8617243489940b293bf6647361f5c85c00bef7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9566ae8c12feb713636de759ea6ef1f599b249c1428aa21f9479cbc3343f3b343e8dc450b46b01deb38b3715efad0f2192097d9a5b8b4c4e6c5081cfed1b4eae82dc083fe2144c593f2a441135c2e47e92f8e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37d40a6978b454a243ba23c50860a364210f094a9d3ebdc076b7d1016d12933ccbab214501787de314d1d14d78197dba03d0631b645cd26ab6c83252f7824730633bcaa4dd79e4408d51681b057fc1b695abdab82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4ea1136aabf41262753f6f2e097b9cb8abbf26db8386d7929861d008af968242ee8b4e6988d74ae643247a87bc4db6c2a80e3126e7f53b6e78ed429c788c996fd21457b62160c497d0613f32e02b252187470323;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5d354726f06005132068493109ed3d93ff945c6732860ec4a78a787d26af43d26615be4d57c1194566574fa9e23f0b171637d88657aa1370b6f39f826f2333d0a6b93eda5f8f1ce994e134f49e5c99f8330212a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab039e7c15b39883702446ebf7eefab5c149e072db0bebd2578b7b53d0c816011ae06afb3580b1083df16ae03bc3813ad44c305c8794954cafc56c11563737bb80bdd349452fddf5a29e7eb14ea73c60ddd2221e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa6ffc2f9d7d6aac2ca3ff5d5e2a524d42e56b4381a944991bc1070e96102d84878f4f52cd6eb374be5d0ffd4dbf6c499c0033c65bc834862f3f60a4f0bcf9c4e55f4d9846238c4f18d5b4a8ea7a5c41c0e533b59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82d112f2724fae1a600a6b46b010a93306988f8b1fc2dc265747c127bf336464e74aa6e9aac3df1b264ea4218dfc2ddcce5217096f2956b61a4b8d4d809f10b7870631a09cf66f3da52b5895ecee292aba86465ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbee267fc18cedda0cb15b8c24a0bbd0c25512dbd99b052dc2db4aa3a9172ee385cc2509e95ed7a5ce1c15b9b46b6c2afcb1d1ae8cf1d2adfa0d5bb0678bf067e8e1bbe4d8a0390b9b1d9ffa5c3d9921162c3b7be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87d81ae543d2f567f0f3c47243ffc2d72b5a6674fdbbb702d9df36b570d44e9be4d17ce00ae458625c44c28ae9cc9c2335cf1c81e4866fd00d216f380785e3dc7523e9bd4fbc19368bd6ec4a66e2becc910663e91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeb6cdaa0194e6dad61515fb671100a1cf3ce30f83a1aa27152ad0018966856ac764fd5aa9547607fd95b81268fd9a750fd363cf8ae3103ac888a7bf2de70426c81ada50302a328400f25443c636e7d315d6c85bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h346958dff928fe3bdbb261721e4a8ecb7068a18e98e772a2c626540ec4ab6e5a0e76873dfc4a913c8c6e4502503db152720fa21ad6a8e0c92c5be59e2f5ccf905ebf67abfda6b4f67e4568c3006cd33af0715dc0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84a962a5c25889d71d11799856c88a0a41060a1fac63df9af2db4bdab81172ddd5805b65bfd8747c1883ed95c06b4880a546818eaa42d59166096fec562f7137193613846c561ee93b464d320b04c8bef52aa2f62;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b0d3a6c3adc8406941da7834c30f534a3347ac929312676ed88016180deb556041ab1c967f79cec519cb9b7e0b85d1094c1b88df19dd8189c3146822e0c17c4974adc2bda81b52aa1362a82807001fbd3285e435;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a94ff2ecd7d91e682b1b2dcc25602913951d27f670e1916c45b55b89383412937c45d3be7879da77b6753b700121f047555f0738031373b8f8eb0ed56f7420faeeb6f38cbf0319fbd31dbb9b216ba5088122f246;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h839661656e238df579b25477224fb1633ed9330fb8ddce0f66efe47779de54234d03a7c03d9d95bc4d4b28bc05545bf82e06750b638e5197c00a4e6fa9b3375dde26796fd14d54dc8cffb2df6ef11dfb5c65bc3e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1951beaaad0f59d73870eb30111297b4bcdf3e54f3323cb95f4a1a4350d707a9482ab485a7c652f0afbce830a4798dcd401402480dc1209d9cf8901da3adbcf6c59258fafdb74f7abc3b0e56f3a56f4c42be6667d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b93385d181d03f056a663820ea9f9b0d67a1eb02d1d656748e6cb7dca5605e539e92d1f3a0bbab0a8e05c9e97050b27a6982f3e078b9404b87410f1c40f20893ee7929842b468b9f6296d27ab10652405e2e348a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4764b805f5b373f1502fdb03af9ddd8862829c3ad95284e5757497a9f9ac95d1359fda37dceadd4e559115ef2d91ff7c9fa518d55b38614cc6e2ba9c2ed926e3648f7c469fe4b2c662e33a878ae56b4842cfe22d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80db89e72d953a0df37dfef53f165705a84a65f15ef49670750d71ad290de90a8374ff674b74f389c04b9270dca982b79483f8008c7ff4dd1e246b41173299095939cbeb546174e364ff4e8eb09d3bd803466f22d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h158e0094178e07a6fbf55dd22cfe69444c726ba6df5214db529f21b19a2960a6ced06a20b619b041dd7e7f55da18755b562ae94ebe065d412e10e59142e20ab467605958b54608cd16e6db3ba0c57b5971f55092;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e84923de6e60b7e9a32b50a81f26f16015457d18eed2a016b28bf15e3d860a803abb0d6aaec9c86872078e08cb24f2ef77049963ae64ca3bf4419f13a5f98b31e3e7597836e874071d781d8d06af8fff001fe8e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbddc330e3807ddf4a5887e275e01e4ccdc9b4dae2d68c3bb5c999178e0d3d145e5f53faee4da78e514a612179f614f611316c8eb0217cb7b0987832cd680a7a103b8f6b8247a0314eb125b9efe83bf5554a2ce759;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b64befcf0cee07c614828dcf157a81f28fb0cb4020e3f98ff9c852ceb9a0fae427565aafd99f5069791caf906d4b4ef0dbcffa98b76686641f1891c81ba33885bc765c5027d4502ced6a46b563695d9793804372;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd47dff68908ce46b2e4fc9aa67fe005035dadbf65591ca61998831db9c5fb87831bf65a098f9ef9d3e2adb143fc411f28619201796e95d2b0328be381a344577806697a469672c1e4082f4f092c3b765caeb66156;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h126ccc99d851b273ff3bf96e0a26a643707db40802c3b8d9b74bfd965327cdf10b96800c3ebccde580434675d7b52a682ec9289fd7891643bc163bde8ce9dfe98fea2b756b78f6771f0f75db47e68d9ac44bb463c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd27f73541c5dc7032cedb88d89773e3c91c05dabcefd3a1fb051981a1c39434e802c04ad0002620d3c60fab4980ef6a51c968dc01290e1f294a3760fe166c4cd054f4c01ecfe9bc4858bf3f8540684bbf609b3c45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb83499fbd9e0a8969730748c177b6551e71415270eb4b5df33b3ed13ff6e22f9d8c21d81f8d7c0f1e95544500ba2bced045c2c7497283b5d623084e21fe6f42f3c6140d3a4d13f021a6c8b046da9cc707f1e2fd56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7f723a284164fc4eabb5f614cbdc29b55a97548f93104df37bf4ba6ee709a165839426e2668e43222f235d93b0f23560f04eeb8322f4ea1dbbba2be1cfecff1155560da0d947edae8fa387ea9b9e211e6e66d813;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc04583dc8722a1e27b8b3696027e57d67937ae3c405123358d3606f89597b56739974e7555e7e3eae296a4868cf1be187c9607f2a5d448a0434d53794dff9fc335de93434884099d40fc6be5c47bd4b246431a7fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bef1c2c927686252cd2d71af54109e718b66cb5b4b68dcd25f3ef68e187da316797f98ee2879548cacba55895a340295600094fd6f733df4ffa60ef6dcb3d1203971d40fe2ca1fe3e7fe6dd0941e409095dbb8ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ffe3caf1d0dd3cfa8f04cc13ac485e5566ccaf3e70606b42ea41ddbd8434c2f83e5cb3d96a8eb056c2217020ba765ea8b21c3bb1d798fae77aeec04437dbb1379ef39a5e526582bf74798f9cce1a84f29a61641;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h900b4e798a7209d971c5b89703cbbe6a04af2a6e8607d92cfa2d3b49415b58aaaf47a3e5f9145338d9a8b313dffd3dfb3c3963fc4fcb047bfd6ad75e3bd3021ecf807433f971d0a6ae5076f92838614a573a5ac30;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h169e697df471d1c00e8d7a4b240bb102b7aa1a36cb7dacf894be325b0d51b8d4608152b241c842fc512a2c7440ffc5c2d84eb36af02b1cb2eaa79823990ef04f2c4277f0ec5e7693262d36a367e9129de59d0219b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he654ed3b83c087a193900dc1619f92ad42ea7558e1611757c356827983ffb86566e1a23a460d6b79bf32ab15e404395b61a5c2bef90bda847e7aa221fbc1e02c846753bc5e8318e43f35b53c4bcaf368a86b95b09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf9201ec7de96f9ca308047e247a1d4e6794410c1196458b2f503ade155f6155386f06a978b3b20d9c6652165f29d80263d8e93772d62da830e2e279b3c70c4ec7ecfc14425b29154b37e6e96da6c7c681260945c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d70e8c82a82d3c81254cac054e21f749df535625eb925fd5a5660411345d0c78a6f15833feebf6b68abd783b37311f3f50894974d0e4608814f5c8ebb3c632744a4dadff971d7f6fd6d5724967741aacc62a2120;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5ffb6d4d0bef54eaedcf4e29c1adc3280dff336e47c9c67ea6c1dbd8732786b4665690518af127a314f5a3aae4218cd3edaabbe82ed2a7bcf34d9a86d8f078cdb42fc00cc922d4c31e374e78e2b1e696b0b1ff14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f166d153e7a0b7d6b593e7df3c24b1479806fd1c4e139b76d2c0ae3c65ad53c3ba12139a7b6068e13107fa683c121da21f3fcc57aa05c7961c63e07b631fea3a27d1c1636e8569b4a03155faf1fc82471bc735fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52e9d6bc676e6e93f9c5cb39f9ef402edde4fde0351acec1216de14e5fa6f2e814ec6779f04b9b575e4c4f0457b695861c7be114c93d1d2afdca5654eec34cbb44b1b411cd71f80ffae62ef56a6a6757ce63b7e67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h492648b2e40620473e4cf8704b8c6feb9e963545fb27ed9c8d78abc16dfd5a5570bc72bbb849be553e5df657f69a1c1eae6360864d86ccf16000a0e6e888a1b39fbff76e116158ba8a2e0cb5149fb15db12d5b1c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb547ab410fad4b24e358c9bbf5cbea1e99f391bbd08f54227306ccedb7475a11a372be0fd654ad0d959185dcd67c5a96a2be514522ec3db25306964ed6a583c7234d89254b3077ae8cb11905909ed295b746e8c50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bbdb49aa1f39257ad11f3dfb40aca8fc630086c841f9716b07259ee55adf1d095f3f79f5f81e6df16487df3e8356ef0ed0655cbf6ea5f0608a2b104870a2689a974b00fb699cb9f50b08914f0ee9b9655d9222d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f96c1ec1390f1056ffe86cee91c4c00a4806047915f1a33a65d343e0d54a39549bc9ed172cfe594c656221f8d09bfe84b79e4b0149cbd1f337dce5832c237443d82b72eac51c82fa46c441caf479972d7020902d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79b4e732b98b40292ef121a929547063ef154174c94041f4a93fc56bc56680c6b6bed816af2001a4f33019ac02000de0ee590978998667c8e08924f46934e40d301e4d2e4fd38893ccb00b4b2a8b62d314d4de826;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfacee70877b67b99b57f26f16216e339ffe7032fda3de0dbc4a8dfba240f1204f2f78528e43c05260b609311c458a9a05bcf386c09b034ac4a2f78f7c457e7d01db2826079ed8d25ce3707c26c96164f8740786f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ae066b9259e4940fb0b14deb5c904f79bc06d418b0d95facf285ae04308e2e60e74196cd634da5e8e2fffcea074aacca09df82362f9e4f3a470cf3bdd606d1e79e4fefd4236cd74d4c966c603009a5ac9d170671;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf5ebce5997462bf6ee130db8c4e4ae3407409b66cfebe0889d2fa53e04c52aa51faca480490ce7f356d7475b3f84f540a1157228d1fc775b70e12bac52f6ecf4e9eca7f4e56b9c5ddd8103a582a37133d0efe88d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca33351f95726d6cb8873bdd6d20c93878568d065959632467939064008a9ba180a8e4c3d8f9b9dde624d0fbf8331c2c6d2af38684d4c881b932f1aff7ce67346bd1f5114685f46a69963c6bc7465275ea11408b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81f5e853db12e8204dfad67903103bdad4cadfa8ad7fd0f4288db9ee54470c68beb1b7148b4e7311fc81e585fb7da71dde125a4e18bfb983bd406d9b1d5092126387d06f39ae8a13011d5ccf9a3b2afc4f187650c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8773de8be0957e5fef138cbbb6613a96e116f5b405e125f000c1233d4fd7e910977636c910e2ec1dd09b03485918baae77ad7c97efe5a462fd3b4263529e627d956d7ac40ce04a54d79a746262ca1509d955a5681;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc500a1e36aac54f754e79bba1ab8eca8fda1d1e04330b48e7bd72c9f67c3a36c5ebc18ef42a7ccaaa212edd29ca2ec0921723ebebd6f58f8aee214aa3c5c099354f0a641ad7a29c6e4e6ac6b4a47a432311d050ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc077aaec928182b5d51f1be1b1c4bc55af72d654923ce097e80f3f7aa6fd572fa6314189d9ef00e70f3b4aa787be1a2c6d5d9cfc46e65c26bab47c8a40f5e6e30ebf9fe65f760b0ce130b957cc23fae4bc9cd0f3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd11cba14783ebb5f8f58045412435772638d3e1cdb1ab2ffc37f45f79d8a8e68e9075a39888322e819c317665f258ca242c979f96b22b8113e5b45541615825e5f97891da35a3c8b17606e45c02f077329cb490c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e50ac502c23899b5237486c9a2c0517800c5ffa244a9c563db67f8a3d223aabe54b431e9769bf1933780eb12b3f4d6012434524514f7d113277493e62787d632d59cc0eb11933e5bb3e20ef4a5938544aa055040;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd32c238c88446967544d6758fe4ed847e603cb395e110561e9b2f5d43adf960df56dab8a34c721e69301c41eca74807ce27e2b024c66359bd8999193962fc16d15e9f27cb7d76399f40f303ad9978d4231837d1d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habc755097e31a6f6e7408582aa95b3d75bc45bf11ae992390ca104a7987c074b590302ff921458957bfaf1a4c582be536ead46f4ba2a758024814516e6772c690ea646398ccdfe883952ef7937fa7b607fae96b82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88f99b95db69275d0ce08d00d1c2ebf7d0fbc3d87d7f0c9257541d242cc75de52586216a16c0691a4751f9deeb5cb62b158c0db2f9ea4e448118f5642dc06651be7808e67f8fbaec83dbde9ad51111ac5fc2a6d39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95f90ee567ef7f64d60ea1a55466bcb8c5c54e6f9989dd41333ee86a9bb57cf6f2abd6a3d71e73bc659aa458e3a8c3a8776f16c4a15d513b85b892b4f4713674841027ee47ebc6bb3dbdc4574d7fed23a001e6ea6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d0c17503a1081b69fd7a2a5aedf585e114dad2df3e0670944c760fb28b53c8800ee300dd393e750dcaa302308614248e4262e45009748d4fab4eeedc68b97be71445b92fe9d349cf25682d869312bb78b234439f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3107f1562e54e450904b9a9f23fa0df969d70a60b1b49f032a183aa1613ccf7e7a84adfd7817abc96beab6993731bec0e27625ff227589160d69ddd3c4e146362f2667fe6a113b5db001b42ce7fd395d824151265;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6950255868101d789525056034825b759716c4f3e2355c95d95d7e8055859abb7f3347aacbfd179f2009b68d1adcf72891b0a4321bcc66c9b1a5baa38098696de80dd485e0376ce54b3c845aa36e707c8c1e6bc94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2225a76d405bd84bf6ecc3b5e4efbaa6d412698c65e4ba0ad93f85325afeacbb5cd0eeb76a642ca4bf7710041ea57c8c1ee13cea7aedf5eaca981771783f1b1e8759ba861ad6d3189ff4e0d28ec3e7683874467d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h926fa1726a0ac368555a74b43242f598a40296c2c543db6695aaddec7ad62bf70a36fd7a6f21ee777f8283aca213c994756eb33e0aa139b18c34ddea2a73715845f5ab9fbe4e32eba3af14a36820a06e9c78a65b4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8a9f8f71d92439e10a8eefc45e6cb2f2aacfc4a1897eb1e04ef8ce31b0c3bd7339b5651c3b095b1d1cc06242e5133b24693fd5ce15d3357dc1e7b412da6fdb0055e9bb426a6aa0c268e7ec229f62b8631144d831;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha71deeb6457c5498829089c85a783ebe7f6cdbdd9d842ba4906322a74f15a7f99621aa420002a9e107f675ada02ec28435a8b6902dab6f30566d4c560bf8d3b6e8f39d3ce3571b158bd3a357e6826fd882007a45f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e225649beaee0782b9c920ddba83861ce85bf54dc3fd70c2fd53207d9025d0ccb2834da2b3614f9204dceec354d71404f89987f28a9f8bc498bfb966607372dfb448bfcba4fa5bf7c0abc61ba8ee06ca8cfb7c90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he20c1aa8619fd5b744d8c7266128c36f9c35d51d2a5506a53e1da688ba8883677740a7adfa6b6efd162b4e4b3152f0c82aea8643618ec658534716103775d170f78bff16ea494e1259d290bbd5bb7e6043c27fd4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfce0a0617a90bc9436bc84f56a71b03a25b678927cd526263d02a36f250877dacdc68c5922caa2d1b2b1adb1fc05a017b5c8b7aca0e2d98a5c13fd7f01c862a06bc39b5c49fa7dc67ecd2faa741a0f97293c6edda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h753d7ab0cf415349af57fe16a7ac2c77efb8c6aa7f26e32113dbdfc0ceb36c77c92fdef2c075c2000a120c4cb4e33656a4d4c1ed8348efa8c81a94f113461f18c2bb653079794c4449c8e4071e8edb3d5762815c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c61ecb1ec2147f85079c6f5c37539382caffd1e19a900790b27d5bae4fe155e5782c530d448d463c804c041f99a1dd5aea65af9c2b20e15f28c7f931174d8f393b4bfd7ca49e3096b6b46e676b4d49dfe57d50a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5dabfc0fb8bf63bbed94905ed16b7a7314da77b669698ba818afc80e9ac1f611320d98d0f31b41aab5ca99bba679541ded5f5b3406138df8829fabdd5e23aa603b034f4d21fe417f46a999444b2daea664f4070;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h488e3970fbf61e11f7bf3ad7b3b307c8c78685146772a644046040d3bc367219d4f5c559d8be4da0e71804fd279080d64f9002b4c5a014bdf9012df94c6aeff69b6a452cd1f174d639349042647187c0670858606;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7998925e06cd783a614ea76075858b1bb0f10670d4880a45742d7f58d9e4ca88dd64c4a8be67a2aaeee60cd5aa07e41aa952c83c6fb5b22967601347038f5e7024a935a01ea0a9ee42025a4c5c8d8fd3a2cf8dacd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb99bf013c8f7a56aa91b687b51277e92de8ffc9c24960adcab12c940505b707e4fff68ff2495091d78e3f165809ed7c6ad8a1a32e7ec6778e0e14bf380ae1577b7364ef61df329dcbf7b4748735db198819074622;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb1b882dc50bebe7cba60d3868356f435a5312e4de0740ff831751eaa9cc17d6bd62723b41d3989b09a0667387929149b7565ca414433d325adb1603c2fdfd8cd3dd17bfd3664d5c5fae679d865d30f523ff011eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6dc25586dfebfa49d74461186071cad50cedddad1ab555cc436778b94a3002cd06e0a0ed093ccef7be5e62ddbd8c03330e8c8bece226ea1375d179bba2d0247bdf51da10f7a6d10f6cb956c04e19bd0918466281;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dd13f4afd826b2c15e86c54b14232c4d8f0c67f60f9841f7d80d9f5bfd437ef732500ab4960d9e4a183aeeaacd784f305698198eca1c6b0ee4e61992b1accb09a01a845b0bf089542cfb3f273dcce8042c2a76bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c7d06b88440f2c0c164bd79d13357f6e619eb1dcfcfce8f06abde4357b9f8c325544d1af7f200618127c15c7d20bf8e792ad138e1266497036fe2aa79c5a3ac42b406e1bf88a7c80150d5ed882398548e7950578;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31da4263ab2d6c0f7cdf592571b867cb82a57bcf01dc53bbf0a6b1dd8fed3480ed15feeebccaa2b37ba2725aa48f526472ccbb1596b745dc4064e701af8f53f2547480bb4ce1218a34590144f101c528472898348;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65ef85427db2e001150050a7a5c38eac7c664003a6260f6db3dde0c93bf7e251baa04218573eb6b78e09dadf22e0246b604054a93b2821ae0764ca85ef957f242f7c6f835786264193120a923bd767e419099e83b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80ebcee049a6766974f2fa42444c9fb56921ab64f57f229101b7bc2902ff108a5ef2acba8d8db4deba6687ff075da560d630a0604570e46be502af09df91d73ca47c07ff76e6a2dd296844ebdc22ae7110382ae69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f1570cdb31dcf466ef621d71c44f40f5ae30662a006b46a178cc9df7bb93f4344640620c9d17376413be744e529ba808ea20714388d09fb83000e691698d480a4395a1ba9d305ed90c54da58ef96ed26529d6301;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h621e050b918b712cb7ab9120e31855c5bac381a9d94895b7a17d1b61709988379c7c65ac0bf12f40cac7e481fc0cce69fb2e469c699441e7d9ed3840ddfa7fc8355f879f5bf1de90ee81e92730d2e59f1d2f3bb5f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7598ce3dbd858e8a4a3db2eeab7eb6b6e999eca2cad655db3168aff0e56683e4cb6658b9ace3073dc66665bda083158591a2da8306f9761819cf7f34918724b45f05bd20059a467aef149fffb2c15e42cb3aacae2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0f5c0c65784b089ccf7e29b90253c6eeaf1f20af78834b60c641b982b1add13410881e4e561ec87ba30a92599d15e123828cb1d8bfb365b6d9a2bf72f8ee3e06c9d1e44c40724de4c270ef7c563e1481dc5c3f85;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6d2aeaa8e673c673b0f808baa2a960cd6511442cab478d0f8391ffbef8a8477b3e3f20d70ab39eda6f8052b5db090320ed93b2c7b2f736d5a948974b03876fe1c84b18c6280e205cb49f1968639c1e9448d718a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8712954150b75e90e197287d3722e5e485a6af5b7a2bfd348a21dfcb6e147d757be043929734d4ac616544f109e96eaeb641b2b6ce66c4d363c4548460a8b26a9dc04d79d941b58d24a6c69a16ca66788eabeff4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1bc63c3b7eb925374de78ad210f04f9eb4d50c7ab61f97d4f11d8590312b15102215bbdd2eac665bc33abc4697904990d1b3e79fe769bcc86722dedb1c5d0198608332eb35c68bf6c5e9386de0b39d1081c3d85f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha41017fd5545b4d8e89971cd7c5662198388ebbe38ccc52cfa80072bb14605df2516ea416ae3ef10964427a79db0650f1e70f8edddb3b2fb520cd791e60652917aed113a2e80894c9cea0786ce12e64728707f45c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc05ca606251c745d8bc3002f3aa221501e1ad6469e81a9e8c074d21c85c90782e37f358d5b8e32bdc70f73980d1d2719f73c40cc6ceb03914a25199d4d185cf2440827b4723a8dc98268af00d08120bd75e69207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb609170b6c72b5ddcdbfb57be693bc47c6801b6c71927e92e32218b22f133ff6d84c2f253d75433b60de803124e7e39db34f016f424955ad80916f9b9284a77374f0e0a19129d277c8211c10b70b855ba7343a1f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaed94cc4217cdd4b9efb9d110bd92c29d3142af17e3ccbf160b17e550faef37e95fe18728f14a29e0ba10a0123ba90b774aaa5d98392396ebdd227613bfca59efeaebd4cbd9c07c35e01c45232364f3ac084da51;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1194d859c025c003b70386124e366491e795fbebe9b08c505058cd5085c9045295d9666a4883ef7cc3ffd0dc7c2a04da0bbbac0f2ff770c2f5e86a6a55acdd6b3a068948d007bf515d3e4deee01b1148632465d68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heae919a09bc576768b7fef5d05eaca65245482e728c418c8a9dd097f2a2c4c90994499e97a52f57f1159bfae81fa977459bbc6ea4c9bd494475f9620c937615aa02fe953870782d8a9ad018883c7f96f3590598b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3ba533f57bd5cfdba8cf61a86a015578cf86a824b9f20e58a752ed80756ccc10a6b96aef8fdfc762c36da5426e5e243c995c4c9e2a8117a2f1da43d7500311a58d2e0f5707925ca02f67ea99813c4c0f8925bb59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2472985aa129c36c1cb10457e5b3f5ebdcdcc01577df67308ab442dd9ee70defa1fc87455e73790237aec07facdc45fc15f1756099663b6fd38fb811de20f7e8456a9c66bdd2dca0aac04309f65e00ebf65633607;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7be2c84f1963051adc3962e8d76fecf824020c198a9ee5dd0ccd59ab33be0dd2eeb4b845eb30c91bf95bf1955633a0e0e6ebf4a1d8e3a1679c49429fb402aeceb05634cdcaa5d1dece640199388cfbc0ccfa2e66;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f8f294b3a64af6af9185e37ac1059a3126628346ed00f22734c2070eb82dd4d61102c35ff98592c63bc558eb344f4cdebe6f392333d986064b82f9eba40467043ebf6ea2d918c34901c7a2d2a9fe0d1a01830329;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c8372418e5def96d7b34d776accbada48dc207c6d722a2fc72811dd8343e032ddaa9afd5081b00a03b4833eb4dd0b8d8348a17bfc1506ddf0219c9faa0e98c863e1eb988451dd143845da65fcacae6b4b9466e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25e5b4852954c8e4eddb0017ce61cfb8cb9b8d8c094a09ea90acd0176f86e63ba707a41b659f6e5c012775f5c420d3eb4d80af67e894887051c137476c1ab2ede17032a74a536ddf754901e02651cd31be7604f4a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5030da18d0bf207d45e28715da0795acfd7c8df30a5cc6114404c468761968ca6568dc17f86a412c3f0f283e62474bae47c53811ec72db9b46033f78f743998eff1cd7b4f474dbe44219f50396b379ea6a5ae2159;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55ea447ed1d8287065e338a4a041709a514d3f1eeb7d062ec8facc1f543aabdba7a27df2ba3730996528680c31f27608a8cc0ab23e70e659846b97197dbf9febeb0744fd4c90e64f1284025e4ea082f4bc34d7807;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3a1bf7fed04802d0378fecd02eff97ada71d69e30d6ba573cba9cfab990f39381b813f3831e77ef3aa3a32948a2bd11775bc025e86da991813e36e35322c0fba9adf68835755ec360dc662117c0d6e1f3433afa6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b0e1db81e02472ba8cf5c562c8ca026c140fbabd3862ad99ce9eea177460241356dc0c7c248b38c3bcad4dee2cf39d9d3002b4fbb7162e120b1fb60612e5f67391ad096c2b218323307773957d8a3a27e2247e16;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52f8e0abde1acfc9ac75dd93e961defa004c21892da22292ebd5ee6f20e4e72d2daea88bf29ce6098988048cc76369d1b99bdb5736882c1a32ab4aebc0c74513ef9a7ad1112b447a34088224ac85959afb4f10db2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb315e3ddcd424f0193cff84ff69e33aa2e828e8dafb24371815db89313bec3014ce3269eb05d5402319e3123cbbd22113e9058dc07ffc9a63a96f10e0f9ab78c8cc49a216cd86f8237d4872529f9cea059b315241;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43cb6fdf4fd0bb0c334fcf92dd7a32e8d00c6a9a9dbdea8ca3dd72eb7e5915fd5c408656cd7edf9ddca4d2a03cf6dcef91871434e607474b0819078503534ca91dbab24efa0ec4c5f8bf27d495635821f758b0cb3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h130690fbdbca68a732e9eeaf0083c8452ce8e71a9e320331c99464baac849bbe68c4a455800fe90418554a57cdea144d6b3363d6e84a778fbd4b72897cbce97304ad72ad6cd2cf0426be6c3d2c6640ba2560136a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd26b628c301171d27c46e22b905803860f03efdbb6f96863a3b8b167d4840d141c84d0b4ba42ac24aadec087bbce325595591c3487c0f045dc369cd8954527dfa7d7365a9550464ecb5a5b5c77ebb081a5f82d7cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc523917e7ee9f222d0a28809bd3e18cbcb5414bbad720bc62d2c725d211b3f7c7a02f15c2d2b05c0150479a2da33452872fe71d9962cfbc8e101b1d7ffaabc7d443202e2569641d0bd5e4dedb73d06aa1c4855efb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73b05d2315418816470082f095ffdc9efeacb19f08d3a5d0a879524a9dce844df601bee8fe69638427721385bf54b5bd53f9db59b4e2604c953e6830510234a9b704a2f3808f56255e75610803b66c2edf3d77c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f085108cfb77e29907271698488ccee25b2bf2a83fea212c9c226dc2eb2ec247e56cedf2e42db7c441721a507d289702b302f6d9034f9c6bbdd4d31641e9874fc7908c698d9d9893f4024ca46d9636cf288a9399;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb33560b1251dc3fc93d766356aaa2bf02e0765ebdcd7b6b2438a1830706e19269c14abc8e00a8ab0df6628b14d6b56a9d1a08b7288cb8aa668ac4c51e5b641e793a710b4af8d4ea8029ac0dcf469f7b227f2a41;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf321df76556ca40d45fbabafcbb2b9dff5426f62859b3c3c069308ce4d4b485db3c8d05184db2ee70275a92163a686391f640854b5f434d5ec140cb21dd85cde6e0d16ed72650c34b7093611ccbf0c1430bf67557;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9972874cfa1cf887be3de721c7bc28ff00ebbcf0de905f63f8f9b92d876ead58b60a60146658055fa043e3c06826edbc3d51a17dd535df9ff37af79dcd11ed2fcb5920b80e7dc8098bdb80b9c22ad068fe808c24e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6b80c2fa3f9cac305de3e1c37b8cfeff4aa6920c5647ef565fe579818d92ee9bf5a9dbb4d306412094047d6b7e14fac5812b0e1eea8e692bd1a42d661e371993073db79cb32ea058ed6ad573feb05443274d667e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85f3e82f4542fbb5f7a4997e863ce6b6f0c6dc38a5c577c4b161686d3ecc6c7714bc149d4751ed9708faca72de2704a6466feca8deb514ac7011c5e29e99bd31a2980d3075a8fb3d8aa2e6cb86a8e4f1e05bb5798;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb9cb87949c22502529250666debb60e6a2ad29c87ecaa199a0e101e0b7a6ba06d3ed23b562c196d5e3c093318bdfbfde0a67c03691d868ebab55554cfa20364ae799c5eba8f4b7248c180fce5843f7645ce5565a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h288df03449f3242f7fa4824ba1ec470e260fc360bc0843f9df628a294e9bb7c2be0392b5c26a988a4f11be70d559c9af337b17640f27b0a20697ed3d35e9044aea4053304691284231001cc9198e53ef986a35993;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3ba528edecf3a5cdf93ad0bc7956b48eb4ede41236fb557441dc3ff6c324cb67810777dfea35fd731492103617eaa61a286bdfb7ca59375f56b8719f2601f837ff68fd03847e973ef894c4e8b8b32a8a70b87d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb1ed6ff0c173d28b8fa947338a1e6483d0e8e5bf2c80d0236c62e108580a4955dd107552af21d731f9a050862f7fcb1e4be31cc934a8561c24c8e32517f87fe7fa02887aee21fc24454445c87e2ab46747d5e466;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab9713b3f591ec7b0526188232b48f756860f5ba1840060384d1be37c9d9493e9b509e369bca6cb1d4452a6fd07a9fa7cff7cb8911863a90dc6d7dbb9a539a759ba9e5020c10ed4417eb2661012b94e9d46b63f55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61307cf890b7bf0f3c026658af8eb283b4816a9764ea1a67c316d781d48fd9aadd89576a32ba7e0719780491b7cdc879edd3c42d1e1ececd09f3fc5de2c220f225a05c8b11162a28760a745fa53b76956f1e79654;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde79a24f7222140fbf209d90f7d8af83794096d8edcce0a458aa9c7696619defd63b5a969f593a24c821ba6ad2a22af7b23c995c511c735ad7cde76f485f1d96be3b7c47015dc27cde184bf0f19072355da98eaef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ff2a3c24bee873d03ea6d0c8b18413dc2d31df05a6bd702bcfcb45800a7dd59d677e5c321244059e0f270ac248d4c357d6e176fa3db452b6cf5f5c6d53be18eda43575b611ec08d97c02f8dbd19eef605864baa1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca75a65a88d5f354f0bcaee9b130d7fa1db445034c174bf67728526cb05b09bb43181c0dab74d640fb6af237180b6598343c4e8e2b3174e6ec709b88e3c7b5337835f6406a7fdee813b7ae8edc3a5a225bf3ed486;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h984c86459be9d5276badf7e3fd9dba4a956c0931c8c370530f003a801188045e1e323ea53121b098c506b2d6f525547bfd2452b8d156d827c7963c4f2f29222670be187765a56662214e7dac2489010ad3c4dd54d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc04073b07d65bd9b43f578c8473d64f55df542226a4027b7bfdb4ad652d4df84c0977808e23acc0cd76f55b0bc18c2a17f268ab069150b253e6bc08f211bd26edc2e8ad0ab6cbc3648e5465bacccd3fdd5b896e98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22dae388f2272bc664d2c6f446d3a1ff4337a2820279847c69e1da4d8396506136b48b7a3312ccb0900081323abc2af7578d9514ff813e68d7d205cf21d41292ee9f766a2b190eeb75525062c3d6d0bc1987f04cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h797988482a6292f0da39e3c3a933317ec38dd9d9880854579f73c9fbc7e92aa8823645e70d790eb5947b58479b133b027e3ce41534041a2f7d6859a61b7277318fdccdb89d79c811c3caaea09e177c85d622fb362;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd325f6ab40946fed6ba19758123531ba2a2abf5804853a3d554d3a3e113763f66dc5a7f2bdcce79bec1a792e1b804abca48c98cf397e3c9d0fa5a212548eb4e6e8bc0f07f97a6d803bc155b482702ab717093937a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e884340cf79515d548f0269b37a367e6aca2dbefbb6e1dffa22962ecc98600dd7ed0ef9762c43a7c8c42bb29ed1cd76a66b1cf50a757541ba18971123cd790c8e9a06761d8da0c339cdf3f651f6c23a20a4d5a36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b661a7dc3d4ffde3858623807b1513c886fd71b09bce2cfd031a6a08ab48d6d04377ba058361b6aca33d84979035474d9ca7827b02787972472a4d80b33b40f855eaca2a77adfdfec5e7729cd7e7e2267a368909;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf4020a8da48634e5237700481b163cd9a2032c9c07856fcbb51157b8fa7bdd64cf69ed00c490121b02b4817381d0ff791431d006efc44196ec07da126d44004cde890322a36ff4da74fbd07d0540aed0228aeac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcdf8a796df2887702da0cd8b4d0992a74a6d575bb54de1a91cd6677a0ad2a5bfe5ca3cdebfbf936dc84cf386677816f593b7e9b1fd596761c73804227b8cdef945becac4c27ba756d664c6d53dec454ebbf85e5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ff29aa9132c0d4b6c18af5ed6b8d77068d438f79cbb8681abc87493cc5ad30437f1a4e25db1095204f9a210b671af11312a75b6886dfbb0b6a321cb29a261640868f3590095e53c503f2a1cfbd1b16cf88e631cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d61223f8ff325abeee54ad8ea1ee6761de8fe583e0e1ea14482aa2cf466149d58ab4ba2047a5908ec0f91e95a4b0f115abfc9223a31972f767ca83ee47a384df5961fdbc7d53dc6eec1174bc0f16efae41af4185;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf294ed3f3671cebc859f95017e967e103489890874c1c1fd161b4b8d389ad4c3d930d46d88283c82300611b47522a86fb228d86cdfe72c2951eb93104a055d0de3bb3b7f014347706a734e66d3391617718ced52f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcff8b84cb1d2770b8b75c3aa4235239e98ee46233af5c5a5336b8c29dfe81b3652b2b0ff985fb526c8adfb451746e6bbf2b38b43867a91eb3793b6d6d27119f13168f09cb3f19c3b86d38c9bf1b824c922722c387;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h560cd141844f0d42d18425c95a7067a7dead8ba9028e42d44a11671847f10417de0b004d026a2cbb6ef7ab066853db204d859904b229ca0c0cbe1cd6d05d26749758564c56aa81d5f51335628ec847134cebb537e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc116cf621eacf952ca65dd296294f8c0aaf11a07298eb3b6ec3b29b1cc138775ae6d472d0d833c50fb78154061d868132b3cd55ef0f8d23bc716c3a3f6d107ddd9e72a21d46de15c91f314ca2ad2f0e53c25990f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h183b3d7eb54d040a95de4186f557bc991c14e1b79fca7fc51908bc68131ada6bbf97d9ba59309a32414dad76a7ed6e9a633d83484292543809379d5c8229c9c9d6e85d6dc911aedd71ef68e276cba666ab7ec500c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b0963e5c7ee0ebbee351eb6ebe9b3f91456dc75bb5f0e3b28f4f940cef57c5e836ab941fdbbaf34d79c1e097f2b26923ac1010e534c102bac3619b341522257fd30a7dad3bcd263e93e258b063d6e2766aa39890;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf577c05c12294c441fbf0b7386228e790e1af4f625f3abdc8f7496fbf3c6737a7f5df16745440dbd8622f9118fee1d7352fb56a3d47756dd49a0c2ceb06497d267364e15238412b8d9519b9ff56a842cc7e418e87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18ddab4ac4152cc3de3814bf889488e2b2f8cb68c13a1b7b4473cb7bd8c249cfc497763e335c03c340d36139360cb0f77ec81df65758741ecd462f3ca929a6147a62f120b3855e178af4539bd508917741bb6e124;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2fb614c785abe80e146615d553c95f0099172c9ceeda0360ea162f21542c9b16e4ce8bba55d812ddb4a4ecef074be5337e74cb6239b6294795dd3b455e7962589d49ee493bd67689643b6adcf3488615c10e3052;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he20b94e112d65147f3542c0eb8c08bdf4c7e338d5020ae77b8afdce099bd4c771fe9c2dc13227caaaa0250d9736ccbcf1bf1113c48a544c0997cedc6ac3c70cde37b3b4bb75d70815c306413811e5bbdaed517041;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h771604aeab9752e32e25bb679eb21312a2f6283a8ecee2c480aafdc61749fd4c4f6e921bcd9792609f20cb2b36c27b8ee6e3c6036498158aef0ff9a7a156fc167e1bf21d3229b9852feb12770e290c66ac5169fc4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dcac435c7fb7768e087572e9f531ddd82d29f9e5f5fd7b33ccca7284cab0fcf0b915ab94a55a911a723e385c0d71c66804f3f7f358d91c74ed1ddf73bb8a03b72f37da1984d8b4871a02393b79203d23c734a22d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cefa44df580a178dd0c6f8cef95a2ebe6c4eb835b1f7e2d10de86ae0e0b6f060c9297f8f9a236e988f1e80e392400aa54839189574788e2d64dbdc5c2a37ba0f9d07bac9451010319fe8bb2b8d75a785790f9964;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbef3a97391ccd5abfc42c747780601b2319ff630963326990129bdc12d84b0624e2aaaa79a69efa35974fa8eeba89b3f6129f205874a97f552255eced3e6e54d9de39190a7caa34d87c13a788fd9960b29e8621f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b3b6135b94861a595dd563ad1db075c9f85ef1dc5725881e1cb42010281816c9de03ede2335ec0b9ede2f536c8b992c006d5ff311c70f8bc2ecc67fd75ceee980042f88e53b8ae2c623cf3a730f145546c8da518;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf78a51bc27a01cb0c7033c73d74646ec2320ed7117fa6664d4bb41eb097cded44e38e7113da726953755bec04f5cc1a6d5f68c246b7c42e293ae06faa6ecb369c7d2119efbdc98d9fa498b353f0f8289488895baf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88104f6689411f0b4ab9fe792440fe27d8af347088f81cdd9b530ff6171276b6193f052bf99eb2eb59465ca186965a98dc22c1cd6c81a309ea0a0acefd267979a75b0069fff2ca357ef715882da4ae8e3de0bb2f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b43783ca2edfcfc9b2452889b5bd4b386de897ef7ec8eca78d74c0c8b3fb36ef9783a26ecc29794b862dea0810b4b182b7667f8df6d5a668467ff97c36ffe903d503055f2155fd6d28936c4d28efbe6d534cdb06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed05b52a1478270213e7e00c19d8e5cd49c6c4899fe8f8bb1b1b86fff0766afc47287a6c2d1241e5d3311a91a74187e80b459018fd4d3f52956456c5f78afd9be44a282a8d15db021f141dbd40a9909db46050487;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf6f2643109aa4f6de5bf89060f6e2da00f79963a65aa59754d1d60107fd41321daeecdf1eb0193e74b39d5f193043eabe69f813cb93f59abcca2afb07951a805159e73b563ea704c52139522d94ff8d6d1877146;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4371059649c0895d9ee236a376c01c37dd9ea5e2818fe3361e28e11d15cc63b345afa0befd8d926b7b138057b5806b9d8689c37c0d1d39f6b90af8d9706740c788500ccc99365d2da80632799ee75867c14f28e26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfc8debf4c4d3506f5f01dbbd25b7d8e4c97e223167c732993ba2b06a91d52e9969e8554fc8f2e73a812ec5103873149b2a730338efb8b6bfdd6362cbfed0d41f7b85090fc83a3e36c0f9714eb3494211826352a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55d4f0817b9d8b2d9c804f12591aa3d9e7930c3b0c39ef350f42b449d0e1d357ccb3665535284efc6785fe74551accb6170f9dcbf65ca435b3745b6992896e968a22d0cfdd0324cb6a65ea143cce48ea7b353f18a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h928efab1927949f00926e0d74b2f409e93b8ba4d76a4d688396be26195abb48bf2c0fe5ca6e48651c3698c2f191f43de591cfebfb3ec962e320984184f7913867345c8b19071b8e1c32619cfa94f42b5a5a383b85;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h424a540ebaa67659c35285ff331110da7f7c33b7a7bf1b99956510f44b5ad571638ed16c19479fa045648741abd01a2c9c399c049c5d37b31c6002c2b6fe03ba4461c4431dc72bc091c7a3f613fb2dfaa7f817840;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he23ed6b663e0e7af6b294a2839279c55e3f0c3fdabe1cbbc26f8a6492964ff1a798c2e8f5df3cbd7da038f807e6a4eb55404a5be0d4b29768a504574f2ade2bd319514914e859cc111b68a0354e2e6b6b6ac29bce;
        #1
        $finish();
    end
endmodule
