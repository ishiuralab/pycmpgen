module testbench();
    reg [27:0] src0;
    reg [27:0] src1;
    reg [27:0] src2;
    reg [27:0] src3;
    reg [27:0] src4;
    reg [27:0] src5;
    reg [27:0] src6;
    reg [27:0] src7;
    reg [27:0] src8;
    reg [27:0] src9;
    reg [27:0] src10;
    reg [27:0] src11;
    reg [27:0] src12;
    reg [27:0] src13;
    reg [27:0] src14;
    reg [27:0] src15;
    reg [27:0] src16;
    reg [27:0] src17;
    reg [27:0] src18;
    reg [27:0] src19;
    reg [27:0] src20;
    reg [27:0] src21;
    reg [27:0] src22;
    reg [27:0] src23;
    reg [27:0] src24;
    reg [27:0] src25;
    reg [27:0] src26;
    reg [27:0] src27;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [32:0] srcsum;
    wire [32:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he560a81010755d75e38e90a5a599558e149ef87cdcdbb323a8bdc9a25ef7768a217f7e36b1c0980ac529520000571ed063e516d78943f3674c166d75f953c3cc7756c0a56eea13357f019fa9872be260617807f6d1966dd472af3bb3a15c905093f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4f7d90e137aba3d731d972cc186b1566c82e11d0f4ccf6ee34f7018acef86dccf96c4cf5d73e8e87048da74c1fbdababcd4d8a3377ba054be0c54207aa49e00008153804331e3e835b7f4bdafb609cced6afac549796e627568e555188485de6c92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8248eec1f0ff4bf2d52011f210f1158b2165714d69b23a440d43cb0b1cf3c2d1cb1390643bc523f3ed9a983edbe2c9b2792e43ce13b77b8e4fbd8e5e45e141ae59e0c66779684c11fc5c348f996c8b24290c362b5ebef50c4ba1da91bef1aab8beac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb820450116f321c6007a5b67f35875e4a87b7f20c8230d990b51c0e52ed11f39c7ba8df2f2ae32731061c105981d5f8e88dadaff5c0ce11cdd130f6d7dc7ab140fafa9bd0e1fe66714f84903049091faf5006a144695e95b845c2702526c06c189ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18c847b12dc19fbb7fa63c749601d8d735fdd0244bb512959afc8b4112189990ec2a0a7b6b64ed993788cbb999bc9b157edc97a1bba1f312d2159526f26b66b48b7948b1ad19d8a2da2d4d38c81af160c82dd6c1775c4a4ec2386eec1ecbd528ee06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5395d80c7099d84e5756141b4c02b6927a55d1d6254f6e85b560482009d61902b13fd0690511b3a5cc77ff2327359902e04b05893f6156fc6d2cc40271dde51f9bd030bc59dc63b89d44f4e632e07aaf9e956cae9ef7e3cc414ed54c9b598fe0b743;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d495a504ec348a09ac93850ff65286079e302c64ce3e6580bcd9d4f698bc2dfa41a6140a9e0ac41ba47ab9ccc53fb1bc1b4242a087eeeb09f8659f11d382301b8af52a244eec5b5575a85f711a8790b45851ef5a1973116ecf18f7c49a609260543;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he25f8c2d55b14499abd4a571c7dceb84a56b7a1c0b83ca28db10fe6a1d88c772152129e834e843e578248215d790851b4116df73dbde3ea24016b9be9ba51e1fe9b7e849db44df64791f6c9315af40d07c63333ad1cc29828163faf82abac5c86dd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83800d9ce206b6183b9155858ee33233a4d3330f382330b76370381f3bec57359431f27aabbe56681de79463f301a8909856a8f86432adbfc8dd8ea96cfa8755cfa29f5777b8e795d0712baa02200f69f095b98611768043b674087b28a29b1502f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha60e5a3e3f82acd7b11386339b01fc78ef802ce31c9e1d6105d8666bf158b5379b39418cd63cf1b4185b67f2b18bfb141d144881e90ed4a103bcd662a6e1ae5e29d861f684a0ff5d5f39b25b331939c666cc697d437b923b540a17a204d03d411591;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8fa8095ffd35338588a4981e4850430c4d41baa023e2c54a7417c084ddda0caa33200b3e546ae9008a5c4428fc3905e8207b781aa05fef0e1f4123113f157776fb9c5765d16ed232de43fd416429d3fbe8f5d0bb248d71b131fef19ba2cd79a62f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3316d4b2d0decb74bc5928fd058832ba24eedddde7bca198c202c2d3b128c10c6baaba57a658d9b7e9f87c07e0939bf03488e5d13090c098a42d30313538047a0ebd39160cf90694f3beeec7f097a1ed9232a2447c7df613c792bb69c7d934513add;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda7dd7e315e9334cd8902b2eed2f308489a2c1d129106bee014a999d5f5d459df2b1c0003410e269c34641c65acbdb9804b5f358c02430c7b31b66bc1ccb00114c2938416f03d286d9cce305dfd418e631f33dd77d7d7ae9f8e47854105896834614;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dc464752935d914bb461e629adf79a6a221d33459a4d2dfcaddea692887537d7d0588a415a65e34cb62691baddd6375222db442810f5c14ca959451608160eb0687ce9c2129587f211729d24b070165c2f21939b8831704aa301fc9e2bdc04ba555;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51aeb32735f15322c9287c97a8bc63114df71b28f81bbbc648421de526b2e921625bd321245680870b05c44e26cdf0dc7527548655281cd5d81beee1de03b65a5797c4a670ff4a6b5b001adf0236aa70211f1f5d6f16d2bcede5429043b91f4c7be5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72acf4e3441765efce05daf78e13033a41cf73138b73cbd551ec11766045d23457ca9e3eb3456a63fc5945531f90f48fb0498f17c20088e13b2443db82b684235668c69683ddfd18202db41543a2cf620ff3661938ebe0551afad3361c470bea0010;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfca01edfa1716e0e54e351b786bae24ac7e0697fdc8d4bb8a0b46ac7dadf69a73b54a930115a983b410f85871eadf82ec420bd9b77f921fac21f33290c9c425977252ab92a4444c44d654e2eadc8c979ac0fafd6f7cf9dacb818af1a3058703a33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8ca4a1a7c7c3125c97955a756234b6905a323f86a52f8f4b9d4bf91ab6df887a53652c6a23e7a65ac45acc5c51fa64fd685c1508a5e9a359fac7a246512977019d7e3164d74386e7da702b71d65140dfbba3b0fb1a36e29f4fe6701a0f46caf5438;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc6d416554a15e0d80f972a030ef88abcaae9baeeab96df6142dfda53f1fa862839e87082d017b4e90306fd8184e918b8788c54a86380377be08ee65acfcdb657cfed7b78f6c38df7dd062b41e5879adc77f37e0c619036d1477638bdb820545ff8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd41dbae3177577c6145d2d993ce858e592ec2719c18ad5dab3c1b71b0dc753e0c17b9c4a6ce6930b9b1e71f3d76a36c7d988954bbee97ceb6f92dfc833c58007e529d683a74caad5a02c804b993af2d6f64e03989de6e22d2b7d1618d1b0c3aeca3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb790faacc500e8ebe23065ee5c48847b03e5d67f614c27c91d0dfa8e3b3df3bcc847d93440e6a1645605de7b2e1e61e101e25872c02b23dde91b09000ff9081025e699a97de3a420c1a8973b729a5a4ecb6082e35b9ef450f2611c8af2a4fffe5759;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c7c3167b8fd325280c93e9984c2488e00a8ca66dca142b23039db142157bee02fb2a21bea5c70890fc77e01b800137c7d3e3f6faa08aeae23bc5db2fab6787c91d6f4bdde7366af668bf827d2b60e9dd76ae56e7d23f79938a3d2db09f15f72e6e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96f196ec33a81a49c7c00581f2bca1dccd476a39679da16a3e54dc29d4f1b0714dc4b3b558334a096b73086d49ce07b930ea6c069b5b08326e7a4c87f3cbca42960511189a41a277a64516fe28867c5cb832f7505d23cc859dcd3791097da74d14b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc59ee0715d46b574ed4e279178dab77b402492f05bc54b432c27b13b7619da71d05770a5fd0e0e20b5da3f2bcf6fe9799430ecc7d0bc3dd11ad49c670b48885c92ef04cc4fe088f683f4789237afa4cb5e79cc0d6acbd0f6fc79e868769f2367c670;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc9debf97931915b8e665922afdc6f7ed01cdea83e93051be50f3180e2f031c623d2f1b02e7c08b567fd437e241376e0bcf6f6f4166a15c30afff513e69bf02d24ef72392f87b05bc5e58a94b26a2ca296735a451bf64419d6c64ba96abc06015cb1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha523f7746ab7323b3b5b4e9e73d5d3694086ea4740cacc1b42951002ad18b5c7ec6ea4ba86110f849f76a17b237b6d3442d636aa702e7f525de4ebe132a0993976d70bfe87d4617912c9b32972ea8b4cf2cfa44dc8477781b0f398381bd8f6ed90d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbe2ff45f58c5c1940c82b32ad4ff28e48cab859c015a1505604b89265b35f7add47280a71a4c13262a3a4fd2ff9450667323426a30781dea3351b6e2e647e7435a68d2b3d1b762fc8c02c64f85646bfd58928bb06e60b6e9f1fc4cae1ece8eecfd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f632088dc43af9dc1a3978d71cf4220a1030c044903e0bf4d715d22a94dcb45b7de464dc15870cdbe9a63437496ac2af770292ceefc52dd4846368c0424f072150fbe0d419641144dd58d0b9e262ae92e8285b51167bab00ee4c6ccf74aa72537f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22d9c24088b5c0137b8f030caaddf055680d0c7727f921253e36355d7a6cc3d5566a23e47572e18d8eafdaf837f5b898aadb1709454831522848fb13e53bf44a31237a801ff89df55cd6659acf08512009e56c337d6ff982a5adc8dbd4e2a524edde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h385e0c00dda7654bdb7b6b750a1078316b5b47a907a2b51b36b16be0ed4b450657eea6c7e588942a20de5b00bb55350fa8c6f2d2f8da580870edb40dd758b319b063360648ab6c84437a7ce1a91ff1987e580c107fb77225cad24af24b6cd4939aa0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha52d03a9d49c96577e1768979d168cbf00ad0c274a7b62c9e5dd2787d86a0200203c419c7216b2c2078969ef59df4ff5f727469461364b54ac54ee9a1959775400e19b070d1418fe77c66a8c973dcb8c86ca8eb3fddffaa34315dd633824df49156c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b69ed168fbe2b011b672497a37b10309dd74811e258b40bf0f90811b92f10dbe469946efb5b2163533f8dc6f45307787701829c10a91a6b128d54d13dfa64f3cd5a833a027f6206828153cc1c34a3a254f0f3cc04a076d431bd4d907982fcb770ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha84b34758364d6a06129cbeefb9810726cdb22173c22aacfdb913ad6eea5cdeb7a92ef5cd7472d4d06d5d638e2cdeadcd4c1c80b4c0c99b25fc72de6a1596db939033c67ac10143d555f8009df05eb2ba07cbc24dbf1153df1f8d90d69b10fc2f13a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha129e348285d2180cf02ca5f197db26b3663c86f8bec6953f4219c6cd73a3e05dd6bb4309b90efecd9d11a7f092666b739b6834e4b10597fd0349becd35abb74c572ec19ff0451953cab6858690049084781ca9438393a1659fc7fbeaf93c73e088f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82dcc01362701e395002783e0d27b90063265aedeb85ed33bdf72c5981c0fe500dc5bb4a68d3f33b6955fc6f61b8421085e076130eb07cb3cd6e221f987b11785264bb297c0df59abe9497e800837b83a4f8e55c4a5d4433a7a69c156e13042c3883;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h101e73027406bbce06a40d6a9b14f000717d98a4ff1310809ec7098f224544b39b216be53662aa75f1288fb4c7087b10d82dde3a56f3cb96bc750e0a93224b9db85de2da73b4042d698e9d1fa9e0092e41b77014ece19fe2ef8a9d279675eed2da55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha87ab91ca905b4efb1b1021716a8957e67f1ee5dfdbc18ef9efdc73c9a8d255b69243fec340cc76f870469b53bf3af114a7887185010ac2896f749a470a657d95865f9bfbb652070ff734223222bbae741e8e6181ee5066552ff3c8acb66b0d3d2b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb451dbae5d9bae8c596d4919a37189d2f36f7cb9ea228623036ecf47d971ef69ca30dcbe0af4c4c4711f602ec5ea90a9fa64a5062b5d807167b8c05839008d602acacb3bf76e365150650cec02dafe361cd8ac130ba31fe4aa24e9c6822c87afc4bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb04108a12a340111e8db2c8aaf1e46946757a4331c09d13b0c5a40fd7dcaee7ee9500362d39e079ed0c11b455a127d7c60a7760dbf8b7213bb83f243ae6464a367f50f8db9eea75c21b201b0b175e1781297b9e23c928cfb5b3a64a1375b0dd072c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b767102405bb383179c45566e2a73ade27cc0e0ec2afdab9f266ecd360daafdf50eabb8e51533049069729c7b06fe14fab83f453700ed08b40dbbf0977bf4926dfcdd3c01530a35abff789f02604d9a6320cefa850a773e6633075b7444ef18158a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee14139bb19386f3e46197e9cee8d1ff1c70b292b0900ccf165d124117a0e1d8c979af5de03108ba315ba415a003e7c3044716f0efd25c164cbc4f4f2801b1417e090cbb16c61676e177484a59357af033f3ac980dc9da74107375370d223ba1e636;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6991a78adb5d584b1c8a4842602539491ddf12904d123139e5a13071c10f0646ae90c50492e201727d55a4ef06cb0a88495bb02282bd7914b02394f89f050309ef0bdf56a67e8346a6842f12b929df48d0c7b67fc7397340b2d35cafbf0721448f37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1eecd3bf71cf3f7dfb69545ab319300852278df0e02a61a071c5a3c74ff825f4b3bcad293d6522d415bcca9a4c80bc63470f0d012227f5feadade0bcd4ac34786960f862f0d9dbdb01450d290f895bb828d2529978b4b8075bd2da3c7bed9766d93;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bbdf5e97fd3b3559f8fa6a71e4868571adc120a30ac00007ecadd03a4983f163204522af32fd4dfb6a2d6242ae226914f2c4da2060601c26ade3949de97112a367092f2bfc62f2a445cffdfa7279be895bf54948f4e882d5c567be11c64475ac8ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4b99ac75fa41f08e4e8478c282f9164f17920edc97424240cffbcc46fa2d16bb384bb1fbefd10d385075590497e44e8aa9f406ab176f743257427cb60981ecb9379819e8d73aa772c0afa022b5d050a264cf74f2c96d6d75d4e8666e5acb074cdee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b7b658fdac3ab1e597c3d2460814ea67ab1ebc95b235c37d29ec5646586aaf9b36487a7a4181e6ee83157173201a53704a1d3e84bbe5194d73f113b9cac67409a1535ffd8d5398a6c7f6721c5691c32641d615a9f17408112f38204f0f797bbd009;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46b1c35408aed8879c2b6b3b7141cf993e80b9614778e2e8edbdab0fcc55652a7801950604420161d5f89bad14b4c77ec6f30a11f184c4f7a589a68d00c239d6b59fe8ea7da2f75d5302e92b0946dc20a013f52e0e6beec87471ed04e6b0dc7b4dd2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h110b6ccf0cbabaf2e328054c3f53cf7a3744a9b68125df9579eac630037d9625150120e13e9b2f0634fd65efb06cf115fb4277e8291a3056d0e94dcf5451830916e5dc83eefcdce1ede483a20fed1e82dcd554cc47a67d3ca45a124101fce4413c34;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec3f9690459b3e4fb7e34a1fcfa7f58f255eb302180d0bfc976884ca1f4575118f5490a90bf761c3b5e930ceec134f382c4af52146538df88b5521f1d9d84f93bb2bf64aa038c763e7c91ad8de6e2097f84e57c5487ef5aa792ea7318fc7c0777d5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcff4a093345b214536f66cbd5e155a254ff83755dd441b247a695a69d0c9bb171781def50fc82adb5a026f4a13a2db2082bf563d2888792d8540216b4e39bbea8c17979e89204f077d4708fa860e68cd70a26da3b50a30b045fb64147a5c9baf3477;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13e8c747ae8195c798962c23d24c620f2af377d104effd716935b2d3d9296c9dee9ef92d8a0ac346fd39f2177337586712474f3bf6b23f534f7382a28939ad21904767bbc62f0e0e8b959e884436c275fccfec57cb29c075b26fb5388974dda147cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h114ebf5f118d76a1b256cbe7ef12c72c813175190dab316b9b6f132bef6a8baf9737578dc507a2d533251c51c63a53be6dcaa66f42f682ebe7b74072b0f9e3fa2c67c4b6fc535108337ed1b44908b3af69ffcdf1c10de2b57b6e9984b1e12329a241;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52d62e15c910454132aa3a47c8b8a4bfc6919fbbb2f8b33537ae43ee768f8f1cdf60cb745fb5017cd0bd53a0467300650fe3716b1d91e16c1669886d0ce274b967db784a59463744029e8fe7baf6cb7d71ba1e9aa50d43e96cd4c96c324d65f20e57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd78ae6399b9d5d2b69f4745d8a5d78f952509f310262d651d84952050118c9c7133da29588e88732861c68ac20093f58f48f749becb39c7c118d027b894308bb8fb4047d1c40092a0918834f42eeaa6a4b4748e6dfec3d8fe1229cd1bd8b94b23d18;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb411126b3eee7b3f63aa0d342575463fec4a8ee93ad9be50ebe8f70fa0ece1285b339548001add3b8aa6ff23dfb78588b1c847f831a58b364e69b0b192601801f340677550895e9f97d579d39f602c8d20c081e43046a5bab0c3031ed488fac2cd28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b2d737f60cf6957581be6825ce6ea203485542823276e81ab74bbe9892c012cc246df9d10f04fd98c410ab7dd438e2632ed84e2ffdc45d6fc77e8a3b6deaa9b6b2ee4aa76d5072cd804dfc0d6f1f607fdb83ed686aea464715eca57c33262ab35a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h606f5816329e9cf31dfc0675682295a9ffa43b95457c3a9f10de4932fee56cda14f2b61dc076d080e5a056f835613053ac8c7b6ef569e648fe4a71011894a13c421be04d59b096f77e4a3529b7d1eeaff153e473a70fc1a940130ab7d5c6b5665fca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6793574afcbddb02a2ff41e683bea15ce12e46da2561809b18d826d05d68df86b3f2a30a1a8144670c27daa5e64f3f51fe0209dae82c77fd350e7f5cf0e535860a44f95b4435001c49295121f9d3944752910aad86c48b85bef8a918b9b81cab695;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e7c534b71c841f6d146dfd2499d9c47b4bc6931d3e4b302ee26473c06caa5e6cc54bab1598dfad9e2aa5c4be5e08a1f5740f7950704e95f5f435fc4a136415131e3535a349f9d7d2d0d652faf17e7ccd4ab1b876018b0135245c1638a2893ea7749;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66adba1814344d267230d752e5ce8967cf4877fc2928b9d70543d53769901627a91aca710b3c049a6f532d5f5fca2cc4bf73f367cca2ff22558dfb4d9a0cecc4d739301b82cbadccba920d378954d21678eec1cd724ae541db6014a6d39acb0e40a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0c297ac7b6224ac89409d7e31d3a4bd4e248aa87620775b3406e531ff568167a06f2a5b1bd3565c064f8571df1264028af8118dbb108c46ec54c42286fc59ec372aff367a08be1c6ce6bf894d776c1f2cf073ce071fa7dc7581b600c2071531bb8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h211aeaf1058c06997a115b5aecdab571890ae07c95d816b76fc84667e2867a7540a5ad19ace9be2c4d13b20dd086326383b81292e2b17868ef89f7506884e06efc39c4644a907a4e2425d70dbf4139fb828cbd36237ecd431064db1075d6c5a69eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h741ae5334cf4093a6f7dfb02f7dc305f326d9f5fea4aa8b4d034f5027ef15c3ee99a6a37d096545fc23c7a238e77ec92ed18f84f94e67710618c0007fc788b4f42c355ec8e583e68547207718f853c6baf1b7a0a75d29014246230f30395b7f04656;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he11c26aa356ce2e440d2a962ad70a11695e0553da78fc13b4c25ba502e75012a786f0c0780756d53b7fd3495896d3ae2e1a79766993ebdb671d7b7565c5bf42001ac154a14bab0f5fd296256c846ca294679fce072daa756eabf5ce44929076ceb6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdcfa853553d11f3f4d7087a91c4e2e60b85b4e23390b03cdce1be91b793f7280a81b842ffe1ff1afec8364125bb1b68c31f4d70c3c8384f0ce7823381ddd7d7d9e978a8028cbd18f8abb1745585e987f3b3d9014b34d41057ad8d15eba233fa6154;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff24e77bbaf1768609f58b400b47af683cbe6e819345e1ae5ca1030745d1a1970a3fe6d652399fd85310bee7ebf86ce63780a8a3fbdcdc947901382e9044d09074558469247f7d9fca15502ddcb88c7280557a64693efb478d895785834201008c24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2ef702f0ffd660631d1057f9d25939574c233b833ecc658463788213054e38c7c9f67335f24e62b275f26e638882ef84a00e1bba0bb6454efad9d1c911f7a50d82e44d9542db31ec7f536164afb784b506e7a26a5e39c79f13dce60db205d86f786;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f61ee5f06291b7b0ceb063ba08ffc7ae407063c38ca6de231fc56a6db8fc509ce78e5f0f656613a3eb307cb38de77b2985052819c31ffca1ee2834bb4b2d870ae8c3d7b8cdde1447b03d6ba3983fd8cc869d56a89fcca9c740854a3f9881ffd173a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h263013d0598002cb3f8c9ea60e28e8c7111e01b501a3fd49945ebc0fa101fc8cbd325f98387d20728439fbf63624a46586a5088c755432d0819cb01aa740cd46612a798b77f1c44c6bcda0f7e7a899bf41884698088843c79cb987c46606ee59e289;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57cccf76c29aa02bf21ffab219ea95d4fe8c3ca6b449e88672b46486f27a0a3d6743beb66ca1a7e3d500fb58bda9e966fce1fccbb9b7809a41372607c6aa1ba01824e2020b1fff215de51b5ebafacc67451a79a84753c15d7f3b675e322519716968;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h718838c91a120be33ddf860d29a68368a81d84dc401f75bff6c3f829db3e2bcb7880a6ddaac17c2979648aff8dda8c98fc5b52bd6518406a084a814ef0e5f330fccd295e11ac979119552ec05b9c619c8af53750c9f74b2ba61c61c21e8fd8bf6078;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79f4964dea9a87e0f8b55467beb865b171fb12fb939331aa7beff044db49b60fd4dfc6f74a7794b412427764cab463cfbdd9c6cf6a05b466864bd11661591e3af03f421147ddba288591405147d7e9b7189ca3b7706013d8aa3e0272d8d95d1750d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7023720b00387156b965222ec28ee5ecac036770da8cd558aeb212c03d10a289496e72d4e383cd7d99cdae91d8a50a1445eda90e879f4a641709e969cdd71e7f123e6e12474f008716b5409a5a9b3229744ff3c1d827b3dea34d3bb6178ea8fb3bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee765f2ed41200155dd6d25b12beff0207930eefa500cb3244043bd9111c432a337aba066a09ec82e034edac52a6d2c775c90b922313fe21953c5131d89a731929cf0172beda97d4c2bdb9ae0eb0c543ee05b74359d2536c0f85079525fcf02407ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb13047a9c91cab1bbc0fe1dd70ec062ce0b82a4f4f5068aaaaf010429a70f56fd856c718e8116d12959ce7002a77894ca3f3c0ade074bfa7e8063e122156033522f83a7ea7efd8e3b3cc31c770a81fa4084cab0ab81b4f9731e7207971990aee9f08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he819eef39a63fa2a74cf65adb77cf84de59db0131a25c8b606578c8fd518ba06d6342b7bb51942df026a4cb7fb8efe6b442c4ae63aa39fa488548496e6954e261b88a7c6ca167f3ea7d21474fe5d1a43a731cc8f346fe90b2a1b0cb3613b34bf443d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2e2f10c49f0ed158df6cc072957c9c59b6054b5120e50d3e6fdb7c3716ddcaea6f37b731f53eea765f99e5dd3dfceaf06dc3255cef43ab00dd8e9138a9fb5f6ece0487561d870627bf5d04468c03baa8ab3bd84e68c1558e49488dc4cf8faf4a5bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4769327558e9772d1d4127218eaec7d5b73fbefe094d50aac0169aa6361dd287e7a7cd2b33ebb70272f5f66ad02fefa010a6599fe89686a9d453726babbe26890034221cab3f1dd6d3c55727b1020b3f005e5f3675503ee0ea3a78f9e636df233b72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446514b42046727c0cebc988c89ac9936e12876a5067c982e37bd6f3f123d545ad9752c80778e756b1401532b6edf0be25bf163400fc525743a9ecda84eb8be728b82069a883657720a9395433dfbfd36483e132e6376988072c617b6d40385c1ce4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82c7a5174d4746daba934f6e04c847acf0f0d7de1171181aaa29e57a0cd1a15c9c53c5aa45e755b051e40c4065374981f2bee87989762e3f4ed1720bf3069318cb87d8d68259722ff2f70bafc3ea74e5e1302f6517f1c60dc2af731893b95072863d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5f64a6f873d450a28262585c232d313ca6729bcc1e594d79bbc2113611f1d88e51afe3776b438b3c860180e15595bb2a7a389be46e1f17de654150353a6d6b52507df16844413d7e599ffed13a09e745527d9a57161a2c8a125b1f5c3197f519a5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4824f22e6403ba2b92f5102b8ba20ba047189dba37bb89a065062ed3b8bec6b1586dd889a6e9e2d99e1122f65453a0ae1c9a7ed7db277d9fd71bba030d47ab1f062e91c46548514d1786b502bb19273e838f86545cf73ee991276b66f1be3fc8a530;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84f300be1c5d8130417e95cc3b709f7373cfc5e25b7abf9bc55679fac140833ea78f81a98bb6f51ae3b00d49d2874fc8d8c7b46691baf68ff5f8ae73ab737be5a367872278ae1d6391e5d72128a0d140104cee57d1fe91e1c5078068e1a168b1da20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h422f2977efb9c375c5f381f82cfe6bea121536c25a4f7e0bed5c48312007ade64d0f8875c7a0df965687b497a9599b3c18f8d7113a845dcc0f90e8903db676d646d42e06fe4675d1331cc408b5de08ae48c9a3e12770d5e7df59d44db910e0888656;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3a720be273daa200020efc10194190df89103532d21b0ccf27d2bafc72ed78deda8ed7de81e62c377d6c4180386e3d2b9c8fc6d962c07a8b966bd97668e15215c224e79d467b6c12decf4fa2a2f65c18141ac60c703b187a1b46f20c5a8aca65a32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47b7550b5afad22acd21141b12c0d85058e2df5fa3e2c69174bb5a352fff8ad6b008b5c5d22eb007b6a786b603ff3047388a369729c3a1e7fe5b4bd7de715eb51533adf4d15790fa79212fc069f1c66f2083848233c2195848c0c00c6b9e595ffb55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h562195d8718da240b96e1ae2bdb8f04c01b6d111e70547f2872701cdbc4e582952e84320c2121d48d62a7862d20272fa523d5d17c61920e6d616caf6abbdcc8de39a16faf8e6567348a574007a4e8e0869220e5fd78f57815d43326f5e076a4d87d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2dd3010d3ab6188446195ca5fa1919db4657cffa0ae4b5c5643910c471d683e2cf55d16b0426d451f6fcedccc139a4244516b50830c43b678c080b92707fdcbd1194c0a8f0fc79641da30a0e18286c27400287c11fa4209039a12da9a9eb0b38555;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69e0d286b4d7af0ad3ceb79f60dcbfd5db3b2523f23bf3b81506ebda70fcf5de32f7b83dd549b40a2cdc454b85f59e1e2bb514db4c2f3e3b69a1eed078ee1e7f440e008679cf47b16091b02c3cf8c74c30345430a73f98b192e028c56676916be69a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc755a3f44e8464c6f53e2a3ef86e49fbed6717603f4e54d8c43be4c8ff4bb71f5c934b3f60fa2ad0f65bc3cace9c9bc549e41136a0d23c8b57a6b77dbcb9347fcf9ae4f38ac4c77974c5aba316e66d67a60edd4e801684905bb9086181c6c74982c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he32fb0443ec50448396ad2660b01f311f064e0fe4167e810d07b8718304584629d9c59b604ed30c06c302ff990cf670272251a668dd012c59360fc52b34afe8a886e5b3455c68cea04d08346fe019dc0ab28eb5e6e0f394590f4a511798a54953b3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h188fb3ebe68129adbdfd5817ea6a95af455f6214817f0679c9fc69c388895e30bff7d3be58ccbf493143317b97789170255f2bc4e98bc87f830502b58f24f6180bb0e38f38c57728f921667cada3763f8968e122d0ce1c34662fe074557ea2ce8f4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7068424027f7d2015e252cd9f46cc89f9495eb1d7642182ec685728c444769f35195f72193fd3f19ddc4bec8049f6b6f432de702ddc4d8387ebcefacc98179b9736b190cf2ae0dd73c9c439dfb47beb6176a051f94f6a743c02d0e1eb8d3e96b2ffb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5ea52f6b8801c4e11770b632d7db9fc460df2dcccdee4b830076901064ae5301b798612d6bb2a4856c485b4f7273abe72c5d5eefc3fd0cfad9fecdb98112625e405ba36afc6672e3fe4379086b698221d5abcbe296e364b3f9e35efb7bad368c41a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf96f4f34057a3612654b0ab208b1e818294ade44c8ebeb68536acc1a79809f6287dc04f4e40ec5b61580c6e0b1638fd249baeacf38e9ae2088a11d2cee044831f0cce6424b89d6636ba80135c17578649e5c34c747373e2cf96877d44545b0f3e09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbfdb9a7ad86a203bb999fca9a83386e836bb2846e34d876d7f7f60934f6f6a0e45050b70953918194eb00a41dcd77e2cdf8c27e3290f96e451fdc7144cc3fe2503b4cde05a013f35bee1a10436ee71dad3f51943561568adfa4dfcb885f9f3111a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1e77dee8cf99120db52e1c7945a47ee5a3ce4a29aaa8e26d63bfa55a79c82c168f83da51214018cbb906bb69dee9632ef6d154dca6eaed36e5cd2e6a82b32fa2b854fe47de1943e088d98cc170623c745995c9d63ecb42b1c05cb5d1e85c0f8fa0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd697a5e1bc09588c835e3d2cdee60105990eb2b0f1af45b0c7f6cafe1d916fb44e9cb26a40f76a53bb92a394351e0f20e35c71e7eebb3b4f329e28a33a8b1b6858079d146cc55f747b76192bffa0b7b2221436c9ce2b2eca06de5cc7400be6d63d06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h533d5aab0bf2f5b685045f20b5f3776117844f1992c0bcbf33551b82814a1a55f500e61862ee99e5c7ca7f3a74d775eb184352f12603a903a644f58de56c70ec2461caa15f9973df62a2f24a74891aa44816231b371a36737baae771ed206a6a19ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fe4e2246d632cb2a434db9410cebc014b6eafd7c21757b44e5f1ba7853311540713f6841c0ee0c1884982dfaf77a3ebac63ad099a5d07155e295632c7add3775d37e8cae35249b237ba980764cb961828734a92b336184a5af034a12e384392f3db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3502590dcea8c5094ddd4351e876fe9225657c6d6be7b36bcf9dcc42449e6ad4dd469516725dd03395ff6cd65ffad28a3d673646ce2fc7c7043de21712f66f2588e041ed567237fe072e796d854b5524fc4fee3a86b724cb974a17d898995165bb41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5568479476c4c9d1e84d14214f0c91f42e709657f37df2178ae01a555077104367839e44b145b2ce8e65a4c223e97d012d80d96117b56590e4a915c43fea576accb480be0f2fa80f8cc7d4a2a08e436fb36bdfaec04cde3279ca3599a4cf058c1f49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafb5818e7cd701b3f5707f60fe256169e62084c117770d87e34314eb92137a629b67a644a8b8e0e4467c0da0092394505d2ab63ba4e68123300a2d389b4991a5e0db130f0d5963c05eb819e360b65aa186e9df80674d3016934fe65aa0f7a1a05603;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68c6b01926ddedab80cf5363a1fc630ddd698ce3f6e8ba33e75a3743e7917773c7423c884f1165ed53fe14dab31f5b274ec96aebb3295353e78949d5b9b34b38c46655679a5ac97411a3422c2aaae9251501bf44c487c073eb38de0f8282613b0772;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb598c280224b67532e86960dcc2a1a70fdb9ae6f6a744817c9722b553c63d0c6f1fa61dbe8ca707bf34a9ebc3d846601bb04a17e09d54b17574aca91b143c1d7f03de513f6e25a249dddd71f1e54380f0a026387ecfb0d506c52119660d0abd94a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f96a294c2fe238f9ad5da60d5ed24137c25ef9017639f51fed1ef3212ef2dac7e564c576d7efba8c667e45ef1f226ff6c3a2c6d7a8b472b2da2a591375718a570a513e42d57597b8f232984568b113ab5cc6ab55381594dcd8dfb6dd1907b300e80;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5095183eae4a23afd4a44347da39f990f0b1c18668af86e0380a149180648206fd9d09f1d2663e79d6226c9ea58cc986a3c274874537b92ef1ea6e710c8f4786a88fc5d684afdc3c12b1b1c3900d6512d88d6d0a70c82206f10fc6ce58e3669049b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b03924520e2d721821c50ed26e2765076e0e3362f86bceaa17a3b1eb570dde847a8afa70a7a82b23e543c55db8892812eb0a0bf78fef9d080a83856a7c682f66ca51a8024791e0cd8f0a27638de1b6e50bd1a46ecdb8a3a837af13343d233cb470;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3f1ae08b3b9e7a7a77e530e69fa4c6635affa2d6b9f4f33412cd01cb0383fd37932f80f40fa620414d667706b7028fad59a47acaf898ef7d74e17abde1f4ca1443450eb4e97eda0301ce83ab434ae72b67a11d72eafba34b79546854321a1248393;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0ff96ddd84ca9fd9ebaffa3e2932f87d7cb7d97cfc9a5c00bb90d60233534a572bdc44e60586ad8be39114d91a0ecfcbf4c803d0a5dac8348898ac76a6063d84cf9d31750ddf9563ff4be91eb028ad178732ddfddb966e944422166caaa2c7c142a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf0ae710be1c546eaff5bd884243d307e8852e965e1759680deae3b1d530a099a3a5ad6a85b7e2c2eb97b9aa62697ebd6f8900feed123326cf0c64383cccf24776fb2ed54ddb11f5e77b976f41e6068629d46e122fba4e21f5bd47216b7a3b9a8275;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha26b5b3f966d4ed3cc74291b67ef2a9beb9f582f648418482888bbd9bae63899b70b1ac8bef0f97f02695bb8b83398a5edb8f997d3f5b909504da2fcbc3110a6f077d92fa550317ebf9e2a6eb57c0d22f8808fc91f4256581c616888444e909d946e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9351c83789de5ec0056b454a1db4a366226cef536fefc77672ad03d7c26e6a7a45beb13458cfefacb0d6ea31313aa5a9eff90713dc0a0b4f5b11189f00de6f45f59e7738bda7c022728b704907ee5d05afa0e5a1538955b5b6cbf4c0c6a760cf7d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c9d9ffc105c5360ec568afe625ecdf35b1e7fc467be1616b9a923140b53ec82f25700c2f1d5f0a6ff4eb89425f5e192a88c591679936a0891688759b75c63191fbad9900c12f271f8fdc118332933d752c056699d50c8db40d3e38c08e079f0d209;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9d0bf40199e7317018f87617b29f45a0b828c670fb21a6ce073fde2c0828f0a686163f6944da6529ff3702d029441ce8dd050b89e1741c0a9b088693961c21d29b8039f431a854ab4190d81f3623bcbc8c981f1a778939e70ebb7ccc195d2c74e69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6dc2e14f5287c9e25d5c97be0d0df00eab57eb41cededc81b4632dcfb626f7e89a17432312b35c9f83e05d5b54f547a32a771525b3fdca16e072dbb2506ff5c0a275641e5b4a64018d9b1cd2cfd229a5cb17d55214b352e0f2bd97d33087f8521a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7d934c6860abfa0ffda22588526ca6e57d839280faf40b714dcbddce175d148a29283439dc2a25da2c582eabb2ef8cbb73646ef8c9b243b621d61a6122c9f39afdc3a362d3f4ce52816311ea6e0a5c223d8a07707c5e5f018fb14b52cb07f2e84f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3045c9f240a5d9efe8112ba01ce68acf7940e0b2eb943f2179125a9a5490b270f16b6ffb70159ccb8000a6db6150a4acc9de8c750e675840ee5539676efaf0607032cc0b7d685a7a8d9a70d987c4b8c37af757e6ecea98077007263ac5ad1fd81ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e1c8d2a26575680a5ea97fc17aa9108b3576a521d4b90ac09584a9a4414f5518a39c4f4c1d615a8f528a820590314301402bb81a2abee1857e5407b5ed52673da56b488e9e7cc9065126ea323662ce24eec2b307d762e24d48195bc63ab7fe9a56c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69cc1afb84cd063ffdff4a4b7fd48e4e01e0f0f7cf3d5b145aff37ca43887046f2fd6c6679d7d18a2b568dcefbf6ca982329e6d55ffc144c3ae72e8594949acae0849c1774de872fa8ff59ef3961790b2ef92a64f00a9c15b0d59290c773b68a5727;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76e348ee2d9330bf6e887bfb29b87ce36c57240b7fcbfabbd015a782f7daa31161e2cc9cf1060d90b6eecb5973a8b83f6a49ca4027caba85fa1507e064856dce9003c48d95bcfd3e0a7184568b0f53be64f046e84f7d483ccd32fc8f5b8405882a6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde5cff356b9586cff4842c89819c9985e13a60e041db688e6f326e78b67b1098eeaf9ad50b7a7e96afc761109e034f476cbfac848e8e7fa9669299850726a061a780671c178930b64e4e8556aff8ddb27fdf2834e56847ac7f5f513b4a47f881bf6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9df0717d9ef5198a999afc50aa53d99caeabb8f8a192320e31b998fa509a9e1eb97e8a4eea23c91bb7bbedbe92f98639f2557fce9eb8cf6474484a7c88d4f0fc1326c243c77328f91e6cd07219b4916eb55d40ace778df648147b39770674f27dee2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc16a5116f4b893a1aeb0325b142499241dbfccdfcfeb4a2ba3b21095265d74dea0a26ce622d9220ad0a6160abc8b5605fe161b2947c844c6f5635a8da5caca1e4c4bbab4317d173a10fcea04ceac0e6fbef4101debce6b4fdb218579cde100b64e16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec7717638500067cee2eb0c8eb41f489b04c36e57c080253d0c8ad7f90e14d9c06fc41fea9188d95b2135f69dbfd5ed221e28febf73931728edace2ec2d9c684e979ff9a2e66b9fc717c86edd99fbf499649d5a2be39736cfb45c30a4bfa9548f08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42f00f4a86140c4f1d43fd2858480d2f31fa9a9b22c81e9f8e110eff1cde8006947a3cc4c6ac5d388ca378a7e417154d5adb2eea55277f121f952bab5cd7a2a04d6e367650a07fafb4b155f6c6d10f6c512019d0de64bf9c774b280825a41a3ce867;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc69823ca7abb04fe4537a26d5a45071eaa7a44fbc8f270ec11c84ed8f0826eeac6c61a88f104b30654776742befbb9b9e11be7491bc750db2cf156edd0c6d56563f9ff7028e8c9463af331367ef608142106cea9c6233a4d01b8982e5c98f32c37b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba29456094550c08c69bfa390982439ef3ce5735cfa37ae93d3a3bc7b567e6dfc2899c6c8d5b5f25909819b706e3dc8ee7e03fc5ec9c230d5400b7a619f46428a62a42e756982666bcc942e9f52f66b3c3412a8a8838f6036215e37b6331e6fdd01e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b47346df2a74ca40c3ced19ec5bcb6d3ccee780163f2a5a6cb64853b7a6e2b8f5d590a8af4f1a5baad31adcaa607b3fa9ce922d56d2bcf92515768aa806f05941f5945b9d77a3c92ef5c767ddc27f278bce62aba0a33ac0991ed569edee0413d9ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e2bfd597a749812f7e5859c1519718ebd3ca8f9c4fd42ab0f82ff0124abd019522f1fe816efea7c61f387bfc059ee5361654f4e6f6119176e93672b83b84b2bcc2d11c32de361dd1274bf4de91521f7fe6906473cd925a510dd5c448a3b8e74be37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1865d3f4c767801a21a0601e30193a51c4611cc9c272c98fa16d741f6177324bf3089edefb9036ee929a6b1b4750fb21a20c84a607ee126a9e84a09595a3deee7d866f2bd531e71d5bc477bd2f2ba1189434d521a24293823b3840c87b755968ac4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8591310604492d0e63196c43d0f15a01acb7d4114abb4af7e3136291025c2232171e798174e1f100a4b733e20ec935a79ce8571da42ec206a4ee351f0a633ebf201e18731541ae4089482c798d04bed0f484392be5ea4d0ea2a3f7615afad88e2178;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2f0429564a5d93dc107acf0c0865546f5311b2651a95b472cb5b0ebb8463ebc9dbd4bdf3e5b0a2b96d8fb662947ab38c04cf81b64816ebdb68a39b250f8596eefbd788b44ae411685c75327560f384df90423f4be31425bc5db4c7abb95700e1f1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h208fbc8cf3e356fce116db6ef0d11e01525c08029cd11765b5c41650756e540d3e12cc008d85132935be3b13e18c63f98d6b3c828bcf1c19c7c8d544bd5509d8b6b081b464da00d032b60dcdcd020e67dfd72d7d787687da2516e514b8312d57f74d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fcab2ae9f8ce60f6f7d4b27980b9299ec31b9379104d70a9920759f13d01b5b2007f5cb8becb79c3d7cdf4281217988d74e0ccfcc4dafcd6c281a649b48fff3614393d9650f3c0fdd7637aab1a3a9a2f04c6f251e8ab8c7522e8538b2da89c99894;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he18ab465eca4789c80964e50b70b6a508101bcf3751b2e1e73b7060548286a87c1cfb402592881c9a7a4cf14aa5ae7710e048e66b68b0133a16079ec664585c083d9c41893a9c9b0dd48c0f250a3ea87d08efd5dfb71dc285f7ab648c6b970bc4625;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h797732c3aa04d474b227421d53b25674068a1993d27c09c150ff74ca329f9dc3e8277f791bad86039c5ffb2ab2dcb116c692725814dcd53267486885adaf0d06fd818bce155bba53ea39b56b89a39c5bbb876f4ff0e4768897d51b3c78fbadc7820f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91884709611c1726b9f5c124d8f24984640f93c258e974058e445bbc252f470b7902b3f5ebee0e4ce2926ad3f15acd0fd47171262800567859b8f2f7561c352c49399446c08faa7a7c6b38c9c8310d6adc7b2a9f937b5538960d4bc5ff66a285c77d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd04b72167b6821577550032adc5cb45033be162a05f14b829ad04fed53fd9f0c93e110fe22369209eaa9eb0146b0a384f58a32141d68059d6b0e4d88ec74f7c2be20a1770565386a2618a9e09858ff062eff03344748a0460f19aa2b5ef3598f239;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9130b8b3d8f934d25ec0d2064d79084d53e57c4962ca45a2b316b983ec3acab3068d0de10ef3efce48c590e77ef238da29d6656eb5299260550a11d2e7668dd6fe6e678e0c0756ec1a67cd297d218e11034ca4fee0cadcbecbf5e0b498c6e67fd45;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75203d200c75c08135eafa5afc76360d1df51ce6882e1c3603e1bce022ba7dbef8fea2d611fe41b2ab88c5d6531f3ff2987ac443dbb4d3de1f75502ecbb641b08d8b560664a07593341bd45c785399f7cd6ae8d7729b0354c7771d936f97e6b6661d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff49bd65c2de5457086f0d62dcb82a13ff069ccca9e5662060152ce3c30ec354b9f3395675388449c59a152f7f9c902be15e0f59731cfc1645b3e6173e42df5eaffa5e93e1dd7c4ce17cdc2ad4e3faa542ac72614726cfd1641fe754236c7227fbde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1568478f7b8d27ee7b2053ccd4f2abe7e3b50374e1cae39bdf7ae3b76c8c08ae2d549b168c08e824dea059d819a6eee18ad277e63d73be1b3ffe9aa2fb1f69b292af010aec283d1e78b33d9698efb4ec9a20c6515cb0c128ce0372f0b1c28bc63348;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha95a498a8beb3f1bb0950eabac8d31470052c094665ff7d552d11c8f1287443f1afd6ac0a29e25750790c3887cda383a158da76783db55212b4109c38219c50c39f3b347a5621ea3b1659189f6b417afc9d6422119a3d7007bab45547afa8af2a65f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d2c72b7ac1c98cd2b69b3a16fa9909487d01d3f3330e1a6a08f34d32d863304ff1dfd0921d9c294998a08cf5bb00c553b85e47a1bad5db3e226d1981668e41eee19fc25fdfad9bbcab589906bb18913d18fcf220cbc815ce4c820a28697e53f84a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ea53d33c9689b877acc30d4897fdadba62f87a1312ed9cf310b0fc482782d0607a44abe5619574416035032ef88d30b30fdb2b25016a9ffed20dda547198854dc1ae487ad40d997aa61f7e76b759c5521ed0ed2edd85eed7f1481349fd4f67e36ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fec06566951f827ed27979b751da695f2774794e51a814ace58f7cee70f8570c2ef0b9168d444cded68907e22349d434dc1a13d0db3dd24281f209f54077f42e47cfcef9b1d7c7234d243507d6237d58b93187cfa30a6fdde41b24aebd56ee5cb31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa5d938d1f62d3988096c7cf33b8c22cee794343130d68552f7261839aaecdaece0f69f2a94a8b06dc4e97455838eca039dec10b5e176385bda5e3922e7a32d623d9c0d639e8edaf440288a22ceebee9dcd9c9aa1d538d10ff83e32133b9e601a905;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7be3dc64b6a62cb857a9e91eb191b6925510c2065c7a8b19796bb36038adea7a3a78ab6e02fac96896222eed6d0df6683a3d46f1694e076d0eee6d6ee2c4a1d2fb817b3c34e78a0bbda1cc115eef0712e912cd8b06e0b29993a4af07c85c16088d20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d33fa98c1377f1ca4f5172489e197955dbea1347077d557de6ceebc0005f1cb25788ed11c42ab642136e2ac2f43f5959458cccdb3552dc61f31b4af524d1342b688b6f1719584aa2b11a3318c7407811dc537592a5780452c4e508d20f7ce8b9947;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32aad856e0b1e72f2394b6ea3339bdc8f28013d26a4733cfebff8e136ccd6c99ebeab899fbac04de4e69cbff0d3095a84ba48571da514e941720fe5a7c9a636a050a873713c6751551fc2ddd0d7d6315102c4e3457b3f5085079642f6ea066e3ec08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1c02927796a7b9642916bff8284c94fc16cd17a81893c9b5dd3087511be608bac30583221ff7317818a0e3f894eedcc095657f9903d21dae0927b0149495a77202782e7fc3bee893b962f54450393fecd704871125ebaa6067eacac3b35a6db970;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78044fbaabf2e11e596e5707c044b8c30ceccd9042f82362ec05dc77005a30e06b09947834db575dda68f9356d7550f242b53b95f0144ab337b8d44f2d113db368cdc77ff3018561514ae220869b2ab6f4b30241bc2ecd326304265df0250552af6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a322c16a0091a531056a4eff2c39afcaf2f72ccca7faf24642713c88b716cd0138b3d6b8077e5a933de8146c91c9a49fbe3df99b39b51727003adf889b3fee7b04182f39f74059159adcff1144b314b20ee648ad30bb1513bb42459b9aeadfbb9f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cc027997b99130cca24a0ec88964c24a05cc40620a28fe9cb98c35d63e3c77653901127e77a09cf4a008aef62fea573bcb1ff360e5a221f8f13a7fc8e90c5259b9cc621a0f1bab9e47d7174e7ddff32649ba09977155f5425ddf8d3e97e2608011b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4dd772c01d3e4938d68b1409cea9b13bb608fb948423e00a3cfc2dec36835224d911619a44d12539afaadbc80ea4d71eb042a32e0fcd3c8374f9f5b2fa1eb1dd9cb88d04fb22cfa1d820236803762d626b1312d74932713f3e4ba4cf82177507513;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf37f1b216a81aa06bff3c2bf520746f0a58b378e1629f2a1f33fa5ee6a7b86393d070cd46e79c2f45ba5aeec1e29b8bcda76cb9ada6362987a93ececd169f9fc45bf679e67b33a9f09a8e86c90f00139e6237d58f67da78152940b5a009adb523732;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6354d11d69f7b3f5defdd392f292299fa0a7bf4edaf361615203a89f3942b97b4289a09a7e0b04738011fe7d8abde3771d53ab6e63e20840f7d3a66bb5d920327c5627ba56f4616ce7064278a7285d8287098a01a8b2e2fe550b29b1f702d84c0f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56be7ad05f65dc5275d3aaef61e9658893549b551ffc756625148c8e56fdd2ab68430f9f48eb0b63dc5f0189af7dd47b26585dc6594e5127d9c18bb56b559b3de721cb470dbecf7befe0c1b2a0accdbccf8a86694d28f23fcbeb6ad7488a3b8d6c10;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f7c29723d33497a40bb3683609be69b03ae83c8cdd5c78601365c9134ffed1bc90ad5f0d289dd0bc1f79620216dd675bf03aeba757aeede7d195bf2d74ce0f7c8d5095b8348cbfd4bfca1e80cc7bfc5a7e8a3448ea4673e16f57333c75bc174110c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb9234b0ae14f1dca1b92539af92da4229f5cb35e922362df4f8e740e9d974139ddcef60c554c166ef2e9b11d384a14fbba65db9760e400dcf3b3a42ca8ec11d729896653202b78d19c81fd0892172d0bca7e3e9941b5f7fc1505fcf47b58c0723d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba96d650474ab00b49cf881b4ed5b091c1d978fd3775181501d543e8c558bc61e5573fee0d3d9b1736355619c4354db273faa91c014360e856ebf31342f706caea7a6b2537d7c9bdd23e5d706bda5b10c638e7138cbeb5de2c94831f46ffca17d930;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fff4ccb3366ade4021f833518fb430555da787cbc68842eb199f5cc8f94be66baeae27270544bfa82c0d285ecd49affb7be102d1b4e8c560717e1474b838f501a709174a5814a3d131811c7a4e40186ab19cf0921951fed524441f44804fbda202e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfabc680aa31f7fba6aa6986ae0e8d6a13dc3fbf83ec5d3d4d9d3018865265ba2d1dd623f0cde15cdd03796245a910129fe5cf71d9117717d6c6551cdba91c70af7b15585295196fa8d41a173558d4802d0cb69556d24f0eda3d7a87c73e9ee7218a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h947dd986a171682248f61a62fe7eb6b7ae01d9e00713855c883faef83ad4b392ac146f27b3d726741344095737f5b0cc49e1542a8c1d05a88735912131106007c3d0aad02f1be1ceaa239b1d30d8005a9e1f5bdd4f9a130008247c665764e532a9dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfa41d0106c8b0242b0991bcfd225c0e065a8f67e6a619ba804b8f2d2f6d796065f90bc67041e24d5181ee1355a726b953b322a4c0f2ad8d3bd5e07e063e339c84daf73958ed88623144258f6039d830b44e62ab2f1cfdcef209a44703ca55f281;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1a5588c65baa05863ab2af2ca133744f6da33fd2610e01f9a62d28ff8a2dac9c6b977314de552f2c02c12c3e42b6f39caee6b63f3774f7fbf413a77a29071cb704645247a32bf9a37be67a80c6e20097a4d47749bb3795fc1c035bf20fc7415d254;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6cec871d275d44dfcf4ba7353ae75ce46c7a638efb4867c133ec985a67fd089c3fbbfa00efb4fd2b6d9ec61a478d99cc4d2b3059ed8e9d6ebfd6f44267cfe63a7d87f2ad3ed4a39097048958278cc2540e8eaacdb46d43235d606f3f89f66f44b3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43d54e0f3341fa44881ff46664ac256d1213080afa5dd99136fd21c8215e3709b3aa349800ca3bdd7535041de71073ac72b47a37d13f95aad241e5b0497760b0d3c732e36054bbb29ad6ea9a7bf2985db3326b6ad65761ab472ddc7d0a16f03bb9ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1133dd32b6d9dcaf0f9a57e3116e0cb07f4c1516f6206e952c195630bb1c1436f9d8b87b6809a41e63348d90fef295a4b57d6ddec29b7e69f1e77aad8a6b967d33a2f5b08d10964f57fc0f78583b6895b626a97bf3401ce83aeec1ebaebd1c08003c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2a38aada6f5fb539cd94f9376bede3ed269e97296c7a23308402fe43f15ecc3622f637f1d82f7c1c649bdd68b5dd354b8452aa751d62844c122f19e2d9a406c94d547a7d2f604163583c09250436bb228368b5eea8a7747fcfb3191a6d92498646d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb575342e753d0d8d5881f2c8d13d7fee9c6789cf3297273ecd06233e00bbfc117d8f2c45d597320b192011cdd9d15137af142b1f4ccb38896176c471988f67e4c1412940a706b4543b56fc4cffc0e882f54ec7be4ce0730459d818b200ea40ffb13c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h812b84987eb20a7b6a275b3aafd56afa485adfe30e713f5f16d9bf2ca4de4e0f66d7a12deafc163b7edb61844a78072972e2ad8c7560ad048f8b4f5d9663a8a06909d282accc59c1d6112d65ced563ddebcb6781bf607685bb1d52a09bf4b297a151;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc839174102daf90a092eef961c40449046c544ed94ba3afe99e57bd5a1e5e17cffa6fd0ca6fdb5f687b8a39290a88e4a1ad4eb12eaf4e8c187bfcaed2ea671c4a9d31374b5387803f847582ff29490d166d0259671a8c9e9c1407a256b5648bc363b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h877920e0617d026a8d766262f66185b7fcffeb26a77ebe1b70e84e2534e04f6ed9913d109a968aae939a7afa4c5d4eaa3ae501153e2515c852bcaf747311bde82bc0ab33c3efc06e28b77cbadc74f7e167b0410cdcaefb144d3215143f22cbfe2df3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffff4ed90ab2179a49bea2aa57942fc8e4b42452fba3a7b27d708522628a0326e9bf83e7cd061405c4b33dec0aafa27e4183056e0aeceaf56a7f323f728426d19cf773eac8f716842bcf589218bdaa12e48e2d2b80b69bdc042398f43791d4aa39c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14347153f46e0399b222210df4bb06826c5f9ea6579741925a7fc83c5ba99895641cfeee0e697393a60db9a3b43a26cb5257c6fbf1397ca3332623aa3517a16adb1441ddbd79ffb6adac2df9f6cd233c2ceec86098e63f62be6641abfbf594e6dbb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d763f23e4cef1dd03d1ae2c6dd485da69a00d0bac176421c07f73c446aae7434ddad817c954ed1d5925a38acfa9bfa966da98d4cbdb3e16f60fc8c1518c7c7f3368f292ee1ce9344e03707d1ca2e7ff396f7adcce10a77f445e62ddcbb3f00a8304;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcd586b97c3a27ba1b873ca2e5655a41c6a680e1e5ff4ff9c75d06473b1fa0645a5171cc97026610015ce259f7a5b2bde44be25d1c9de7dfda80afdfe52379578902ec24b3e0fc0453d0d1c676fffa2e706fe306b2ac16abbe5c08c2e9ec426cc95d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h710371e1a2196f2fba10d828969fb95680959b039c6f62987ece4a4c0e2c67a97efb539107e71888c15adf1ff8a32dda814e3fed632dcc6c4fa5e9e8f09cd3576acf9bb045db2db02b36908fcd1d8354d564f611d81e2bca6b6f8e7aee1122b646c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d482d4e029369ff509cda5b71a76ecf121c00d9c985276eadf37f68204b23fd06858e39f929d7df30d26f6d552248a67fd9aeb0d87425ec0e125443c9d1447b2dce6612fd702e31d4473ae32754cbf2da24d93d459cdd05d8adcce2fe14a6249b25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a15a9af0e68511ed884ad5ccb6c1c0830f2321a97310131020a258d1006418f9c698517b5e6aaa6db2355127e39a83d3389035e79df7c44bb3b60594c2214913b0ec2a5d1fc009be17412d8812614c0bba22c6e8ff7b4246fabda34b05ea3f14feb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had1142176923b65b623bb9be9625d7e7c2d13ed3940b6842cdbafa8660ee01127ef4990c739ee99bce2fc9e853fd24f31ee4ecb0916100b9877a2afc8fb47dd585f0f37896fb07aff9eaa216cda862015941174bc66ad3c42bcc6eb0f68301a3f8c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a2ef36cd33f78fd37a76da66134194ba1e40a6cbd0a682f0ad1e646c8b194288aeb6ba14b60a3705ec8795a05b671f8293a0e871d69e384eeea72a1225d10d9136ee39a4825fa60f33eb6ff239d679f2aaa452f26160d87636aed9998e372d35e96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h961cac10655c6302248167b5b8a95c76a47b03098f32fa1ea76501bb783a9b2e0a7c057f69ebd775ed81e5b96de91ac7727a58ee6fbd7f25bc93e6934dc9eb818570a8d902635fa21097c2ea0f71897b8892f948bac106fdf82ec6feddd4e813ea0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha75e7a5d1fc37584f89036feb6a1bc8e3794fb5547dd9b7707f8cb69d09ca94cc44fd19c98bc165a90dab47ec4f452e776b25a3a815167b91579ce3aa021605a3fc2442b06b1b6e24809e42dc53883a3f1b81182caef7a84c3ac938b7814bcd46acf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e5276db4dcc93d9bb51fb2172d0a129da4ab198d32ef5ce6f43bf68e9f49491a081c6d979bd000c05834a749c7bfdb22ada9a85fdc8c1bab9456c392a24ca400fd252bac4807ea7d2dc07c7d41b974989fa52234ee17d4b80e13833fc87828a443e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd1bd7c4e5349b747319d734c6ea85c7c3e304f07f330eb206268fc523fca29ffdff21cb2786d8721e6a6c3ddf4de400e2ab1196d5d1daf7df2d25a038bd50cd05fa58016f840eeb9374bab6478de6a5fce42458a10af1bc123b6316fb471cbeb0a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72339458a244230a547d41c717a45a8c79b86ae01eea09b039bf17577841b60b29cf8609f2375f635a7b860e968316669ccf43912d2e2696c0551989e28636aa82119c2a6417189257620daece05b7b71e7797996574209b83a34d57e9578a311687;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h261b70d62738cbef82b15c0d0846e6b01f3cfa09fd29030a1138c2f9bda01505bc4c220e0065e2ee8cdc4d334910b9216e693d12e8bd42903cbcd9bf95d53e22830327f3bc02b0d297cba4021109d377312e639aa3332afd1971ef89a451dbd6900f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6eda24d02648d9c1fc32c12eaca2a7f967c0ce511100b2f0eba5b3151b696a3e626d0bacfdf84a72804e4279ff491425e8dac6137f39dc46e9a9ebdb9212821f62c05e387fb266a114b93a66732d055c749c7819200af730d14aaa331e25a4b5b3e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc092206168c2e1617df1856dcd7855407e644a947b6bbd8757e541137e74f1deb4764a6bcafe901ae56a42de84c4401b48e2639fa20dea2c0aab0d842a3a89dc33df4982aab656fdfb3b3d6098c2e97456fecda1c87f4cc177861ff7ffc3bf3acc8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e549d2344d536e5c3e7c47b43175196ff520d53db73b92938df0e0db76418723d73f7a328b9538dc60e050b4e65f6b374a744997ccc22d9a585f1ba2596d8c84a64ed376f0af058744dfa105c1c466e4ad2a4e71a6e93c3deb7730d3b09ca85a386;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e6e441873ed80940961ad14cb1545a95500808bca8c784969c41a63f86cb293655a52568bdb672a5d7cf890ac3f5e865d1da4d46d1e07dada8e119480a610e0410d2be284258a680736d2a3b16b73a3455dea522b9db2ebe2dba6f576d9158d3d9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51da8685bf5df5223003a68ef329d2f925d11ce36ec68f2455842ff578aa8acb3b817f7a8419ff114f471f1d66c740330b318f03950a2cccf5ba0dd0d517c262105460615cfee1ff7d841e6bdc5fe9068f76e50b17a96bc87fe68982bc256508f19e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf3fc2c338f2123e2cf649b9887dfc139c6b6cc8f2e6aa853ac699bbb6019d2c51d295b52af908dbd41564f58b2461ff7f750dc073a3f7d1fe0456387f6db8e63d63df4a64153cfca7a2f11d8ad0a0f4b9c45a2ed89b358c973c1d3f0e8b30fb2b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c007751433a1314516830e52e4e6d2ef2ea53853b42de099bb29d1c24d0f8505514df2bedf709bc9db28104f918105d1440003684dca3a4fb6b08e0742b7e854472eeb2460fd5cc26522be0f3e9ae6a6ccd444bf762ddd01117a29b8f226d5399b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1521a9bbe955add18886f6e268db15aef430823e83983f8f6b95b2caaa74b56a58bd3460fed2db0be2d0779440f35b0876e3603e7985b64f144fa012d2dbf4b2a93c5fd904cc51be551564faf2c77d66de3db7a940bd21f250da516c2a6ad03e88d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha297b2fb04d00976453bc112b99c6245e1775f2f24bdcd0d11190a3c8e0ec22f06b6162509f5a9c993bdb32043ff8425814e0bc471b1125cc2913bbe6315b8f7a7e26dd13d5150add0b9c03a40f662a7a21b66ce642fee847094bafcfbdfe0419737;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe5c35b4af5fb9794aa1e8de01e1512494aed4b30269f1c2d6ade4393920182d9bc61fde415185423eeaa308c9db0fcacb64b883aece02478863681e90a77642fb2b83ba41ab8bf74deade10c44650daa13bd9ea663142c64d751d4b76646ca86a9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f91399ac70333d0721b30436b6257706e4a19e3c8eb63cd1cc81103d0a28f9d6e115cebcea4312b1b655169a0cae29f22836079a392feb097ed2dd6b07301a2418bc738ff8678aecc05ce4bded7d2e5e5c58c1c7346d39b9581ad0fd6ddff97aa1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4729e8b6ea57717d1281141007a1e37978fabadac3be4fd787948d79bf7e6d0e5c3fbb492884766b99c72d1eed4e439f92e018c203120f90f5f8e488ccaec274969622164644f3213255f28dca3bf47898ceb8e54f2cc97e8af2930618f644a5e27b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24c3db1826934948c286d04f28e1f7df647fbed9faacf666022501afa49bfb713a3fd80238c1cbde9df20b7ff6e364a162e894407c6548389e327ea52d5738c5a468eea6c57aee5d4789bbc216bf9cd64e93647dcc26711e2a55b46089c450d58a75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda4211e2e0991347528a6b9a321060aabfd7dedd55d31e92fc7599db89c545274b398e137a6c52de054005dfa4267eefc39408f0ca0427506563b4fd2342fb324323e1cef215d1d5ab1a157d0cdd7c50814bf5a67c74e94d3e5dcc7f37924397465b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1eb7b1ac6ebd6a85f0ee6e5b6451c597c79a4adf6fe5d69475a52533be0b6b1f3408fbecda0b6059e101c46d6d7d84a5f434b8b94063da3b998d1835cf779cc06b960b298d8170c212ab287f7abd82b56a49ed7a38d476d5bd7ba2464afaeee69cd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7580a5abb4b721388ca06467042678db6ac957fbba1cc64319e709373114fe44953b8a3dc01dce94f8c9fa34b2b0d1eaabc9dd690f96f8f74edef7b7ed6e6a396b4ca78e82b1ce50f3726233d0de75797a5ba4c6e17fbbd7b99da62c25eff94a4e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb303148a9d723cdb25d06427675585e5c647372d5ca325e41b3a0546c5ac461f0bddd54c617783e9dfe5f1e8d6d1ad0ff1995a602e09983103eed3ee3aa9ddcff0af844c78baa92000d5b4c5587df2c2d999fd9b3dc18008191ddef149ffe65fa13b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf019dd82c24663c7f0f9d206597ba9c3257b787456b379369781bf3451b3528e7e1879887aefa1b7ca54aef327953c348a1df548b2ddddd247ebc4cb79dbb5e66d1fb13c823b4efe3eb2e4c1abde73d43337ebea917b5fece1442f1bc0746ca64cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe222b60972724cb1f31cde82617a325d9530283ad24c944241a6d4dcfe9ebe491304e33e9c6f98cae5b54b54534fd62275f05c0161c40ca2b036c74448a37d9f010f02fcb5a8429fd7f408a24943ff6287fc3551eb7c3cff147268cae75ca04c3e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd1da8719a8a4c11dd89b2ebfef9a926f4f14812970ef2fe11e1f1fc8722b92fee9711e8d5702d39caa1ad7be1ae46e62a699817a4eec8fd2b8e66839ee57c970838a1e8d88cf2bb36c3dcab6a74510f19baec17155b9ac9618cf19a7619aa933e7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67353bbd6cebc989811586cf83ac36de082b40637a413cd3fd9313394d4c78cb75c69a261c666bd8fc74737cf1f4397208bc7fcee4062f8e993257a521faaa730c184846459ff513f74ebe9c5182a0561ce46551db32e58b33cd5606afb80f9ac7a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6af96990bbb7d7139c0796d00ab659818f40fe0522b0d239c34654bc5028deee58ac1f138b84cec49f3b9a4b0d08f5337bf74f588f1b98acc55df85c420a72890fe9f07fd21fcaaa6cbb03b45b7836e1e15b9e1205b61d568bd3902b28aeabed3ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61d0a8f28f44863d437fb67db829675c163c008cf2aff9f5adf707253e24969a2a992abaedda0a6c04dcc3263e961372ccdd205b4a5921343c8a8253559045d272e1bc319ac3ebf262cfef4ea1a87c053e26df4e5a64a4e908f800b9639ed7c37a28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h670bf64bbd9e9e644e62df9cf9d3a474f5d83100d6ea67b616655086b661ea43d8a722f69ce101983748968653a33e0b880839070a788ba528a6db17c5295339f7cca6277154a8cb35ec896dd96617b3951c27bfc1e2655f4f67046fa666e16716a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc0fe127a2ba8d8b560d7c8d590d9db17ea41a1ffd0d4370d44e7b90af2f3687ea9cc80487511af79d93aa80e88b5d02d59a16e74ef93d3dcc224a13345c06ccab7f85f46e139e3b7a31d736bff102c168bfdac68701817961fdfe50aa91f4611f3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe49c8eca03b13044c5513bb78c639b6f8f116573ec0ed2127f3ad425869ffb202795da4965606c0f2af59147ba4ec91f3a171e88279042130f463a1e28ccedd60a1bd76a5906cdd34fc573128b702047f212cc4092b23a812d69fbb3a974d344c3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h962d7228e285c622cfcb749cc195a822ccce3c58ac2119feabd82477f16d014663789905128f590d4ecce7d55a62ec869610bb2ba09e7e617f413b19cc2ef85d98ce010a7a521104ac6188fd488855f5a0f2bbe6acdc7c77ec9959b67c6dd5ee2e30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e0f1cabf63c9bc4cd0356ae14fb4b8ef5af015539bde0704d689c24274bcf7481d8c0261dcb828dc45895497118d54bef215fe83c1e5f9874a680e53132bc7b809a87bafadbd44b379b0c5beef24291b92ddf835f7955eec3ccfa0e0f976e8e2e21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf961f13cd949104db2437a82a4684cb59195ec1523f4b5f575df6c32ef1f571c542d709f5bb07bbd6017391c278467405855f5124658ff374cae800af34666f0191402985b78d5f4d727c438f275939520e521e0e6cac91eae1964adf36f774115c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e8d273a7375c921c6820802ee3ebd699253f33e4af593157bb1d9c0fdb8c5a80cbbdf1c04a87330921adb50de4d5029926afc3eb533f1043d6a675efee4de66e60d0dab8d7afdf3873b64c87d8c06818523c32b0c1bf1c294049eb3903adbeadb65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c56765b6960a0f1b887ca8366bc1d74f3a680ad44d8b8a8a8ea794d3b874becae6350f3e20334a377937955380943ff1fd30c6cec24c8518bc43774d6d59224177a596cccf5d219ac9d5bac3ff52bd8568b34fec2587025ee2487289e01cd891242;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h273a21274ec6da7228ab6dd3daf9ff781e5edc1388de72a21c334c69d8631c08198404a32ea61e8cd5e5e6faad7749c2b99b9954a5c41c9bbcf096c5fb07ead52b7768c3daf6e1f8f6319d34fd007e394b358a365c2395fbc850c7ebf38642704cbe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89c9c6fc0bd78b269368ccb0335d28e88a76ecae8734f905164f2a1de32509d3fb963f9326b0ffa34d79e955d3d8dde7bccdf9ff839e2f2cc493b039597417feca7610b3ea17094c4a9f287f1974dc22a70e68f6f061be5fd5afc4b20dfb0b5e0646;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he83de15b6aefe32e25e343fec642892512c7375a4e33f7c3306851e04b27620225cc044edd67a40b8c5f5f3898da49926399463f5cd2485d93114d0f720b2aae1b22d37eb461abf4b25373f706ea4b6d210fcf1ca1d9375ad7587273b4cf45f8e3a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a9afcfa958b26f601f86a9e33886ea188af171e5a20c3a85cc1aa7d853d2a41814878c85de86b4a8139e7b4b152f08dcbc7d47143737609d1836feb74d34cf2f0f8bcf64b608a234dcf670f44167109f54109081b9581e835cf8bbe708ab3d2a499;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h534db71d3d23f146e19bc0767ab58cb8f6d9a0a289cb1aec93a703680fd1144176a06c5e8e875cae226e8f5836ebabf1ba8b6101f2c75b21f38676d80cf2af434b3d1f807358d8d512d77a66c29f18fa6ab2171ab55060b4939a407f1b24155c18fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16c71cae8f4baa08d9863f12f2ed448255c94bdccc8617cce95c8d449111a9b3048ea70a1473caced5e55ad58874c935ccfdb607c677e8298bee6f17949e93d48da51b9cd6e2db2c7efc6c9b0f6160d2a70b37d387bf110e33e23ab0ab288e9f666e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b4873d6654012442b7ed22d29a9433052b5efe8267c084da8f5e017d82a0037ba43cfb55cc1e3b110c5a25b1b651b3fff07ff077fcb305327453dd388a9f96fd7901dec115109d823c7ea9044fbcb6d610cec7a2bd6bbdc92664930e031b6c6acac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfea939a4422d2d643282345e9fd7fbacb720cd9b0e7453985f237197f2c35a14b2eea5a274687cadad1727ccb0fd97bd1a969b30aabcadf65245ac9a2e90abbd2d289f73cfb90855116ee3ba44e5fdf19cf52423225258adc38eff6c692e4e6d852;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dce0f8b45c2bb3d93134ae752f6b562aacfc05d9adaa149f82f0aaefbfe28cb7b042056455bbe850767d2be81c088c53950c1589e14778d1ed050e912726b892c302763e3722f86dffb6e6561434ed70ed12ede38059a1e4b4a93c8e62a9c8df82c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h493b2e43abbad219947ec9ae03cea5e2ce6eb1cb95bb56ae957c2739477a554f5a3ec183076bfb646c715180d53fc763e853dd45effc75d2286a8b5d03333bafee78608edbcdcd1d352d92ad1037bba09f9889f6eb4948807fffb670b94d5fe20bca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8bb91545df2eb8e01330a0a8700624d8b7d1b12a65022713ab008d0a1ea8fe9d4facea9df771d3e6eb72b36e97f33255bb08f17f8cf26e2b210249b7d4f476e066b6843c18c7a0ffe8a420b278a100fc4af2ca3e5c8e3d0977f3eb304ab941ba6e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e8235de28cec366d8dcea28002f0a8bf1a1af25375fb5a2680746411bbc83c4e054b4a87346a65848c7054f5f9b4eeed0b4d8a1c97f77e06f98dcb37a7e7f61eaf3b0d82728fa6c8c6eca3fae85c29b3fad57b9afb5d997b12d250ae6cdde5b6e48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b6de9f9bfa18a9c3f0731f65e436e70cb7fdb504984823c21570de0c9c4fa4a327240ca31fc5defdb158f4e1e3b3bcaf4f042677032f2a5cd2af51eeec66a5e56656150bcf01569d539c8de84184d430e078298d2471e4f8b40102aaeb7a8391696;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafdae719fb4392dd8c6a41b7ac902eb59beab3e28b7d648dd221782352ccb4323f6ae8c4673fccdfbb849b9ceaa906b789bb46ec85d98f5cbed73afb4be01d2ae7c53be5dc5843cd8607d94924bb6d9ab6961c9f6283331259757d2b2aae1912b178;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbfc3e9b519477e56500498f67d3ad7a2f27310e965a5c8f7eb8d83dab06ce7ce1121c81a8dc18eb7bcbb177d4685c51c4bb2ffce4f1b66e2eed4ad5966e409dd3a65a38e242965613cc9231396ab3ca8d74e865f34916feecb16b2449765c75b1c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h267de51eba04015242c9dffc72464a07c6e7451a213fcc0da04c76c5e8d7833d9c18108139cd7e599d5695c0f84b2d1c600ed066716303c231679f059308724bb75c9d1791d337b1dcd97b9a6ea282372ce5319b7d22195a3fd4923bb3a4744d970a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880f07a1ddde294840a6d33e796126bbc4b7d34e0a778d157f3477e06eacb79c4cdf857cc602309afce0d732d44536bd0b366c88b25bcfc2c6f2a31e08db861725c3d06b0029c8993b69aeee27aaf36d1de6a00bbc57ed41f4df29a260cba4db8bff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18ca38705187ff54f2078efc30eb9b147e4339637cba7626623eca1dc515283f93aeb9b9bbce23306b51699259e58a8cd56caeccfea5a904496de0c03b65e322ec38d64e9a21ae12a9f6c66631430244f28ce8de7206ece5746f385855374e2fe6d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18e172227cffd0653112c0a4b25a028776fe31e579382fc6ba85f2ae268db46a9f1f3949f25d84f98db4109f43d2ca53101ee9209d9442351d9f9935eeb296210266e62b7e9500a792fadc68bce8b9dceec1e194ad3e7260baa4e9c44ddf2c25042a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd17aca65c2dac34cd71e6876925a99ed1c36db0326f0b5d78a5d239bb8660a7928bb278a87f014f600a7fa63b1a53b4e17928aabbc03f976e1cc03b98eda8faaa9a95aac246f80d7c1332f2c7a794decd73e7ad56e3e47bac4bacb3ceedb6f6f4f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bc86f65e508e0ce09b2889e33390a3117a90cca5082c05e253a0e18f9c88f78637881dafad94f4acc75cfdd30ca10a5f817f5f8e4cac711d45215bf0ad4699b8de08d652431f641f84fc7c295ea73c65d10f9ab991cf4116ba27c6e07c43ba1702;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54b85c078e260b9ed7837ab7963cbf00be928b9e9597a75db181d1189e3cc4c894ab87f8d4e83bd370819b8ef1fbcca5868abe7ff282a7b4c928873ad11c55ba10721305bf6add425b11bd6382df65cd99c75a96482dddb50c7901032b1a9d501c3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h518d6217722c500b6bd58a0d5848e04541b7a76e20f2e60e6cf84a28ad53cc8df8e74c7c7d12e9ab66e4f5b9727f45555f490bb8f065aab105553ef40f1b755258af5bee388474f2a709c27d79dfcbd830b042d179047d7bc4ded75c56565faab719;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h465d4b126798797852282bda9817279d1c1d65fcaf10fc268ad36bd8ffadbadc9b85362468e3e3135a5a28a2ffebb4c2cb4bf73ab925cfb8fc56f15ea9b66ec2fb346d59a2788f868a4e9c4445024e0f2ce508d6f42bbfbca44faebbe49ed0ca1595;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd45411cd988f9648d4f6d3bcba37aa64c235190c6fc1b67b6cf57647e8c12b6b3fef9bfe8d43dbf3ebbceb233dd48c2d8b0bd94b3f7f7c4abe5c2df6fe408d48ceba60cd81f936a79ed3746d5e207be15eaef5f801c84acd77820498a628eae3e72d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee85d7c094139e59d3b9cb3f91518ff84f03c91d8f85ab7edd3b94b833fc157d3006f41185ad1db1b1519b640d681ad7eb71636a5ee57efd572ad9bda840078fc9134381d1cc052c560950e98866256a8016aecfd9e5efc621e878cecbe31af5efa8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40407c1fac53f6352e55418630e447e31ceb087132cf6652ae24278115ee3fad10abb9441ee9ab79d0a82921d2ab3b1ba85e698448cc029bf4d6a02f753caa2e7da9e6d6c23136dbf3248ab403e6691d0797b14fcc77305f198a64b810bb7a3a860c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96905c3ec72f52062db07442092d2d3a6601cf923c6bea91eb7cc5c59363f6842bfa18a42de8beb8b29aac1f6bee0c30e0842ee6f709992bf656ad55be0af6aa8705a3eefa39477aca11c65762a81f967e1abb3a14c85f417f6ad43cec4649a99f84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6b0b298e93497979b992d91a794e465da8fc45c8c5b7bfe64380813061a2ebe918fc791c45b9ce2ecbfef32c2b61e4c34acb88709d400b54b2a27944d7c327aba49e29845c6823d397231ba91f145b25a454140d275b2fc07f4eb91b99f0ef95d26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd94bc739b67e6fae99c61650c1d5f12fee47ee09ccb2bc613f75d22d29aa3ee1a0b672e2ee17f3b61125e7a4e46bade1a831e464d274fe7635248690ccc619a6726993ce45c353c9bc69575fdfbba2a1e8bffd89bf5c838b8eda434404d2a83cb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12ccb913da47efa266733eb159c99568b7660aeb8e7c1730d4a5c7562d30359a8270134066e19d178611dcd0cbcc9b203f8c4d3d80a1de5b0b95052aa38ab1ff7d810ec7c24756e0559d446611cfd86dcfa1879e1312026c6edf57809a55b1d9e76d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ed3bff7ddf299122b109ae7926c3bd25ecd1fabf1a738f14387ea1446c2b20931bb8c9b8d06162a8cabe6a91ee7f342dfce50963f218eff657a6b025fc81ce50a3306e31986b892c4e4e984e0b4dbed8efa9d297375979a51589b7d636067ccb913;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e552430f6cb69c77a08cbccdfa7648262ff936f63552fc5abc120f5e4ef783f3534e4a69ab0c612593bd94d92d81de3d8a01017bc215cba3a2b75a545199869798dc7d57b32d8c63f7497a8b5dab23cbf28cc5e850faba1ec87a0702239b9b31d5f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e18c8e6018be55dc277d06f931ff49cabc84e1c94a6c5c9fd7b2d04a126a2589e5e125406ba59668da43d7788584e49bd8b90942ed79bc84942072585c7b100fdf6ce6d1f9ab3df2742774c29e43b88884c386805631cda9421b7ca93ea95b3fac7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac118fd73436c01cf4869c221ad759c515bdaf5dc2499a9544b49645a7ba517d8aaae9c49e5b98d99b1f0ae077e8a815ae5e2b5fe9fb1be0fa142b6426603a8a75c5ecf981d810fade76ace3e9d1401ad429800af99eb61f54000b1a6cd0bc405c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ca1d71fd06d68859c0d4ff624b87e42b8d0717d05b2f704eed0a4284b530271bd074719a51a739efb52ce01d54ae80b8aac211e6b19152171322f4ef4c1b1ca7c4656af9359dfa4566ddcba879263608ea3861a68a39359def48b03c2542cd3807;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9595c655de40b34eccaa6e433704a4893fa8cce26f8bdc63fb9f27665ee455acc5742e53a539d46d287fd348b3945ef7067b6f0da27ec435750cf7d14fb1fe8001a49a5ecd30403afb38a85eb4a892415e6ba815da28617c174c696cb436231d06cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57efaf0f3768c768b046c794ffee1be2b90101348feee68d9c0b05d48598b62aed9cd4e9a1cef94780373dbed3d343cf1dab2eb88d44912677d3c9e45cc1ef1dd21f80ddeb922b835cf9e7d85dda5fb0bf6a87a889d11b2905eae2833bb308f403f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e7b354d89f97a449c3052f2d58a562ad4be4927ce98c5318f6be2441a55404404d76ca533f4d57a3ffef561d4cb52120a4e3aaadae6eebc279da5f925f673ba41b54680ac6f6ecee7a839aa5cd2d4ed7bd12988a1b71355ad71a8afb57fe9e74433;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3aae44be9a672e093903dcb5fa827398e253782f86fec37b0d79fee947fb5a34a001155965af1146da30c24093f3eb702614a722d115289aac7440eb165eee56e310c450528e4d97d92dc1546d006f8f02cd6f54d0a931a63f3d6ba96d1251ac2c83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd3728ae57036e621dc8c48033be9d837526c9945e38f958bdc4677491364e35f955ef24aa2a41ea13290e84628beaf82dfad90c24c66c6fce47cc841df42de3ad238c359a0a8351ba5180a03b43fb9ba9b35c3de740969640c555642ff5f98573cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd182c2e28013b5857f35e0ccae35b49c4f836df60fe8df98787da71364ba0d84baa751f87184badbcfdd920410e2df78fad286fa50df397eeb188943065f008bde30d47e4ccb42f97e1d28764744863553ab51391a032951f28b3bf927bb483eec87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h957095000be051fe313973c522c4ea42b606a94635ab513dab96be86bcc23da7539a99934ba2a25f5c10e07011fb5505bf962964684328851ba6d6d9373153bfb84c95862de2b649c4e1f6510babb7580f78015ee0e333b4417623b6ce1a6a880039;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c9eac4fcc6b3d46611a561db003f3facb063aba5a83aa1c0984668cd75dc8f27af698981284dcc098f13546005cbc1cac875dfe093d13b53d85520231d5c938c1ad1bbffd4f18f21f3454b33201a7ac6177974cccb4a3a5c30b99def4e682a2083;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78b05ed48f00147ae3d92a730e40c8c638997021aec14d37b362d42a5e34629532f8980109f238cecc6ae552d00edbd539a33cf3d1e50cf84e9a693b6b60e502fcc52506406b2d1f55895651c9fb19c20d7b3e17077215d1cadcaf1c5f0f599e7ed8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeba2a4baf4dce90151d9d800e33ecad90a72458c4700c208978a67d334668b8ddf67122c01edd2e5945c527579366e41e8dd2670504454ee381231af7bc8338d359520c6bfd4dcf1b222b14f4fef5c0f815564dcbc6dc9c96c6c74cceda31c19580;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0857b5f00f2b8b3dbe022bf66a3ce0385f8e4a95fb5c827eb03e3a6287ed1979d71bcfaf12752f63246145ed7f802436e8797f2cee0be5135585abccf37297850195a459f7c529c0087066d360a3a1a996e7b6b5c1f83c26bf5094414fc782f4053;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46e6080750f5ec65f8b4d372f614721b2c03498d1123a129d0197a4d62665d93e8e93abddd17b8ebf05cc1d5ba82105e447d4b6fc54f2839b3c875744971f93613dba67969ff7120bc4dd05986d579995131615f1fd97bf2b828d5a140668989cecf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7df7b4d5cb638c80c28fa1fe575c4c7d6bc4c3e4149efa10e864cfbcea20c9b907d034843ed1806519309dfad1bcc806038879bdaef745fb64f82b8c1aaa4eec757f95199c154692c657e6c435f774107cf212468a2b61eb718d32cfdd775811a11f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d499d8a2e4b08bb97c7b02242f02b2c3f8c928e96cd984ac9e5a0f407270d1a407faf866e707797592efd57fecf563e54655fe04ed53c7e95700bfd46c8598af5bd8f68b43d8718c5cea6409a40d3740df460d58faefa28376a941193d4b69f56e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ec62de597ce6355c7e85c7b90184af494b334981eae75751af0a2787c838df801eb380d5d123c8678949819e30efea8d67606b42e8fe876e74d9cd568ec0ea93228798ee01769b2e8f4638f540dcd0440ad892cadc1a5d8b4ae6008c77f3c609172;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h991dcebb986f8d0cda01c8d84ca20b74705fe8fea82b7c276c76a3264fe996788a4281d2dc53ef6d1d8e100a0eda5f48f997b073b83692cdb3e86a047a70d2e3c8f3a30ef2467d35a44c0530d4d59fc98317404f4b8cb12baa7ceca5958cd8a2dd9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf03bbaefb337549efc2790d794a8b60317b231e7810a4d8b544c4d78c388e413c22b7925c80bf44abc1485b5e6c8b410e1ab88660e208ed481c85fd65f961335ce2f1eab620a789cb69dcd3e89823d516582f9a33e1320668f17bcd0e219076e03a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce2b751c73727af89084cb36b857c07fc0edea4e62d45070d8209e1ef5c623eacf1d008ad2200da24a7b573f7b68c20ec5f4377545e1816e26bd208eeb9c3420962c1602d99040ffc564176b0ddbc92f2fae0f436532fcb53dc300fd34da09c8e303;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa3e41b90b4bcecf7cb721f9e8365dff7fe4334ea7c0e01424f2091392916a83240b9e85e4a9840e8732f6d1a7279cf8c8c66dc0dff4b4bda101c2e5073d264a227cc514746985854d25fce12af837a2212da9fffd92cd031b35bc4d0f1e713013f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6178fd4792765af6475bd08573aed79baf4a178530c086707cefd2cd5045ff615f07756f95f0595e8ed09b689707eada31a7c4cbb57f0c13e5d764e280eb39217d9a82368ea0b9a6f47c1130041f8a7458f842ef587255f4e61ef154eaa899cafe3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha880c004d389da0e9c5037dcd180497dcb6011df6cc05cfa1832effafca0bca2dc774a9675a0f495c5d5a9bd5d95fbebe3d9b01daa951c04d0290184d04941e2606b8a879940456fc78949bdf8b248284fc7495e13f8077439ed50248d305397b88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8da7d63dcf83fff75c4fd7a0ee730bdef90b790a8a2122a7ed39580c0f07a7edf7b3f47088fe4fd30fd731a35a57de5ae91276c3d2c72b1b8e97e1dd521b25b3ae74e1c3492eb915b4b2e4f48f36907dbb1e678d1ade21e47d00bfcbcd2c8a9de710;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc42d580faefbceb8b7b867fcbbfdea056807d22def9cb279560914336f8c3fc5e275bc02f59a235acba2e059f90273b73536e48f4ad1c22c11a972eee2d60c2d9173cddeca8b1c673ff76c3522dc735bdb32eb6374870b3c1f9579d2395423f4d14;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed41c8de91af665b5d3f982739e10e66b4d22d987c66d5bee67d53dceb04bda3c83d226a1128a9cfb7999ff604328fe439571ca8ab956b68f3c5a80c62c0a768dd20bc15ae126f5bc49ba3959c2757dcd9b3fb4a12a9a620c1a63b0f71f52fd393c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44713eeb710e50818c52ff4fbb7dec748c970e2cbb822e6fe4b13ada06b84b246d3be7e9bb5c70a4e8b51ae966149418b40eefecc380170b72273f0ae89dd409e739d3e1f6c2fc13c4045ef49ae7201292e9274dacfab1680bc01cef29c79535ee02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6243da31fa6f42e27be4d34af058aec437499dd0f173393fc9c62d3d27eef99a3373dba01b478fe60ada415e5dbac9b810553566565937ab39d9128d6221ce0f161910c29e03c571b5f1480ea8753544c5e8184fca41bfe7f435d30b9bab15d736be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16ab0ae614bd1fdfdedcbb5995e8a14d6e332f3211232dac2163815276cd7529736ad6f4fc4729d9e4bcc9aa26f4aa7138c4f6ed5ccf820e5b7a9fef2b71a6991a56ed75bd7804e550b633dc3f8b17aba0e29a168998716f14629faa3a90f5f892fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20061ae74307121003b3f9ca98dd3d1fecd25d1178c8d70b38259e09fa524d74d3b944cf9303f0cf85cfb1b8812d52d09acab934c5b1486cdff345fea35020786ed8a26f2f7cfc676879077231c67155904460453806ddafe28f5ed75223b883c7a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha66264305d44df8f025f7346422b9ddde530c49a4b4dba2114b54dcbcf26d0c173405c933833b0664d0fac606099daf897321ac98a68ba4f119e95e30a6d157a0c8962130d6a2324cbbed3abcea9d6ebc9d2d5dc3b2d684b19d01eae73af983c6638;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd334fc0fd927bcc0644e19c0f76341c4a9f75aba5e34864dd0015177f4fa4b09d00bb92397dad35ae9ae225499297ae35c67299d530b35b6d4da7608a3ce29059f62d35d75d0b938c51a5ff39b9632ce56af3fe8747153a9b640dcc2a58b944d21a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86262decf1aef98fdd9adf9657e996802fe3f1d48406b2398ca2db52901ed6312414912f086167d3e053c0b5627b7e9813ad2d937c192a9f66beac8da51612798d037997ee30c3c2d1cbba9ca7c41504c599dcca0763fdca9fae1c23cd5d2829f5a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb60d6090cca429f0aef4a21c4c71a3302c23157afb966c5dfc4a51689963c90e38c6457496c151b3758558e26d2e9ced54efc8b13667b562a743ae51ef7e394d11c98c99f89a4f5fcebbe70cc396387bb014b2d63bae5404280919bf8b0ea4daea3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dc1bbdb70fe57e7830535483a29b70104837d1b0f93b0f7f973c85fc55fb9c0a646ae12e8108722332c044982ff22bc1d07186d53ea320603c4473b9057940bd91f8de49facddaa76b333e1a030a72e2ea12e7eb1267bad71594457624b55628851;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d6de9517ca1bbc85d9beb3ac766f481a3db7d88497a53f79b301e634d1439177acb07dadc5f6516b9fff152f62b76a38e155eae2a19ec156d2580f9271ce105b70b6fa4fd78081c0dcbec9499d91094488aef98d80c233e88949be6cafd9421ad6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76cb5a10e4c809a8ce06746af798065e5e6f0beb3645cb5ca59287579d8a059ffa1407055a110ac04ab72d61f0c7e212f9399a8ac4d2436ee3efa191a7c664e00f36ab8091574121b0bc1be73236b4ad57853b1f03dd0d9fda5f6dd1e03bdcf9b72c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6525798c99af7e84cb9792f93f4aa33f5fdaaf37b8263fa22033ffb5854fef8eb10dd05462e287b55b6e3cffa9eeb3535e8f900251baa67529a93135a4764863c1c5e777f1657f493d89f22679b1c53ec67a42edcf6cdfcbbf6d72b5ed35d74d6f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e440f4ef9395073d9085added0f11bd05e28bd35f36920233014e5342063eda40f820cd7537fde67e950d8ab7165ecb30c9b61eaaf3f99fba662c63109d9d550f1f94b8aab8820b35dababa794bec84d85af14ac7b6f1edb18c3fb3d673f8a2a3a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd339c6e78d170ea213d5987a6e91c9d4a7dc6734ae6fdd6a45880a39963353b99a6adcf0082a68c934f8d600cd28e3520c3f3d0da396a777a504c9797f330bd76550de985684896c254c4a00145399d4180a5ef2a0486cbf3a8b475260e0e226021a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1213a62f519861f697109cb0b0c11954937f30f074afa71109530b255171f44ae3af7571931b7a1d058d1f01f3015e5596ffdd5f62d4fcd2bda4e3988a11bb16b3db30193e09c1cf1f06db7d892f2cf17d4b3c795a7b5c72822af841d5db74aebfc4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33d8a7d32ecf85c87a5f0e52d0821de2e9c684c3ffd6dc3247262e406a745984205270f4c8d089d0510fd130f4d59e9b33865a6f90a31adb7c089a8076012823a05ed158c55f5fb9d00067de1cd6e615399f2febc084f3734096b7237680fcd0f440;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a4cc0a14e6e9cdea5dba38ec3171dc6c128e29c14e726be9ca572e88694e98bb22886e32062bb0b8526b22103cc7f57fe4dac2e5e2f164b5bf9497c911b9f0733c06d7d5c1ced4a714d5e9cf0ef4703f4b6fea55511388c1cb5240acca5b8e715d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3333d166ccead16de5d364d356d27fef2aed56818286bb55b17890425ce1aee9da08a4d0666a60201582378078df30ee28780b617cdddf382e426f1db3f51c2839ddf14b4c348fde91a70325dd13638d5c26078c159d556d6ee19081474c8d450e4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3321d121d31c20552b70d454e9c918ee53f5c3388f6c9221f2510f012842c8e75037690696823751c6d6abe4d30e86a2ae00a836f5a9c0530ee2c4047118da1527a5b7d09565079f962084161406a45e21acf0964d32d9fbf94074588ad381986b94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d56f28c3fb3a8d9124e934ea65255264de12ba14519c46c07ac5cc299ba8277a7ded2fceca4b4c95d7c7c18f2cc39c9be5ed0afa302e70dc53b65530ba4075cdaf09ec5032e2394098a769689834b4e7206495a2728ea56b0748a1ad5638cfcb30d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6010d4757cedf9fcef9cb4a228c82fa0812ae5573c1e162c9f0353d6259068e36b60d3f40201ee3c2f2f3769000cf22e7fea20eb6c69ea5e5a2a7dd63d7c8e6a49b8c58887bee23d13c2c8683af77fbeed584c13565674305cde5146c4b11f6f624;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2136b5ede0dad30168ad5170b6b2ce0759d35c888d2303ac7f701a9b46a63d0b397688740d104dfdeb98e4915c105b233292572aa541f2f062a4a0de36c9f595d4adeef84db39553332ce7e79215d2d8a97bc38cf723465bcfbbc088fd2393187bd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c7953ef3765c178385e5f6b180e51981a6d371b4dbe4675d750a5bb37bb79383d5bf295bff1a17cf0e2269ba1ba7f1f020381c9ba3dee95f9a0814f54af8a929b59975b71e744fb603068a25021b23a1d49114e5b892f3c5432f2563a50015ae6d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aba27c28fa3ea2807d7f0c6b52ab94e4f6d2ccb4152ab6c367309eb84fb572e72eb8c5127f36ffbd8e77b18ee0744101a8994b7b3ae139391013ca800c1d1216eb352df3868e9574c82161db465b5e032f82aca9ee3798dc66c5046749d3632f03c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73acc6bda2c6d54ca768e6005fe8a480b32907a6b6872d28b7800b0805e7bbcfb36188ee99cdbd9c415a6cf02b84176dbe985d521eba4b94043720ed638cfa8fa0e5632a9d147625516bf6ecb1c9aa2eed01a11b548c5dc22f939d99b34a2db1e6a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12b352e6ba62d505074b6decd42a502e989b732c43b7ca57c0bb6d46884b8d430158210b3a3b446d4a6dfbc7145c6ba286d70e943359aad4a11d150333a5204630c2087188bdfec8c600fa77dbd693fe4022d67cf9133abc7ed4729c07f86911da9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15b171574287f6b0ee7a4a773d3a18ff514a78510b87f99a74a889e8a105b071d7aa75d93d5bb9dff72ac00e1a47694f14cd297d8bc8d15ae76c86ea9b2cced01a1ed36dfc122cdd12fb8ad133f0752d1a1b6ea6f934798c75506560f33905815561;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab7f8cdce2fc24436831cf43cd59572525225e451ce97cacefc2fe893aba85c5a79207f5405e2d47f277d4c273c82056c7856625b471f8a59cc496514b69b583e73c11f4867985bb89d007c4e1a460adfb0b60772add0ee82bf4a4c46297a37492f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ce8a71013688c4523f0774ff8647fd0c222b352e5ac3dacba58038345337a818818057a066e5491064747252957b6101515ca2e1869334108c166b68f6716eca90ee45e667457a20d2fde25bcc3189aa1f94b3b341baf7f3c900f619fc7a05b62ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0efcc1d950823b4b44a22e33b695d25fa643b8484b2ff5f5242cdd8d6c58c8708d603141edd89f90f7ed7d798f052d4addb63716d5562ddb0808518f6280a33a61d731a104e1227efd50cc44bb227dd9257735e5284915908f4741dd5acc7691087;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6cdf29d792a965ef52b5d693ffa2cab710eabbaa240cef737febda2353d1791b0d8e209c85b59b7077967cf205ce3288569b6991db584dd15966298abb2d4449ff8cfdf56932160a0f7795d9d8a176884ef98eed9bf99f7853647050f17114a6b1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4b2d431803979ed2b5fb699d01c68541c6eb8da3e81046282b9dceb941265eac7672b3db18384dbe3c8d1a70f1a708c31d83c84b06f668f2cfd2a81cda923677037546dd7e4fba4c1bd1fd6ca09ce9064e436dcb024c03cabdbd1a51b664ebde4c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc13a849354f401caccb53b16118794c3bee3ac75af2bca6e6d8a1ac70de0d3744c01cb71ad7afeab44d413bfc6d7a2ce3f86e27571ed52af081d790db19acf679f6ed54f2eac5acb2b058748f81e570a3c1b6a8977f90cf4578f001008246716bb7b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d43d7639ffdf7a0b7ebd817557e0ba60d5330362355f893db7202fefcecd3029be526fd29ec095e786ca5ed06250ce03d4f890c72911c96a3951794940b28272ac0d508973d336ab519150f9ec85e177d268cca419dcf5963fd4f6c6170d8042441;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd956a8db96ba275d76bfcb0e80e577485baebf4f94f45bc94c33c027447f462a9bc71b1125570fffc0932b436f26d07f73f7e84469ab9328d0a9121f18ac064381f4f8183b14c051d22fb663e5a330a1ad2b72d6684ea113cb57be4870af40f61b52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha84b706e2426e91822221d2c7f170edab78032fc9700a767df836b76bdc61a24cc8ae17d92f993d1c6915d72c8e13ddea5485e3452cefdedab9cdb130e49660c4f30fc0e3162e1a5c1294043704650ef03f9954974a9908bd75c95d27d027c67cca4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2494e01aad72e1dd2e04753d08364350f5c66f7dc695cbe7a7221159600b7379fcf78581cd0845439f4dd44fbae4aa34149506af7cb11bf8859c76deac12064c39e98861400a4e8d5c8729e1a85a4bf720e309d7c94fefe16b17a3673a5675f64c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31430ae9df8967ebb00be4c09b11cee164f7150b9498da15617af01c6b928f494a42a4536672eb8b4323278d4553ddb51245ac09b9402b5ac34a32ab4a2c03663b478b552190f0711fa7c0cff8d7b35f76027b2a541cc843a7618b368f756d25449f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71079403ffed148b0df3a2d62063cf9d546bcdb4d7df86b3115ff5416cea4a469b2087c2e5fe84d30231331f8250a3605ae8fa53cdf1302e29f5611f95f5a2ecbdea28f2a38081829ccb27f54d16cb6217141d745177936f4602dbfcd15c0ac9e0bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5aa2e8b2cc4124f6fa24ba6d8604919ed5184a4b4f9b68027a77681480076006408a27bf838a521ffc9d15cf9be76837360779ae6ed5c71da883ecbeb5ac95d52b42c7f542c52f058317e576c1114ab6340d222092bb829bcb41c83e2fe142d5feb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25dbb75233af9fbf8a6ed2c7d5f4b426df42f40a9a9362963ba8ddfe9ada3b7e6727941ddfb2d217c70d86be877b102c3acee71221506e6286955c4952ba8a1675c4cbc71eb32e0b9d4b150cabc62a6c845eb27eb3f0f2a5fcc55fe315b14b51b6cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb2231d8205f8b51543efd881930c71c19c4bc0cd85f006ed342bd5e40463affa4bf8a02d615aa4eeeeca27227615ce156841b6108d5d02d3cd4b701766197399e6569ff00d7cd9f257288746c5560056c98500a38cd5ade467e5a4679ed8865bb41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44d44b61e6c569f45968d782a64d8ae098eaaf39bd656d4e573429e3ea357af338f512aa3806d661a61a38815baf1dda0885be235f241dc174554cecc5842d1799b9fb6a9855ce4f5ae47676c624f9821b26f32068fa2908a9f33f0b000e0e8f5950;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e3fe2eb2fb8701035226281cf4c25296c552da3db001df0744a9b753ee9c4cb3dbf9566c9a0c52b838d0f0efc99c633b664d77b86cfca3cc6ab825a202f7b0a7e21f5780791b589f7af6db3b759a1d01fdb20acb10742dde9aa79816036051ddd73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16e24e8d9c9f691e2c891a9eb204ee8b2713d7710649d4cce4957053d982cae5d3ba02009c8b3f8fcc1aa229a51207ae5ec9e8e9a5302ca5f7a1b4b27e1dc99387840a669f1c7500e5315ccf06b35ac7661edd4410cb5e89d8d7ec637f67508da6b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55e82134c87b8798c808b159934db6982ec98afda2c93896ac9a1c343fb8f891cddecf7a75843a18d62115f6c5e377e32fb8e961da978cac2e5786099db7494cdbd6ba3bab5b0290736910d248f5e7a387a909176f5b7291584d12c903a12a1ec6fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc2ba813ddbbe08e3292f299e2e1bec49929df0640e48ed2e2e94f0071b020f26b689f74b7801adb79d899438cb4e7dbf5bdd0b0ada278815239dc82e42824d7b4314178ba28a4bedd92036495a062a144401b9c31d7130bf542b3ee63aa53b68a43;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb4987b65f3fb3c35ae75d5999c17a57c2db62e1c04784414a44861d775f0a1c3b9a3d955e85f3d49dd81787f8139af107023ce37e12d6b25907c9191b50c4f7ea285c8e86c1a59775b2c0d4f7f7691b3279d8e4f910f809f9783d9e1903f008e249;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd840e8a7ff5d74631d916bb974ae5081dc6bfe265ad5ca384786932e6de493d116c4e4e4077d870294bb6c1fcbe1f62134b6be2ebd6a5c684d210401966d1c27be65a92602644451c6ee5e0f64f6dce4569a032a1835164f3aadd9333ef2d4553c6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h772befac5e9b49fcc70acc821a3d51fb23b2d5789880b900b79b838cf153a5c8b23b0b473c2d2398e3271b34d6e1c2a429e5f5fcfaf504a5391cdc054235323f6190d012d1c803ca9ab0365b84910f34d094ae4627138acb2b1fbdc5987d92522c69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccb38d138050fa57213fcf70c0474683ac21970150def4db14421b96019863d99cebc42a98c015c82df78f60606db8eec5304a85b28258cc1ee62d3928ecc91e2a624ca246ff935fa79fcd7a4f414fb35ef944bc5d1adc0b5363da8e7e4b3ba17826;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he445b582c79fbbc91490802ddf5deee0c8db30c371311e029c51db05c6c4c8ae53a486300038ee7f03b666886a53a7b4915ce5a8a45ea543e9ea20eecc7f39d483aa3cb275b02377729f6e0c498a1136fee378c6015b1bc0f5bcaf8c78f9a4b99107;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bf4e8bcd708e4e3528547bfd92ac2b7057dc7ec51d97df004522f976c344eb37e1ce833417d47abd59b6dfd4e3855ce7dbeb33f647b58f7ba4b9c6194ed11e1d58f416acbc7f7e7175d02ca099534727f20771e69edc915683a25e2acbe92bf5dc0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h405ebaa57ef3660b7e3cfb4affb173b3204f94c329d97a6d24ad719c16709a660e47718fcc09d7651e575aa14bf6528fa21d96b40ca0bf87e9fd6454aad6ae0fd4220e1aaf871cc20c885ef393a602d6c420d1d38bcf648c76eea8caa100c667266;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9947dac528614e6610dab116c07adc8315c390cd85a4814bd8d2374188f890bd46f978a734fc571fd10b86096981b6f6111e19b17ece96a9a9bb72ebb080824dcad367eb44104759218a39c5478910656ef74e59d116e64ad68be934383e41fcb96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfda5ea8b3adcdcc61da23b9ca4b72324657781de279cf7c7f045c0fe5a605533f7739e30a55f50075c6e1963912d95a484fd1600cd25ec1d781b608d09eb71b64ff745c6deb8b93a426c885fe9ece374408ed6235cfca7a91c071451f0bf812c58a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfee68b2542c0893a7bff76201bfa37eca62ae8d19fe07790a06ef5e43eba3243826516e895946293fbd81290e4824f51d5da3201068858aa446168d5d6f9084e19085f2bc184cb21cd1f52b324b2fa3025fd4770e4b31ba6d9bd79c6a3a98c4ed1da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h807bb62f0f50f26bbb4e9dad6eb80bda8508726ee7288f2720128a8c010b0029a5c9ac82be5890a99f5fdd526d2339d73d5e3ae674c98e88a2b6f88c87bccb44cf7da4ebeae0387cdf7fec8732357f709d18380c8579a159ab146bccbb90fa61d32b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2fded0a88d73ceb4b40fd1200b16319fc46fd100a0412c73e50513966fc9e84e283a319faca99d4def9b04d0a6229a41ba3b96b3f631a736533c57c65c76abfee4f54888c949ab4232814a67e81e0b3222bae3d6689ddb22addb6fc8b0b61e9687f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h219d23578e9de7c9d47776344cd27f14f11d8b045a134880752672d6afa641fdbc8af044e19d3eb6c5977e7a2bfb459b30ae914c454c7ed907f928cbf55bc507d08b59c7b27eb3e57f1e3707a37301ff8628cecbfc1e83a7843b76040dc09b03a4bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21d040800a4cb13bec184ba29c1c81568cab56c0670acc890b6c53afaa4de1b427c1427f7c6e1d38bccdd8b38419df4f8382904bd3c79fec56e70ef9401cadc0276ab075beb6e81cae3227e741fb66fabefcfd5cec27ce86c37ee20797eeb8a46560;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30e8d6466c0673817659a649c7e9a548754f96073b50d3bd70c451bab2fb7325298524328bc568d9387587cf9a60ebe59b1467ab67705f4a72b6a866788f13879eae893af6d9221791d00d2dafad7daff891647544b1743e55d2ec67a2ccf7246e2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd20c08dec883878b6ed134f687c753c97b5e89682281aea63a6eee978e0781d8a27e0c19682044df40acd912295f009990bd022550ab8b7fca69141fcd810e51d285c5002d577194569db5355d1d00de8afbd6e982bdce74eec027d0689f84cfd1f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b2bb3ba648fa2ef894729875504fd547906c52daaf50d2aa4217064eb45797cb5574ec4d3931f0e2dea6439e8d1678b38155766578891694eb571fad9fe3895f562e0100297bd96b7404e2dc1b1a840e254d8212d55613911dd1836ed41f7de70c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbce35c8d29d85a9f496a8f9ed7faccffeb76df4aafe854b4d5ecab74117d1ee27983d3c071153b712aca72f05178b14f67292234ffb552cc2e10c36ad8847eddff26799a45adb0e16d2d8c40532ca002ebbe9135571d5985131b79883ef186996a78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e8682195ed13d2bd3412f557225b173e9d83e19bd6d24047df8fb60bbbcd8e25f0610da43c545df3134d32c40faf7d34ed7e5ca7b0ee36b0d9e6ec138ba2e867354d70c99aa048397823f95f5a2ff4694906008bc5765c8e55d9910e1ab9ec53a7b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c0ef8dd464a3a4bbd5a5ff9c57606c51bb2d1465aca1ccf918f58baa1361d25f7cd9c01a94237b46330bbe9ef571fcc791b007f866fcf4de83731838b9eaba84965feea1622be3949e493167cc7cf1f336b1b286fc7ee2959c83af94cb2a36ad6f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h214353cc6e532c9766026dc46796a25640e3ff9645941424f490fa0a03c6b36275ddb6f34dcee75d72c9e828e80b656ca98283f4b56935dacb7a11acb12b011eb6e5f432f768b8817bc7aa049cc0df00689775b11a3bc3705bb61d95b95b370b53b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63f6b43323d463cb682d5faac23c1dfd631f41b3bddd36b6d70d33f1e5eb6bffdab870ba0584ec9211ce3b78e867765e2c69c5791d57a3b84e711cda749f7c834ab21776045f8db4024671de95f7aac7378040954905a36616baf92b475c6d8bd20a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haee08822d261ace1733132383e4b2dcd21e1f68cb5a29e455d3de7fde61fe6612a4a00918400d0fc785a2a48dfbc7c4fd2962edf4ae0c58a129673adb065fc43eb6c0e172818a013ade8934aaba4e88e979b5daed93e3c648159ef5084c3791bc456;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f5c8e7319f941004654d2b768f7f19dbeb03571a17c8af1f2610a1a8407983c23c8e1f042e87f2c999302f3212e8daf9c8fbfa7e81f0541a58d73913751296bfb054b1d9b63016127bb5a4fc6263feded36bb1a4c77a767be38d95e5778839f1e2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a9d2541f5309314cc4b49b3a357dd88863640486ef6eeecfcf5a8327906e15b978ce11f9e6e0e6c1874c5c4f57e8acecc2393e0f829a8bed291fe57dacb81e32c0dc144b79de28f32abdb8e4e981f1d7a261ada2a745e01722b9e7b5c0ebb3d9212;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c93b1cde891b8c460585fbd547f50851aed57148cee7fc7b511ff2f96d214a45be42a1d625c90543265273d42e90a09768998f2725964a43f3c57d716823a3c477e9dafb39bcd5cb4b17335d08b087ad5d2f506e5561e09def689e3936368e65493;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h684056734bf93aa40aba8ecbf3c8207fcfd5be0c9c76cfcff395bc0f9b4922a02af3479af0e0d142fa352b443519ac977b1bb9fb1b5f3e8393e48d5b8f5f069a9a24c86568b95ebe02d5c40c5b0d5a0264f929416014c7721af9fa7de6ff6fbc8629;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h937bb052a5187f3b59a2b032eda6a9bcb71661a92f769c1aa9993bde05538863d95612ad400f902298f4a923850191dad1d6b45ecdcb5857e02cbddbee9633d20ea76c9284455249f5551c25b70188d8140adf57a613ef66f059234739e08e4a0268;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha856aa4c053b83d9eff3ec37d8fa1ee70baec108cffcca0396c556507259e2de7a7bb1c08f67279573389228d10186b2e056b600a39392ebe4425506321c87682740d3428968b811df2d3d0508482fe5772e95fdf2c74a5e0f65f4a39190baf1da7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he870766fe2b39abd5aa808fdaca5fe5219e18c20e631c25f897fb0f7c0ed25a42fbd4eb4ff6f641cf7d702c47284a9cb5f121cc95ef7a1cfc9bd05d62fe6e84e57ec9f8b639563b08a02b9d5d3da4cc2ecf86be09b5305b84934e9495f4ade24dea9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd19e23e33ecace595631b35f5f3b234717e4da9ea55eb35c27376edffbc9b744df38cd559676ac3ae3bb58c95ae36872665713f034fc88b720ca6c826e4a7d7dbd6a2df26bd2bfcafb13b674eea2b34bf4c412d062fdf97bf9f31403d05cd08a3e36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c6cedc3ccc534ac74d2f673e67ff0998532ad1107ab9026ddbafd72500608c78cf1f271418c8a6788bf009cb5c320bb4c1ef016082401bbb129919a07921544585accaeee2098ee8d4876f052047d7b45ce463bf776db75daebe77afa0a8fa4585d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdef0f62328f8633281cb37fcbbdcef0b352f586b367e17190716d95eb9a89db7d4ed46d7a992c28aa91c2f72411213af7e1cfe4b6aa0e2ec0d4e28dd72b5fa7071a2392b89f6ef770514fc7a6b95f6b2c4afe9a7b818bc80dbe186404264f4779515;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd544c1458cbf0c1a032084290c9b67308971f4eb47bbd1c83422358687c716314dded0c99bc59f2f958c1bb50d76ee96cbdddb7f48c8ca457ddedf024979513a3ed58b222ef8dc3c92b7cbcd6d937cdda7cabc01791c6b021eb43983a1833191ccf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h561ca2c6d54cf6f5188f7fc68874a92cae0b8c42396bb735278dc6bc54560099d779edb2277cc641447f722c0e659fc84cf1365534aac72c3cf141912e3536fb6321d23aac9dd9ae1fae1be89521398c4b1656562488d7a3c5313ff64406274f7918;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc89a2dae08094dc5de802ae5e34ac772007638787ca21f7a6b9ec7902cf06429a6f4df6003515c74e4fcd1ffaa5a82a29ba8705d437b3907a7cc4c80eca334f89248c1589662806f376e97d9008cdae3bc93b539c3128cca9385a7e2b1cf9040ba68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ac50be85d4b97879930fa721925b2620a10c0ea9b5545495fb22674a9ce885aca10838c0879da761d4d94092f6b0fb4153a49fd5ca621c8d901579b60bb80c923467a8d90ced98f5db158e5de0a0c690f023c1ef264f244bcfb9c50ae7b6ee12179;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3db6cae0f47c6b9a89ad645e5215550af222abf51226dadb81ed33e4127996d53db6990ad29025e799fc4d4dff02896cd7216f4c401ec1d80514764a948141cf45bcb940f643ffdab4e01e12081eb343f60fba44ecb063f8fb48f3ffc48f05b203ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab3426a7b29c729f463fb7dd46833bdb100917392c4ccfdd292300db0511c989f3147cc3c755bc50dc85f6d82707e22622dc2fafe4fb20ebb06221ff218946172d7b35a1e2d10f28d110fbbc8d8da665eaa7cce2541ef04de7841d8a6f1fef518812;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b83f11a70886db1924bccdc810619299aa5dd69f06fb66a31922abfa373872159e88a612d52e3ab0915adac88e4e211357882060d13e748c844c902dc8a1f308578048841a76338602dd4a746fe569a6fca5dd44faee333f49b8cef454874f66dc8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bef03cb7f3a8085095ca2fc2b317a56ab2f2c096db1d4d0c1798e9f9c0749793d444b86d8f5e01473b7bc2d301c7a9081c1cb8d46d8abda116af35b1b645ae074c562d617f8a0a09208494ac0b5c8e1557d8194d1240acc57d39c564946cbc2c46f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32813a2dfe2a2d82967b7da2772afc9192e4848a5ba6665c8bfdce20935aa64f1162834712a4991969f45cb2bc2a0b99d1cd5f9753da76ac998a342c4d0c48039e2c5fce9484274f67478371d320538c37c3ab0b71d6ef05e03611d8ecddbf10dd3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35415648e5e2f3e3158797cfb988ab2049584a57b90b60b6e7f62ae489cebf66f49c7c1cef082d07f0efab27f46cba548d9bd1e5668cbfeaaaba5ac10f8f5b3f9be3c574eee006e90b9cd6970079aa51cbcfdb744c1ff767f98c6d4fa4752976a185;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc15ead7f5894e8aeed348fc03b2200839492e39d183569826f94c4a40a38e84727f6ec4a201b9d56f00c3013dc876d2cd7dfcc710556c8fec6525e67aac4dfcf96f263433d28ff5338e0843215c132a47b95db58ed2304d60a7bea116cd93a1b03c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb03e79abc8e9112b7bf590ac5cc610b8d5c66fefc78a892f5aa8155a6f7f17d37e9b2033180d01cbf605d76ccf8bae40f6a2e25acac03177546b829afda08aff8a88bc678a4460889f89ca99cdda8c406974358ad5d40b2a84c3fbac3e02628cb8c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4047db543065c48e477a39702520d3ffe2f52b1e1792ed088d3bd9bba407afe85357489333ab21a93706595af9fe1cb350a4f21f8e809f0e62a49ce0863b640b4316dc0c6e402a98cfbc218e42d1618b785bc3ce41f253b8f3ad407ce6be05d4d876;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc69ccdf0d61ea107d0863b952d50f8a016fa6f0c1328ac0663a5025626be51367ddf60ea2dff49da6322c190bb169711551c70ff6f23dc6f73fe0cfb76fff8d8106df4f4248974972c3e2f15db8252a739a497e7d6267e0cd5e4501fc7f61435e757;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h715d0ff18f283a0b4a9465384cfae44ca0ecccef68e7dfd726d33e9ba076c04c7a2f4ad3c3724850c7764232b8fcec4f278d0ed76f39c6c60608ff813cb8ae07306d2ea26147a385b3926afed6edbc08435895a3d2cde7a1423dc4aac1d95df1fb57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3620ede6b90892d04ea44b235c6511d15782029f56855c9100c0828784fd6c8b625b1c5da54fd4ff36a031ed609a0fe15e72e8fb6b3b65e83e41d1fa5f6b75ef8b4d233487f6c5679ac6ee177dcefc9f5fd763c0ee88a370aee9d6df35f975a5acd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6667c7cc8f0c60e5d85fa5ac9bf6ecf333d0d5eb548527df57e79e42c979fbf8848df4e692018b4e31d7b7fee7974ed104320aad84e48181bfedb646667b12aabd3ec3d5e2b1525601401541c1335b89d9dee9d3be96f0de078c561c27ad552dbbf0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5e40112c396f906688262808dc88f4dc71c80f6165f50b2fbc4dfdb3226964b57d9d20deae13b92a6cd23ea33dddfa40650bd02e323a545027dd2018cc16c96a5330aec4e3381f46f15ac0e608deabf158e9ac2bd2cf4056719dcf96b0948c84c12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe23cba8dc47624b55856e6dece53bda0b06cbee4e20b18ba8521503bf4c9ad90cf5f58f5ec17d06eb3b7c27159ea122424290d251499c7bed16adf9ab16117edf2b8a5b609319961a9c813cdb1d671d1a88af376fb7f13be82682827b7bf9e13b8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4cd8073e57999379e16f28022e5fe447ac3ad57573cc45e827e23f03c6a7e35c704a995e9b36ee54b018f02a5a745b047d4902b589cf756d8748fb57edfe34ecd300b42c181de548bba7bb99d5ab735f5e17a0b686c64b1950e14d248bca3861e68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h708ac2a5c4b92f7f3f73e379b33ed57a0abeaa62eb9056027144f2dc8efddb1f9451d1dae645c7e494fd8bd2bec60a79cf3819d6610e3666d28f01b8a836e1136faee82294b671900c44282262765d2a05d48b73e652ddd9a58bb7abcb03a1a983a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41458d80c60b9615208d4c80daf0ba3415104bccf72ca8ff55c177a5c806ea8e6753c0f06f224f4de489c8e9d201ad6beba830a272b2ec541057da69c38c83c039b2bd45cac12b1701db43e15b44278ea3f1784945c66c1e787f942f42d7d7661924;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72d8faf62fcb19c4306cfb70679822e8a1e02ed1db9405e8f4a0f7b14f0efe753da66b020f48d4eb6059b36750242ccb91329baf3f973170611ef70746e083e6bb02b004b71aeda628b05afe5f45dc20a888797a33e44492f1e4d665ae4e7d0f3acb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8cf42a6b4f10977539897212b4c2848bc7d8dd82561592be28743c051f767b2d9036bc90713f4b81c76fe68da3a410af361e0d21449745bb18bb73cbd14ec251c2e10fe16acb6c11e3c68651de5a9530241970172fc2e881bfb4b4fc81c765f1819;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68a73970d97c8cb42943d0d591c7e3987e6bffb21524175b8075bf97dd56db7bae4080692fff607c14b9b05173953ba2905b242579668ac339814e6d5f3959e0735eb829463920d62c71d9d023bea51ae72d87e60aeb7b72bf3dff69838940b03510;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2952f3a6a033e655d4556f0d3ce6685dc048e47d7a95919c2ed9debe55a284b26c72831808b8c2592886b3c72d60aa7e2dc6b2463c264a5f3238f7535c3050df1329bceb9f7f28209de4ed8b451019a1d7dae44f358cc0634b16fbec14f208ed3ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf99386ef76cc5e4aa365bd8bf99516b5b43c5d30bf15f5f658d8eaa235389863cf86e3040e779400fb9ef7c0a4f742b128f770a052d77d2047c6c7a23c0b19ea1076a66013cf99f58f592c465510b81716dedbe56e9e2a40b429c3be1387145298c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d9d396e5cb385d5c421926f0e1248f751af832662fc46dc769cd014e107bf16fb39b36278f71fc4db6971c00602b26e3576e830fb7cd54d40a0a5653e056bf4ab46e203aab4783d200323f56b9d5cd58edddc47a60f689a8ddc0d64d792fcc94c5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74e07cb6eecb7f1c63ab2352c25326a3ac739f12ba95bd164c79bfe80b0e426255f79513e142e4a4cccd690ab5df201430b874d922bd50ae13e4b72ce5d1a3ceadd771e16785fc83e8716a051d340c2e467e420e7e8686b8444634224e7d638e3adb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a4f88b36273b8545b8523d48282a4fec2d42e2d0f52597e1292ae98dff477cd2368f05d38cbfbf095e2e4fbc29a52137f428c3d8653cb0ef3779e877ca9387fe09ba94dbb304f53454966b59726fd90e1d9777aee8e02790e89f2872c5f01657f26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44467f9847337ca3895fb4582656f1ded036b90430fb47651de53c424c6b988d9af0f4cf6eff88d292084167f7b9dc4265f93c4cd57d3536a41937bbbb2dff9364e1c68aa9ac533fff70cc9e5f7da40e07b79dc2f17a644e355831eac9ef5e1d9c54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb43108f007f46e0b4b01c3e3dc5732878ae577ac648eb3bcec2a0f4672b8118fdafcc47862024e82f5fafd334504a4cc0095a2fe1f79faf21c0c8ac8fa8d7f3751b198a2fdfbe5443487467bcd9979a7e29735b513f7a8abf75a0441bd89a9378ab6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4780e54b4eaed9df092de279c03f43e4aafa96a1759104b281826519579eeb0c8d406e02c17c2ebe826f5897ae912220b1f5b0021455a59a92cfa3285b0674182317207b8883043b01f7b871a472d3bcdc3815a4e8582f2da8d01def1df187ff2ef9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd080b9e19db16d8bb7e7367d190a55595bcc5c531feb825f6624a71cc159b595197cddce5fd18adbdeabcb9862d13e4a5439f7212f638c8d0f92409e946b8101b7075d5aaec2eb4e739644bafea9b189ce2b585a58b258982346250fc8aa881d68cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3eac08a8174a6f605f2575bb92d2c03a3935c270ef8ca372d445af135dbc1f78bedced24b498b139396e8be1cb8c7028c42021d23fcb0fbfdb43a06ea7762d2c320ccfb0b473859973c276ef9bf8d7de3eec83d9e60aa758d6d8a3671429c9b32bc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h836e66ec8456a5f0098b879039c5e8bfb018a3b55d8091f0c9b0d39664d2e00293c6c242b38613a37627a956d3a0e4f9aee65ff93413ac8e02558f319563e69c0174379eb2ce2e9beb4ca81a25732a58180fd007b0d0d7220a85c4208f963b771cf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h403f4914ac558f064a041dd98fac602bbcf5ed2b7b9b4e80b914de9bc24cd5502292e5e4be3494963db85c8d41db343fc60e13a2a0b0bfa24f77aaa82f07cedc7342efd6f0822c0fd16657c0a0ed1f7037fc8fd37cdb60fdbec3029c1eb07a5e7906;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he955af172866743c01b79b423b29ebaa1d563e7e872cb19528319a30d3abf8f10f3d23c9208a42a6d0e0c5887e2ba13078db41436b99b2b0e7b35c6ec8a7a8a221e811a165b216fabe4212036c23ee5968a8644a244b56402ef61056b57bfd433495;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b3f186ccdc7127ea7cf2773966a4674b3cc1c19dcccf8ddaa00e2162178a9b0f923ced1b46940a0538f55c195a14c20dbab1707cb37a1c6d555ad8b2b53f90cb474f4a983a4abf522eda80f5c8e2bdb8ebf3fe821c64bf3bc01cfd6d2759315e08e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cad679201cdea7a139b4370ba60f35002de09207c5f7789050b14dddc1b77fb8e8739c045f5d1e206fd7bc624b7296bd895cc3e413b94f14481b43e420d40d6eb21bf38829df1ca0be5b8504ba3e7f6fe5c5f2e5be329688f59a8d8812997c2c33c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4fe3216cd9098ecd8441a65c826c88ff01d5956b34b6d96048b62394c6612b1988b96d6e6ba2dd065f8a727bf389c702f896e59a2ba7d69c5de3dc5fd099171aecbc3283466bb37d05db3a7f4e30a4553320c8857518373b85f2b11623b7d0a8b99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8abec915b2d6b26e3f5133754b71963f6674a41b0f2b049ecaec9a3f0060178c95f9f2b3059f85c37c58c0ec6335ab8135499d9aa55bed35c23e3fafb59106131267c0c1bb308d1adeb227553dcbf1844ebe9098a1f8bfc5b7cc156a05d29009908;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87a6c992bf8610a01be5e754a4fb2e823fc2529927d16a4ec35a5fbab80a2a3d343d9af5f70114af8eabe97be386a3af6d03cf823526f3254b728041d1f2f8c9c598633d98a7eaf96cc39de8af08a396ae011ea8425b287fc1253a1956e320243715;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcefb19879b294bd5fed4488dd94f31c6e6edcdb4a7c34a9d52325bf1d5462c302a67cc8fa5f6b5e8f263b77cf83d826308b8aa40205db39da60216c6d4b3527275a6444523736747a14cf84a3f287829e79dd20c251da5ef1583658a29e48f939173;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ae356f4e9589077f8d5dddfc6500c70b71a8988f799fcc816bf07957588cc834a7c362c9d1518c40533343a4a36ac7821eb981b32eee760dbb701827bea0bd7eff2275df44b2d0ff5e81f337d5c91d2d9dd500cecddb103dc2fca6c1e22840a8702;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aae547b71cd5565f5a352b466c9b99468bb686460ee6bd4511dc2c968b4e339b6d1986e58fb06b53a0db4635712eec347eaa1f178a6f5840492c53e6d6ddab57cd0284a92911eaa4b26bdce3d341858fe2884fa68fe41bdbd5c4f0e5976620f8248;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebaf17fcbacc85d7e102b834c938f200fcc6d1667a59b9dcf3913c3f12ac9df6060dada208fcc11de0a9a542ad1a53c74b8214a7c907c6cae10a9d475e3f8e00b3075882cac584d494ee9d646b7773b557058d06b1914a72c4821431089a6a23910b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc2957f8c243360e2b5cd6e35b370e0ee2c69a8d403ce2e34d3e7a775378a9d3b22cb06c9ae16d6a9d0d19bf8c7461f4b65670e0a72341cc0d88fd17c0171c314008c606c856ed487aa487c31400c1e9c090662b4317d2177829f1040a04863b71a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb56926039ff98063efac12a7769dd15caf9818621806793305f4539f451ada1a3da58370a20b4910a4362b0e6c3fc2b302a346c296b0f4256a852b5b9c8b50f99ea1c305ef2e427344a5fde05f99ccca763a08527fd3d3be27f61c43ce5e79761297;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc49f98a60910c6637abd4cdbdb755944548f397597a4686d6df4aa4925f8d9ac93a2edbdbf42ee2278ade2d2fbe146c09552ddd036e47ba51ac6aab5995a41b8e7a216ac57b7ac4fbdae2da1f67580549c461693d6687ee0b90200c2ab0a07decea5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59202dfc39c3b8b931d1d47f11ccaf18628c1063b9f576198030db9f71c81e2f53aa4ae0e99b2c470a10e83e41f45b2e9fce1f83d7ae16a39942ed01fa39322816e0f27c84b49236ffc45467bf2f6e74b4d2a5be8d43ba435b4cbd9c3a09a2508bdb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52e40c08fcb1029bf3e1b411404507de92ed001b7c50959943a2c7225997c4d9d839f4fa97a6ef1963ff88aaa3b23ba49fbda302555807d5f464d800b37c90b5f4d3271fc91707ef242534877335edaf8be4b09c1c684a90502a0ef649111ffe95fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4579b6263f10ff123bbe76f0a1c5ab3a5203d53df0942e1eceb44df90e1b32a61e219e4a0e74fe2d5d914dd6421f40a4e04e9c1a62302faff9871cd2c07f8cddce49d1caeae33e9c73fa0a97fb6e7f9771b008a5e2598181c9aee799c633e5b704ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7e89d68fe5e25206d19cefa35219ff3c7a984f06087ceb3a8d9a177c931f85e8d8f2a9f9abd27c110d90a1231186983e63df75c2c3203ef4accc940439697d6ec2988977c2d10e54b9909f6a677b88bf1d775fb181b85334665acc74f70d9f91e79;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d255706e673583a7317102aa8df2217f9f75f479511f66b380a98234ed6202926440c09c5a7f78f4b644c806effb7811b7e101f56431daad69e6e184ec052c72864d2ce7ad266506990baaee0fb9b8dbf25fe484cf21533a2178eaf461cac0143f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce5f09708b04cc8d6e1f512f10fdfa084120f230695dbb02488763489430ece8ef4d353ac665f48a10f64a2dcc67ed28d45df0fb73603f616d30ef9e5e7749e6749b764544c13161d1fb6656e7e1e71cdcc1a96846b2fa7e4a4e2b92d55d4faa7d72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h766353b220b9962d70b699417060c2efecb3888427e4c0b4cc91d823da1d6990f288246dae14add759109e951f1c0c4964167cd7ed6b3e8c7467e219a14a14c3eab437d81a282202d042da6fe724176d06d76e623f623079454d369c0c826aa96ab3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba3cfc7b9bf13304ae36a623936b6f7088a14bb679ea49a7ad8b35689293a644e4c3c5e0b4bf6d121674ec3105de54b9d6a0f098c735f9044bde8fae895256a7b0cbcef0f51ea64ce822d6ecbdcba1f34758cc3571c01f189aad1164820ca93811db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5eb18b447ad5607177a4b62f176f807d256cf14a61b55b234c0d04a4325bd0e71d9d736ec3481080b9c5c5a76dfc12e04ab7e93eea6b1e6b8952a1a465de596e971f699385c9fc022e07aa90a6c148f2cee456ac943f82605a7565fd59c9316c39ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88aae5891160fab95f1495306691d4dfc88354e5534ded641e253e40d0273a57c2030d4e3d7921691e6c937036fd569543c725d3d62199d160023735420762b64a494d6bba6909ea6fd0b0cdcfda65f34f11e48280cd3d8b9bfadf48ed9e6d066ef7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67e6403840ad7f3990f624f8e40896b0d345423e0bbd3ed855340d72a15399fc536c9f8a498744c69237d691e901150f0abddeea733ea4dd4899ba7f8e4d28674c9b98139753363761a67e8d453f8deac46e65ebbb7819c8cb7b8fb571355044c962;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd543650688d8b978458a2f239dc3938a0e859f740ec389a56b8d48cc2d619aa3392140e75aebad817bdfe8f90ee1106c8b105a04ab1b2f3965540397ec5a94e8abb344f9de463fe2deaf0b59230e420478d77290efd0904cd1235d68abfaa369baa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8717c672ab186cf101c92a7b1a45778abb9b627886ff148bdc9ff25429ee91ca1e3c815fc1b0ca67f3b37ce0da348603c9841462bb4b7b97c176862483e3a75096fbf0f330775ab9a625917e4a9c732d92f73f9b127dc3f3b4c96166f6ef659652ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c7de820692dc5879398cb40f442ebcacf518c7c673f6b209fb6941c3025e562bd6f0178a3931e3c8342a36405489c1889e0790347fba5043c2fb7f6a60683ffb7269f17076b174636970f07a56c3338a1c759688e878fc21e4fe1d4e9c92105ddf7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59b42dc886ce953c10a00989145c889d6618dea32292b645a0ed1d40df185aba4eb875e1e366a473daefcaa3ce16479fc5c48adb271823cbdaca60cbc67ef351b0c91d0c4ebae8f376171a90cfae9181e20753bb3f5a7d004059113394ea410abd27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb68cb01b353093e86b13a6ef5359aa6eab0aebbc80c13be98fed3805d7081c7cc4de9c0eace4acb36f8a74662e9ed63f96c06ef9179cf7a77ff66534afc33e52ff94fc69708de4e1ac673b28008df069cbfa132be71ec20be032ab4549ae28ed7d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24c7603908dd1754cc1e4c065f042314ec1ffb8592cd3e216ab6445756098ad4a0887f8bec2261843902765d1712b7eb53f3aa58508b0615cfe69133e82a8998bce377e33e5f3e589d55b54b0054c59fcf37f3cb7ada2cb3ee0f817103d0593137fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a945efa1426682e1d89e2ef4da4a4bc8018eae0eafe5b8f1ffda18847a722015b05ac56700a9c9c04e4d0362c70180a3a491fae885717c7ef96472ecb4942eba99ba8b7f7325ac9ef77e62a11d48f6ddabe37216f43bac678b605a2c1f02268c6c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c26352e66ed88a69bc3032f54cba036b1012919ff94d9dcb94b8ebfe8de1e8e15d4b142035c71b6fc7a4f169cbe8401099c4dd4372c8684f03a830cebbb6409aed142615bece5055ea9f1dc06ceee7ed539f2514d5e9332156ecb2719f418a389b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fb540ea70c1a6d98cdf19cd634bb50b6e8d6abcdfdd963af96b9b5c3379bc0d187ae18e99f8a6b274c5721c04e1c970dada576614bd502fb9bd58a6efffb6319e99ddd05e14e09125998519484cfcc05e23c40396360f416eed52d3c2d139d478a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d632f427dbdd2959839396817db16328b0aa3ab332b650a1b7ad4a3b634659e6e7350f88c4c1ba889a86aa8382f9c18e3550ca81517a5472d9acfc78eeea52b48fd3ea52eab9673cd6951abfc38f2ebe5500dc12d1121a6f2d6184d1593ef605687;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h435f6467879063960466baee9c6936e6243cb81379e086519757e29b9f25318d8a7180e33519cebf7f8f5a76aaeaaf857a5336556a1aba1ae50d30c936dc2eafe6675385b5b20924762886fb2c4736161177302977bea653f6b0df978fb9aaff9d59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69ce20f5f973f106b998a1ce36064f37323c1d4c8ca5a2eb0997dadb3c94039325befba1726d63eec6503c4f2999e660bfce2c399a14a86540eebc078fdfd56c967ae3cddd66f121ac733e91cef73e1822a5ed60bc67582c527d059ed1b12cb59fee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1762811ed74aabb27938e959c7122d060cca682cd1bcdd6b9aa66f0837eec4297ba2f120610ce45d2dc7d4cf9186941b1d9a5fd5b334354f67fccf918fe921f9d3966c188d0a26ec343549fc232b5c89fd2fdbd1891ea00069771dbde83f5076bb37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8e4b213a09193fd9d1bc0b19d4df6fd0e0a5a4342550ef26005d579ec8f0e4f882de117b27e5ce96fc919d4056bee09bce362317d6a781b029fdb79aa854b61b0c99d00177281347f957a01d0671edf36000390d7998d66d79c5c91134b6177a076;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h271db5e6f34c4823118f068f0ea5b7a52ee714bc16e4c20efe171105e1c0e106e02daa2fec366ed32ac039306d8f49a4e6ea71b75aed13f8cc90e324b1f1b4ea7ce9a6ddf092e80f8fb1bc30a46a94b3dd32909fa3b42eafb10080891c96a6680157;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fd3689e5640743fd4f7bce8a3d3b4dd7e28f1b6ad037c5b6c0a7d88772300c06c2c40dce7c693ef39467c1e58cab51fa4ddd204db48c492bd78b10943c4306172ea824b7883ae6241e151248328a50dc8f0719f21128652c6b5fb649f9fa60b80d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb76f79ed103355d0406c56aa4b866b247a0918ec6ddef18391908891803938a005c77d89f9c676574ad242f76193a458109fb005c2847aaeabb008f8a1661c2769b03bc9269b0965a2b1f03cef7ba2f5f4a004b7346b67d8801892542e2a4df3b12d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h770e6a2e403cdc1e561ed02f9e59360d2d0dd0f06b72e2d3e99c69825646faecddf6194e7969ae14502610be9b4662697473f4ef72bf45d1a4fdfd9ce4022bf2657182d710744fdf14479cb75da50542ae095b34e3ee894195c16ba513fcf57ae5a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8b08a50ca18e499045e3b588da35e2d9110f7c05ad3bf2e5b31f48dae121408a013aaa3b7751f9995f3fdbe88be1c06ea3aad202a780e020cfa63fce9e19567a107c8fea15434bca00bd8524589500de413d0c1935a411c102f3a350aafd8191f3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb418fc51d55cb9e35e8f454bb7e8199560419ef18ce20077241b1cefa1025aa393f412c8458e37bb51978f9800339cc9fa62be20ace3394f4dc9cdb2339b6d9f4404558c60972c220c31a3eb3e379d87cd186cc0fb5aa44496eecdf41de81dbd7b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2619ce16a1b22ca8a7b081489aeca13b8ab4bc07aa7a2db291adc9e51c7c53c781c74d4b52b307752481c6c563c73ac904dd1511ad922792c5a7fc9716050c5f267c948678bf6175bbd206e1ca9f6a638ba044838248504e8cd1296962ef4a36bae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bc9f8dd322508249610e576cc5703f96b57b94e1cf1474efb459b3b098dcb1399af92037554bcd7640ed491d089e6929f4a17e2fa7ef81ac2c1564b684fea9a7b5d79b41c603f5b798e4b6cfaa61ed42389f0e676adbe5ad4cbb56ba9237b1e4ae7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd45f3e5023e6e867474d71b484e538b141cd01fa02e75733835c0a424e02c220521d7c9c27559a1494284d8e75db63ac7464b47dec00775f051d3545fdb543f7ff8995c99162c75d1f776d6eebc59652e73ffa059604c483f1c285a647991f90d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfaba148198d186df25253e8c66e28765c8ffdeb489a2b1214b75939781f3a80cbac24328c85970f98b5e487c45ad2b36fb1e74bbef99b7867cdfb9285fdb6c66822e08ea5de401beb93043de7d3551f1ddf41c6c3d18de5df965676a6850f5b8c04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ade28144e0bad1629bf63105817e095419146074373f6c5c52ba016542108174497d759eccf6527965defa1752be18a7def8560ef38abd8c71df37125b2b786b984c76f88ca31cf76c8c568b50e1c06524bf2f0811932a16773c5aa6c7403059f90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e47dc31dec02b00688c1f83c94632914ee49e46685e8221f55e0da4e4f32b2292579f73e171de46c6750207f437348b5445d02ccabe609f577b1c9101be5599b7b04765069959081b9bf1c9e5928628c7ecadf0e80accda63f13c0c3ca2f398c5f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d6ac79aa5d448615d676af544dbd23c851cdf5b91c54ce7e6f2a531de8618c5ad3b19afa30a87c73223e8ee51e11495805e6e007d6e8b4da4f86313d07b4bfbbc54fcaa9cff7ca412fe0893717102666a2d07aea3b7f7d595642a7bb05300ad796b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h996d0767977e3678078018e2c19009cd5e4bc805293c24b33c39b9b3aa630a8b126987e4ab93eec3e6715d36f7af7fd8d001f5d2d9f70da5a968d373f723566c132076628cdc6b32eade802c94cdf9143358f4e2d61be73aadd6d3ca0c4168799a21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4963c003f06f57005dc53677dfaa1d7dbefea2c2b433ce1ac752cabe296ceca237aaf63398e4ea274bb2e9517a99e078828badebe217e5bbdef1cfc19155bf4b609ab5c70c41544b852ccf565a2ae3ae417e779d9cfc57441bf550d6671fc22f96eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc579a47f5af10c9aa817fafd48f3686faa71de5d31790eb492f455df81e875e9a1cfac0ffd7ad80251f74f0529fdec563aa82d8547b8392ddfcc8219f3df63e5add5266f294666c81165a1403dd4e6e8ce509f9ce82394c3d02dd5616395bc3ac44b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ef7d345789c9a604f3e1e5ff07847cf18757ea84d0101da02f7719ac2beb2e3427a416a9db08e1c9b1b740ad4ce28167215b2c9980381237f86d21ae5e3154b70b3a52127d23bde04899b49c407410f2677f97d24803c617cc2b3d7b2fcf90b9f51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21d5e0ee8dfcab57126c89e376af225b592d807b1fd8ccd0477c474b03dd6e920396d37f1e506a5b13987521b2720abc02d0b1ee6bb2bc14e20023ee89bdce059d3a29d4951517a8d06eccf75bae6f45f40a2dc71e09d1807e7eda046aea8f9d622f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93c3c520712452856744cf6c8f3b06217590abb1f6e05f8b3a2917a877de0466b65b6cb54977121f2b15fe5901713b5ed30fe61463c5ce415d6f5a1e6ff507c1dabca109ccf4cf958d31b2c2097b98fb47b47b99bd3874ab8e60bc11879edd320ae9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4a7c8bc6c2244e4efb70df1aded6f7584b41ffb02e52bd5119e83258cf303d5323334c86f23ea496e2fcb705713f4d4afd3a3b8d24c45f600b0b7b41d2731a15890a08fc63cfd2b586999f977180311de0a4648fca2698a35d096b5a69d2406e88e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24039c68d73dd162ac8c16745cc4f31e90fed43f9c1a3157391a88838f45011adfb2647c73e190a09fca42240d1a12cc452c1d61827bd1f462ea38c51b964624e36bdab2df87a780d5ba06c1c4e4206256447525e6f664c044dde6613464c5dbf057;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf70c4e5e459242775c0ff09e9236d286f4e036799eb12cbc4aadaeecd80d7b1981946118a9b3d68588edf3def1156129a9b3bbfb70e37330f6d5858ad02c4f4907516c0ca5bc1aa96734777c10f459651b307765ca11db3531f969fa55f2fe8ed56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff77818c3c311d171461dd8332a73f9cdae0c1caea6e8a00f0c7eadc1b16f814e0efe4898fcd1da3b0c9e3d5bfb5c6b7092be6ba8d66babb9672522fb2a84a02cf3aa988be8c64afe2f8e15ed8bd1fefa5f403dd0d1038756d57a490c87acbadb00a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c1ed4c3e660b37f5fa339dabe0f23934e92c2ef85589e7d5a6a761256638337b968a6bdfd33092d2ac5827676e8d6ba519b943eaab3d9b0a9c8debe8aef360533897dd62ff7653f12038d02bec2d602b4c9f6314136be21ea48b1ea7a312a4d64aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cefbf98ef0697908765933253995172189d1afd59c39702fd8058ee7d064f1db023e10da784ad815f95b6b292505e80c141a792d83a68201254b4441cceb6cd4cef8eb1ea8a5c4cf10550a047c48542a47ff883f72919403cbf7842ed23b479ce17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fa5877467e96f25b6660c773fc4ae69ddc4420094c4ea1dc881f45ee8fcb500295b7d4df6488ee7e4b8915098bf081b57a7170b07b93aa55f62e0ee524de29a3c47449bb0e7a7ccdf809871b74a0f575031c455ac6c3ecbdcf79206159a0eebb9b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he85c1bc1397f4dafeccba3c5f86ef722ea5308c5f400f698ba7e385b90651d6cdc60e2f116c051dcea90d14d88fe5e10b207658a3fd2eb03ca68cb1a59dc93e420e0bd97ed43b15cee2e03a09ac23ccc5514a3390137045558c4d97c34afab08c172;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a12422d2a2c4119befa0334ba78222b20262112c7d649d46e5ad069efb565db4326ed3a01cbaf6af6454ca2f74c1d985204d86defe71388c62c9f4a9709e01cb02b028c0546ad73cdb1a0e818c79ca2c2c61299063d1f339b4515d4a86d32f54cc5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf165d3ace5a3077a5bbd22a3edfc2920ae901e834108502fda8ab91535e355cc6772930c51f3122ae99d6bf72e4a4808cddb4242b9d1b5e150fb9477a21f0e5a18df756403ac8c073c18c336a5c691b40135b67c311f2da2f198b21ffd7b20b0d1d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62b31445ba096626e95a5a1f22f99c32ff62947aeb4c6cc9d6e1f8af864fe050aa93966c0cbebab22879586358b423e6a82988ff855d3f6d8a93b74083491f7a3bb9556990cfe84786056f049b1a90eaec0f418fc95749cfa4fe640618e19bb2a0e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h152c9d5e3b010c59fdc61798a792d1f9981c0c8ee7e00954117688868605e6a166283efd951f1b06ff004eabb9e5942ec375b85bcef51ca2b58060414ee779153c822f92439c35d1f2f68d2536c92c3ee6e4a3e482f3cd8ead73531522fb5d7e6052;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee27baa854c1ca7de4a4566eee3c886d307954f8100081f63b237eeefaadb75d77c789abb5c2d570d36d6014ac520be91a5fffbdeaa8ff1ccfd44deba6dcb7162ec039c4fafc91bb76860c14602d49d1f99369e8fcbc61097c9dad3f9d1a1a0ad943;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8f0e09ee6d58fe9826919e197387a9367a63eb2fdfefbe36805d1076dafd183a4ff98b25220dbfb5a7965d8e51e579ed290a37e8def7222a49355a856e55864333b596dfa86e57c4563af4119f1369787bb33883ffee979148bad29ed46fd2b7b8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77f165f5cac81db6bc2498885aeeead41106a367bbd8f9bf9fdde1409efc2acb7d0ccc2a0d1aebd67b1753bed84e685899e966dcc9d61dcdec7abd1976b522f57b6afd40672f6e83917bccdfbdbef1dfc95375920f957ee9af6a1a130dcf8a5b7a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfca1a56c30f7f95ca8edcdd09657a0fae35c8c043a68363ff5bc411c93f1d10f642db9f77b1662a5679b48f1ea2d2a13e12271ae582bedfd62f326a53ab524c15c16323d79987276d5ed3a30022502e0b31def469152dc16391ff8d5e09475a1f60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d9a502b67154a7a6597bd60538837b00de4bbc43151059fa5d9eb52e514d41bc15ff939882d60adea9027217e33b1b343098023ee734a049f590a75d028128db110fd067b4156dca196874768911e863b42626b904b0692b6f7fe386cce9264714c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2dc2452d071118a44b94b7acf9fcb13f28a80d1a468203e2eeac4f2d693ad461d92ed5c3853bee6a8c4581d8492b5ee479fe2b38c54363a6101af0fdf86045a1a1c5308c5191e6ebd96affd7bf157caeadd5749874ee7f0dd5566e92d789e7091ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cf46b83a8e3b2637895d6f4ed48daf7c04acef7567023cda5fcc6f3be50d16c53624107e004b7610af1d3fc0d865dd725e9d87ac8b5e4a9e4b15b4af4c784b57d1b67b0454b70597defc1b3ef6992085eac98e7229dabfc49da8da1cf333acf2a85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5134c2929ae9a6ab50bdeb9b83b7e19b162727660fcc19676b834c4e91463058b717fb830ee3813b57e24196407935d7c68b669d5c1a640922edb8c8e57dddaff9e0f06c51800473ee2bf0b3a43b175017b4f4857f7d00c95be92a3566e27ad6d3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1c0ebf05c52a0a2fdeceb5cf021490b8407f2ebc2fee898199ceec411a00fe95d3489293a717470c32b97e4f65142d8bbe69521241568e1d1fff76120ac00fe82022a0d6eeab3b70e5e031521e3cae4f7a0d4dd0c3713f5069503dee3030b497bc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a39bffed5efa816f51089c46134f0f1d1d94f0de96051ef16d3b654cd4c54a6f436ac8e0897e88d907d0475c3f71ac18d2f4b76a8b1e59556203cc8ed795e92b86954fb6e7238de795191afa97dcd33bf231bd85000efb52f4dd670a2be472b30e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h117214ec78eca3ecc8aafd244bab7bb7ed5e0636a61cd834199dddd5e56a9b3b7574b0d9dfd42aaa2cd011d79c29cba24eb7efe312b4c338c2b553625e1f69d9d0dc3e12ccb28630e124e869fdd1dc972bd628af67612d680f5d5e6af8b172f8a717;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf08acd4b9412478473f2de049753b28bc3d2b1b36c2dce848cbd2b21cc52aa20a118d52dc42b87a89ef87d14a57a916c09962aba29eba7a636740da7c0775524f43898b58d138b606968b762bc9c6a5a6659dd085027e9f27fbe90a050048afd8fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde5b30cfdfcdc7bf23fc4be11f936b78ff788756f2a05248fbd712005a88c536a143480dcc89d175fe545d0c3f00083b4cb6d5dc67db50121716517d4e29142198904a1aadb6311a0e2f3cd960a3b4c1742e5d0a454cf1d69bd0e0872dfb1a93150c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aff56c1fc6c748e9b518b336ff3f5d185f6b32d9db0c82e8d8914d552713ce5a6b57f2d7cedfbd7f21cad109cb9d949144f275e0bdce9cb3edcd20d712d6b2383a3ea04f7a81a07856c885b1e5cfa872bed71c43f48b2048f5147235d9ff6be09d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4ef91c44eb20ac5f8dfbe2ececea787c395b9471ebe23248872572f489ae507780c4702b2c0be1d0859dccb0c576575c6c277edcafc73030acecab247da5cb323db7d172203a9268b9509b329fce04d099cd7b5d39a535fcc6e0de75be83226068e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd00345da26390fcff7f620c516c305ca89209e838eb40aa10a4072cdd9e1c71a89b13bff03b5a962850ac567ebccf9754ed983073de828c6996950f675e29d33c0f9789792ffeec3e17c9cde93466849f56d8d727da174d4b385094c55f42ce287e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35b1fc9f0d3207c1de55e40d00f2fdb28740075e1dadcf4377912efc6eff854ede8d6fcc921234a64efdaf79e7775cee059acf3ae55d338ddbe6b1a318f162c3998b0752bb93862003cf21b4045407757dbcd5107392df1451236e0421b0611dc23f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9981b6eb93a2351cbc7b1e95a2aeb82ea7c663b9d11851c25b028bb9054dc7badd9b095218f0ba6c8fb7940174be34601fffccf10a097e59e1e3b55d48e81ba99ad88f429bdb8620186123330e3f896ca3748ae255f4293e99368aff4df7cf57aa15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6425ee36b92f16430e6c02a0360ada11f103eb0fec3bff425e0f9f07d98a48769ac2a0adc393958cc3ffa7ff0bd31177bc236d55b7a3e195a54fc3b6bfc03758e18f4b97afe48eb89341598a63fde8a494520959256bc160ac0b417aabe852b7423c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc439d438f7b9b00f033a5ce9372c6af9669e119373bd9da0b0d0c49f10ed406e45e66c4d509bb654d35648060781f889057b0045ef38ec23ed608681d5af52ee58c569fe6312f8fad480ff0f485acc0d6bce22ae535ad3f4b02c78a49e166fb7e6cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4063eeee524700feb5bf517697f7bf2d3bfede8f7ecb782c4db4245c1f513fc7d5f25d3bc7de46abf68e44432ae554cb7591127b59548d5705407b417673792fe25ed28d68016ffe860ea2891d0fb5d8b69b343877b3a3af789dde66f3aba2fbdc5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h699a7140537a91e8230eaa113ff843f60f781bfdbc9e5f96e83fac83105816236cca9bcd20f3dfd03e70cb49d2f90b8f207bc147e3f58d916cad5ba57753dc3c27a4cd0c0e29337fe6a7fe0b5b54eb422e66413ddede002b098af0ea3760fa065aaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80678c7e213e0dbbd853e217ddfb0b72c6e8fadc682e4783ce67e40f1548ee66f8bb677c23deb6d2608f414c354d1af1031d9322f4c23dff2f03b9ade1f5a8b56c80c233623527fefe0286d6a4239cb18da01d8de6e9229770bb153fd36c35a6f2f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf906c7f3afedd2f0567ee17c74a3d78b4830792cd104162f4dc4ddf7543b82482f900496f91abf8b913b7807070c9e371ea0f3305c7f3e2ef4296ba4224f3f37a02d60cc4e0110215e8d68542e92bb3cd4c0b010701e73bd788471ac195c068d3bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78268ab543e5c923a003b8c19ff9b24f477cae352d51d8435f6277de11759973706150e41fc3b2cb2e6dc1d5876151090cc6c330cfc5423392bc50b093cc8c66a5eab6e85d12f3b6f69c7274f53bb77534ec553af5e194df51704f914e2758b596dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72ae31d3b418d46d394f5d24157736288db4d551d2402143e2fa24014235ea1f48fddaa83c5f130f61edd1ed1c62df86e9a9dc20fe281d0cf5a0834c53af96ea7990f526a6c185d23f8d1ba5e9b7951dc5ef45d049f262643ca7cbb9c13d46a19779;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a1a9c66dfed77c7fbc3190159c6ed646bd58430401f6471db4d2e49d452ab010bddda590706464d2b597f4d1c80ba279b8390c55e506bb257191cb38feb24f30c53fbcbae973090a2f5d2569b90f05ef4a3d3b58e5f7d2fc2415e8b304c81aa684;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h487e042198ae46c2853e8a8a64944ea0e6a108e4fa46d50e23995b3ebefff396123f4f48dc9046d413d000d06a161dcf4087e1e1b618b2e580bb43c830abf6ecdb7aecd4c5c1d18ec3842c15b0cd070bc7c860609954c99b50fc04daa344f285705d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd78832a330c20198df7b9c236f87bb4c9907766309aae1fb255abda40420575db0f261ea7ab123f2db43e5ff2cd1ce83be132c359927483956558f3af4cfa419228b147fa432e443cc48e555414af5bd5a4a83cc069e514e99af23e15acec683fddb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62384542fd73b778ce32030e73bfb9d1d94ac1af28a5f30bc8c6dd6200d46a8de25c56a5c2913da15acac424e9fd602c86f5200e64ba234fbfc4a588ee421049c79cb21ce5cffe9a45c928591177ee639eabad444f99a1330fa32e97f88563f4378d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf34cc90f661927f5abc58c3f2ab35005a02a21f47edf6422b8db49476bf80005102d232edc5c1baa86f86ddf53aa5f82e4163accc5afe7b8836ece4c08a0739690e579860ab7b8e2e79a4604a851ee24d7c46070d5e56e364d9f94f2a5ba5941c39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd56a937172f73ea48696e89141036d958db243a1ec1f100defa404b953dca9fff2adeba73bb24adfae6cc84cf670f875cacd63fe172b07f56a75415d31a8f42eeabe9e745696c9cb55c2fc978a340f4f6713a29e2833b1dfc7d73e2847fdb38e5185;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h657047bf2800cd2995c4e42b30dcc8bbf253ae49da06897dfbe768da296a71bfeb8c6fb60e19b3252df0627073514981175b153a47e7ab517a00330c8081017b4f1e53d927ba9af0bde3c82014c9ea13f86bc0501aca2f8babdc8228a2836efa491b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70f71a6c2120181f24d647d5399d5755f9141f2c5e0c515446d25bf16a3803147367c16361ad823ec3b2d473aa899e053b9113885354c451285652a821312b7382dbd1541a57f8f5eb90a8c2c0c6e95a035730f3728772bb7cd238b96933fd35c158;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27c90f1f4b2c9117a283084992d54e24a62b4b97d7b6ae598020b25835ea2a632cec0e982c3a9752603ad5cb4bbb985e1cecd45b41d325042143b3e44b76cacb6bc53e7cddabc7c9a7f7aebe4f08126178febddaf1b0578e6cd72abffdc3429eb268;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a39025e303c443dddded8799c9a509becc6845ebc8137f4b6873a6295462c6766e205fa717250d374ccef8083861d190c8c224688f7d6d93ac59e415ca8064f05795257a88dea9a4ba56f7b806cebbc51f1987486e3942f1a5a20e6bfccfcce1f36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf79b241ed3f6d6854f317bea0138a8fdec00383d956f269e0b471adab66962a1182cf40ef34034b2742ff3a1ab5ec132af14a95277de2517bbd97ac67a895edac28a4151b1964eb4422365ef7984ba42acb7576ef0d2c4658dac624b3afb55f7cdf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6857d410bd15dd8a98fe84954e8e5e26319315ab17a1c96dd403362ef6edd2bf7dc69222877ff70ef0c200990e019b7874592e1a8e9761a9491241dd606db0ef52866a704edd3461aa704b7cbb3438f2880e9c5aa17a9ef44da3e3fd0f07258ee6bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1552d977e8a336292a211f0316f09c83d234ad2d45fa996b3d8e180670d27ed2f6b425fa913bc6b5b2c8aea9c537c5462063d45cf296b8cccc31086b2e92bf4d7994e0fff0475f735fc340042a8b4efeeaf93bce44e03dc1684449f914a658d7cbfd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc91a915ccdeb0c8a64ddd1d4d50d0a497f92d131950b790e0ddfbb3814be9c4ba4c1399b97233669c268ab39917fa92977018a791a7c60f3485e767c8e625a605b226957d9ac78d2f0c86ca413530c0b45413db5a92ba35f35679e4f4c9bea215e53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd44628143bfffe9b7b559edb0d6e2e9f78655c9cfc05f89e3d58fd47e215b469f4b05972528d8d5f01d5183fe4ece977ecb15a963ac78c979b2ea8b2d267f82ac8a65db2f6d1a85cdaa22ec3b04d3682a0c7cc5207994c8110e9bae5da2f300a2032;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddfa64f8a040acc87183200129a929114f9acb798d35338161461463e272e0e9ca0b69e02c290d7f8ee648e509a81589195bd1177758d22ec4b0f3bf35d1a94512f9ff95bf810c1d06bc8a33b8ed572306c90ae4966dd65075b9029a564f15e07557;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6149b753f8f58de771c5f39df52107d0c31aaafeabadc1a1968a364b54ab3cc92628c69d14857a53163f0c0955639a44da3eec8bcdd76c297dc5723759f497300762c45b567e0f2abd461e844a56d67dc0923316623e8bfed3f4d9a6d6b0c43f71e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e33f912c23b1bf9c0e56df8541c3d737bf79283e6171f7b917e1c400a10d2e688dab3bbeb7346871a853ef8cd6c848643da0ddfdaa6853e202b3990eed4ee9b51f652296595ed257e6a3848182f66f048ad61b40a2dea3b61cb296919999dc5f964;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b182f5da161adc74bdceabd4de15e3d281dabf98723bae0a865dc8701c4bf2d22ac0045bfb8fae484ed4da13b5f06c9af3ae549015df0cbfd64db385b1d67ec6346259dca33aa5273246145508d4f3b4409461334a84f010fd41069ee90e68c6949;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h732d3dc73a27b1619c757ef1fa95b7de3ed5e9142828b3d0a6a21cde2295e78941852fa99fb14bc83736893a4253bcebda20a47e54edd604113941d137597529eb1ea6f038a6f59b4467636db325944746d298580077971246554e0bb3b17ab77385;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0cb40622ddfd264f2d0a25f6b53e2373fbc6a675359984b4628d471f1bc49675f89406ff9cd090a4c284f58b59dd46b75dbfa6d043da445f5538f923a31a4b5ba485db453c4b6edcc71c643073af2f63475a4fa3cb2984c507d5090ba343e0afe65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb080cceeb852821ee77e4bca0a5a9dd21826eb1dbdb634480adf3268809b5dbf8169730d793415d740829841474cc47f4eb9b9149624ae75349f1b2f85f0e998daa09dde81d8696be94e7905eb40e1fb9793a9c9f5bea155280c0295adc1bcec54e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77480b210aa1fa9d0834be7dd0100da261a4de50423320476110ea83e278510efa5ee439cf5c3686feec64006d77a4f8c761fc4a9aa4878d587dbbaab21884d6a1c8a3ff5c569f2bd27d672625c2b9915d9c84260ccf59aab09a077592f7315806f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf34512300b1bb0cdecf383da62e3a159877c904a843cc20feba412e0d6aa046fb8fb0f1fa24712803474c48f61834e05e96cdb458e23bf367d17e4d51790f424545b88534993e715d3e812f42d8988450418fea33e793b76366cb6a9c84176c69257;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce830a832bfe7f5b05eebe41bd9089ade1c97fef1c3ea63c344a5f6c3ed58cce6ad5357fc05cd07f8a0c0d2b4fcd9cc353035d246c5af4369a1e6096f4599e0fbf614bdfdfa174a6779eea247c197f7baa90a0ed5c679ef23c0396831f2c8e2e7b1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0a17c8d29455275754f69069c0f73123a111d4053c5d8cda21374f3fffea37cb27b4b1f0de7bc2f85f559f08175cb44a74f5f7b5d6d274a4b483947b979e60f4b03198aef3542fcde4f9d2a21b45537db094a3e4a9b4f72548623d7eff1b639c6bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49d15bf86f0d4f83f98c61c817bdd5a9226b14544f5bda677107aa078bc8ada74ccd8d2e4bbd876f2801b1b136e1f51c278f3c444c97c16216b8a533695c1eef0c094b14e553bd6c7c1abd45cb15533116285db7519cb1b1637071343db78b050620;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5351c8e1290b73e83eb01b6e66ddfd081607e229c124dcdf54e7cebb66bdce10a197742eda57d51e8856ca62ee8224a1dbda970cdf07b39bd58fd4b8d069d028728cce965652511b62f6c705fb58eb4ab3aad15a8a64acee57f88419b17b006db66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbe6822bf4d8c5aaed983d3e577a928221fe2f84391e046e144f55c2608c1e6477b39be2d0bd573d04e3556a2778ead00b00542d3022333fae3fb79731c2312c999ed15bbf3d935067326fdd829bc1ba030f5267c3943e34ff0ba5de23267d611f85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8417be7876906d26f84d859d57f617d29cfb8c810fb4db1d5c90abe88f9ff7cb3befe0f27b8609f519d7b6be3921d017c26bee210f552f9d236a5f0edc8be09e7fcfafddc60318e987600aad8ef3fe2f2ea1316946a7900328b19db6ae8fe2c6106;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1719d0da934b9e8bf0529f416e6ccad84f1c1a7c8faf7cfa17c5a8fd09b576e32a18030918da6d31ddf19f7a9e6a134babc3cdc2274952aae6289603a030d6660734277621a43c76a10fe42030fe2ba67538b5c037e82b6760419e75ac25afb8c0c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h168f00dfbed7e1dddc64f337e88affbdad110fe7d38c3b94a2d38c71959cb0b414d6be2002a25937f5333a3c29f96522fff26e9d198b7428e8135245854591c0e2b915bc4d03e6c6ed4279010209b932d3d1a84ddd035eb4d672f8b3c3cfab993d8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a5951e0723fbc6d3ac174b5ec66e2196f1d36f02bc47ff366254b572db8c310a58b261de0848af6800f00594c78615b8bee275ef1c78775a02815275c87bade82af885502da8c2a16e3da62abf4c042827089916d6a56e9b0c2a0b51e4b007211de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4de9f420302bc8e9b5ee9bfcd6a6d4440f867c612e5fb22c978f8a7aa55371f4fca13f40151c9263abad749d1a738dbea397cc6152214400e5ccd382f3149c9428b97e490226fecd8f302341e6d13f06cbb72f5417aefbca4380692cb7a2dd6a7606;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebb6a790b3a639501d6f4bb90317ba518ec3d85f40253ce3ad8f4cd2d7ee47864234d4c5f21efcbb1728445e08983f308deb780af5ad5be5e22e0a75390457af0bde5da06fb20de9ed862e8be48d1d4b66262beec2841016915cfde47e42154c67ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cc22ec2f5e8fe34fd8d2da0c89ecd64831c934a3afcb2db06e464b33fe88af1dd9f2ae16e7c7306b40fb61a404638db141e14ec7af84311d5b22fc32d3abdfb6e089fd94f311385c400f1df00fff7b71f3b133f4dcaa661dba8f310990a285c7b89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67476e2a184ea7f508e266eb2a9f0cd644f0c521c9dbc92636d465e88e4469a2d53ae6d9cc04b2780d6ca5c8613c067abbcaf8f4f4ec2b17266893c8ce46f6ad3bd28936372e1b6b2a8f27857acb6e11e01733e9d44d87036b72a87a468c35c22d44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a33837d1fc49ce38bf1c612a83abca0fb0a82dc8e4e2a0059e5115858a467983dc09796fd740e738d5e7745da54c73d14c85c0706e638ea3137649077c93fb171c5325248e76024af77c25861337cebcb3d735ed0a11525b2c6c5542a2960a397d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e3354389622037264986138e0896925a6eecc31d29a9a86ce00be004450a09fc3ddb22fb46ec5fc564be563316350ab37fceb90ecf72c2bc716dd216e4c6933ad3d9253efc41578df8b8fa5a79618d6a8021666586039d6264538f00dd385d6a965;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5308956583c1e3b1c06456ea2af6c7264713618d8ec5ad0f042df42d75fd3baac829a24e03c648428c2b5f35e9c09c01e430842ee201d6b2789420aa4aff8848b6fbddd87abff36b7b2527e098f7a25edca46db57e9d5dd5740c4ea561be1f43f55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h792818c4c0f208c40fe200dd163c730e870b525d866a73d571a913b4f765e36dd692cb7a5efc38dd838b7872fc488b3bf33d7e197d50701b3f57f2e304212be0cf74aa8e6184ca5d6ff319be051223a8c4535ce8606a9c72289b01937d5d207832fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53aecd32a59dc9bb9bd396bb5cb3fb503796745cac796068ec014a2ff8e79b05cf3e9ec5944c070056eab3ad7f5231eade4254034fbe6c376d32e88c416189c153763b7535587c0235c16479e7276692f0f88e3238fa355872fc5819f6eaf27eac3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3fd04ac7f0d1a21fe3c07a4281828f5ede52e5f7c4a352c4684ae43e0e7d5a721d8eccbb0903a7d5837134c0a0fc427cad927ae9acf6539d2840dc732f058626927b1257ee801886d1f1d15e3c57adf97e9b5a1382e2cd6a2c0d85c3f7de80af326;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab61882352d4e4852bc16e2c7d0c17985170ee3ecede6f31cac85672f87f874845457ce12c10208629396e93a1fd8e1d43d3447ffa50167ab4ec5a11ca49dfe97541b350a01e7b0b44ae70cd35ce0755061d03311429835c157a11c64deb05d3bf9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2782b4483c0abd5c5483813747019628cecaf9956978154a393834f484088911000a67c3e70a791f71f0f6344727f3de0770f6964c36443a15174d8de2c2d9242859ada2c73213549c500bbf5a68e3ad627d6133978a0cd8fda2fbe48c29dd39aaea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcaad135833ee40e8585ea9c8d1e64786b5a61e5afb8e322317f86534d760941f0c598bf5a058da01d9633557bc206ee6d5741ebf5711b200ff4f88a0aca864341dfa5774735c23283ed6be6994f0d10805fc0f851dbbea0e834af75045c5a0baef07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd353c76e970521ea196702ee7585856694fb58e68062c7dfca4b5c2846dd353ab34afdeb0219f04929ec8eca24d76996ac7641b89e588d5bf9b5a83400a491a001e67c6526feba16f5d78b7d63775963fd1989ce3cafe21465d8e3db7e596bf5d7d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a8c165e74eccefcbf2e2bd8bdb9fe3449545efe4a00c722f34d2eed02d5e0cc329c5b355f0fc1160fe0598bd3e89ed072a206597938f6ad5a8c2a44f7b143c2e6c0fb435d7cf77e0b9cfda921b370c42cfac3506036dc965c36a70c34f980e1eb3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6af631ed72c3b15708f22fdd3807ae78256dd5cc9476347714f26cba0b8d0277126d37ccd9c09c2e77784a900acb721baa1c7083032e053a6cea5a095e4d0ea192a52709c57992b6a5d95a1aaf6204a12a560849b5a80f3ca2abd403ff953e1d8722;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4c0caafd375fcbf0920936ec2da3ec41cd2db53c50c58387bf7218180d260b71ac6eb3b2e546204b36a9fdc28dcc104d9583a5294a6218bd61acf611d69cad6e65d2b3148e95b0dcd86c6a23d74729c6ff56821d9a044ec1b874002b22babea98cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2eff27df2d3ab3656f43405a3b2572cf8a5b2642f5d6df9af6ae34a9532a4f9324ded2a59fca76f6831721c5e2b65ba82e3290044b477754b20a8e98da752e3543f79262c689cada50d5861a2016fed61b684a8ff6dd8aa2071f1fa7d342d882da9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4f7810c6c0f6f0ad7c3d51d2ccc41ca965966c74d9ef75be89e3b8cc5366adad80d81eea0e6f75646e66d8c17c879a6674e3a19af0538b9bc65e827f3ef689f1da2f1fae9b201c1913038d3d72ab541238a7a218c2b1b69745245d7fe4a60b260ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa4b81f9544e48a98de904256be95f2dcdbf646f9801c13bcd47a5474df16f9691974e7dd5eed6b6075af25f21791fb97d31c0f73d91ff148afe2ab9f8d4dc067821d6310f4f84a7c988bcc04224ac56649142b2beec4923847c468cc0f03d5bad30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27a06d8a1203c581e1254d4748b2f814ee285f2588aad3c7f500d3068dd6a2c6c0d9aeff472204fc7870d0e77e108dba211f9f1e693600f8e593826d439459e3452e41ed8e0d69fa18e72fcd7618c123476c6abb925a0612d4abc7d9fe489fb740ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h989585f665c8458e9825399d72032a664cc78fb0a1ec456acc316207c423018a4a0de4e413122f40b409ee59b72b797157f7ab9f174b64065bc182b3f453e79f328207f719099ab681b963fbb048477ad2c13931074ffa3cac680628540f7bca7303;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5edd9b7b64e6523784905ad33abd0338c8aacb942ad41b9e084b569d22a93a91a4eede54af91407f76dc9a9a0d169e05f4c97db96e2eb3f97ca68d6502bdcb653dc897c331c7e77b749e4706e8c8003bee8b0410bfb17362da5ea5f05141cf41347;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2137d4bc550391492a5732c2b785d49f42b73e5501291ffc50d191fa9b08f3d9e49710034fc13b53cda945c656a70639aaa707fc9809bf79973293a558e4feb88d3d39db975ea6ec8399e72784f7f1176e5bca42506119a02a48261df13b03fd13f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbee9925d9f5a35b905604e9b52a7965ad4ece1c291f0246f83c335bd4954c64a14e43c8074fe9680383bf34e2198add9c4d91748c5bdf4a926ef9313d4cd00f4dce52e59099b220b5622abd7ad6516aaeea732f4386c52a668249f0591a274e7aaed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb727e877b77dc147f17af1ff16c7a40581375b94a058ee58155eee6072b5ccf95064df02a0dbd25784884886c502163fad4871b8218ad5f4b363d8f7a190db7f61f8321a1ea807ee179e9079562bac36884c59103004ab8353bed01e32d5f52fc608;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h689b48ec55a3a9e1ff22d7f61a6b286cb42b43b30a64cffb16e33c3a4f4c23df2fac2914986f676fe9978d51d699c2735c2901cd7f9ac4f87f4be9613055d549c2547d90281a1af5e4da5f0c0ffcb7c0182234c117410074091152039d23d19d90d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e624698da49fd033d44e6f6726fa130b12205a057ce2d161f74c8d212cafab797f79fbc66f116ea019b7bcb2ed0a4214f7d5efb66dc7e8a9e401591dbc39610d0de118d9f0ead1a96b5d228de75397cfbafbaf12f10981bfce94bacc3854daa99e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce99ed27045dd3443fa9035ee191d2dfec2d16631d6e635914a412e4402a19884d99e719a69ca591558221713ddca9650287cae18a3eabd3d92a828b9fdae32096bdbf18a623c3796672c350742c8a889cbffcf68e118afec70e6e0470cae6c5d3a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3da2438b2a062e39134567358e1296071eaa0371e45de345321b85ba6fa55936c2960f4c24b5e1a59aa1a1829a5fd8b32f2995d3348f313ba5250d06fa95fd2b33bf832f1a525b94507003bb0dcc5acebb46c837a4c0daeb7f39638fa728423b98f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c5f5641e8cfbd0e79187bb42dc629a0b2e98f17f457cc307095d2f8d71ebf26ac99c518d62fdd7635cef670e68029aa6e691eac41db4dbb9699fda59963df2b59e1e1d9bb2cbb11d21de8eeb8b3b87e9077a70e47682194d74fa71fe51456b918e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e8cccb7a4d935128cc0e932d9117876483534b27e7f1d6f2b67f198f17299905fd2b0b86aea7a0697e84a8abaa5eced7b12923fb5642ba8d27c6593ce58c6ec6d784298b9fbf1b9ec0547adf35e644512583d0c3206951c224eace95a38715ee1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d036df739cf750ab26e60413724df6bf9267bad4393b22c2a0a9536a1d885992ac9b68dd7610415c3102fb30a07d85dfe2e83cc9866bce85bce432da02fb8f974f1d63fe0110e93da149b5f724682f9a92ae988280701ee0613d43a89c7f3a52247;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he071ac15a1946460f1ac52c5cda897cb2ab12ccb39d02af423a58cfd251178a6a95d1a0017074e5cbcc0dc01fe3b6f8152bd7c96236c1359b2f0c8f0416644b0e07b300f21ae71299f87b1d1c2d8ddd04ad4e193c8675aa069a6629bc5d51fa1e181;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha17fc797e33766c359f76abe7ac099e34d4a016e7ff2108e5e97f8dbeb57eaefd1cc127533174ac3b5c9cecef33d40df189606dc29bcd2d43383cf234bcf6c8104d20c57407bda9f8cc894375b73490d22205c9291bf693d361491dbe9783aceff0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14071980b4bee67e0f3a1ddaaaf3739d5a7136cff177496311119cc4fd436c21a9b32f0419dee371c8ba59c11d6ab32c4c0c6d65c032af25deef8bceef943d1b2d86661f8473e83290eb1914e5067537f74f6af721f7ca2909fb60117547d0694780;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdea96745615b09a29702e7c13f0988d670b86a49ff4725b8767af0d6102e40e1354e0a397b3a2ba4e1e063907aac735677b2e7a58f28ca4e226137f28b4226d11a0e72c289a79f9df1286f5346d3bfc8aed6c12aaa34299856a6db7f796e4bdda6c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72d8daf13397ebbb29618ed4f11d18571ae7b682264595b8af00b7fce1eefb98091784e77ea80211c328e01cf30245b3ff5db45a38a8da69e8694cafc244d0f73ff4b53ce6600a7e4117120f188baf94ca42379872d4950fe956d894bb9098baef25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b4ac27be0a4c1ac4b88af9a96d00f576b6b4ee08e6912e6e0906c999ef5e95ad9a90ac4eec594913d6afdbe18041dd0f315b35917dd805301af24b618ffee5cfe6775a86a7c9943e79e8e076b6704e6222ac79b75404cba053b6af678b77fd6ecd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d07273e0eef131c597154c9e0c639f386277467d73a1dcfc4f159bc05c26d943f3b41a3f1ba552b4d1e5238e71bfcc8f6ce5b8e1e148c33ef3946478df0e225c108fa99e2298cfb15f0161f6965adb408da5e770a830affd9d1616099193efab159;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h406c1e09ae065e3ee60200c122d84efe59b06fba22effc1de9c3a1479c29052f252ae64dd11f159bc182ad2f20d9526c02b3a9e51957f0ed8166d38793cac4dc78ad5c6c19f6e2b1264bbb96bb525e71a4d2025c26b0a884482de2345277c87a9998;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e7132a507a49d19758c0ecae9a4f11c1aefec17e37484df19c53460101e454e60e38701b048af73eccf40d8e8939dedb07acd724f224b8375fce67684007bb9444e742f16f94f6ff8855d3245c9db0de855a3fb793384a6ef56f24e539319fc5f70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f22a657972ef4bbb70920f4395ee0ef47b549e368e2e5fecd25bb399b0cab340174faa789a620b5654e5baab0f4253e0cc98d556a7f464a3316cbff2f3fdd07acf9bc70a4e5552c7e1d2a10e38128d3942488f087935c66367cd1ce03cf3dca93f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc6d16d0d756ae4fd58353b50c6639dfc5c7242f89fedea2a54691f1c6728882b2cf244565805a150b5b8ede1c6ac1183281357d4a3ff3276197ff278d8c423512dd30e2365b5d34a9cc7726a3e968ede0ff275ee4d88a02ec1f9822644492e74568;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90da831e0e1dda59d1d94da8010c61cdef19f12d39332cace0596c5c4c440703f66cd1f551e16673af15e598fe99fcaafeb8511efda383f798eb370f95082c6969e8e4878e49ae18bd4ace151336250000d54daf7d2a6fdd9047b737e6999065ccf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b75e8a5ce0253e731641710606ca86ed9367d47d8cdcaeb4c3d3956b828a545ed429dce98dcd5d5bb2a567ea400243b7f118a474739aa2e6d3e7bce4c0b013eec6bd12252f61f0265f114b60ee6e46977bd96ca31f383080d4e207c9ee4f8e159c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h355a3b91df50c773ba91b3784205f456455ccdeadb3de59430f42e321d728ec11e5fb30ad502fec03c8cb63c2da62f8cde45d591a0f9d0c07e6685a984f77c7e739395ab740b0471472e97c38a80dbfb873d6db227cf509f0b35238eca6d5b39b68d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h240f4cccde7db3cb2bf358a621a3cef00837031f1263e4a2b338b36d4f3106808b6c265827e3a8b957ab0759c9f8d0f94cefdf8e6b639bc56406dc635c7e8444dde845690fce8689501021ff5aa81b2e3131aaeb76596c05d36a7a1c15ae179f19b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1264e02d888926b45a9d1fd5018a0dd985301c3e875b48f4ec3494d47380a5aa38a31b856984b717dda019310d0119b36ac581406759f02905062ae188e96a08675bb5a538e0d23c8646ee77390e7e84201328ca8e519f3d3c66909b7ab2bdf0226c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6361af8c9958c509e6dcb06dcabe26858e8c8ce284d3d43e88937911de38db3e14fa177a91aa11ef8bfe2712fcc482289de13d162585c8863ccacda25ba5fc6ec7c4e691ee1df60cad47dfeae2b9b12fcf2d3186a713b3f196a3a972ab3d8c416f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52e16bb3be819df4eb0fc0b52869df525a556f122810da9914308f1a77a596290b8e0136352bc65f7e3631bb40429f147fdbc0a82c8efa7195b0028f825b6e78d1ab4036fa861a4e3e392d66c7e641165f45d30b362cb2d7e9671f09394a2afb35c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h435249cf78eddb22e07e1871fbda396640ee2d27eea048304694a8831f3f12226c82e74ff75bfa33166f78224691e4a0fd2f3e2f34b155bbd9cfd0e72ec261ed4a2f681ba173cd61cc2d780aa5b0253df2e1b128b8daa4e90fc7158b47ce4206f5e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1ff716bce0f0dc5890b5937eebc209e4a3020072abfbacac3ce7c2db885d091c05fa61e76a8dd11082de9438d58435b0fbe5a467935bf3b086fbab15767b6ebafb183d6361cdaf7d4e3051651f15b9a9f49080652652b042f8486a0aad8e5b92b90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70493a7701fd71c8bcb37ad94f5890aa80a82df09c81f52bdacda739b011183157b57c8648e738ad92522b533d58d31d2c4aafdb19f0653a2e7407d6c07c0cde35617cf88d53fa858d5e9090405df8b3836ef57297bb377b7102e44b2b47455332ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b4d9a9a7067c92aac81135bd3c427ea67c0418034888c08e31ba99bcf78be5915871cc0041f44171dc38eaf42824f2c3faeb9f0d99691be459aa458e0220412cf2077d2cac5fbe8f4aa57eaee6d709779d877290b40853ad4f9edbfc664accdb987;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a5458e854d5a8cb1a05ce5f8d7ce79aa24b0144aed89f1d0b21d05f0e35935f3c140a90eb59ec8425096ed810f61a40e02fb7bade5704320e62dc73ec548aff9a39fa725782e3b98117c48b17e41c33f5d51f93e76af785b571fcd63c813611c01b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde0532e5053611438f6cbe079b9995a98afaacac47f842d4242eaed53807f22cb1d607347c9abd20baf8f23bb5bc81c617bff4276d5c9f08653521229dc477baccfd7ab79834cf235d4ec21454adaae6860d1c25c7fc18ecfa7246376b73d5304cf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacedc65e24d15d78c4473cca63329a6fc49cf8a9d1328a1d5c60baec76a79b1f6efe34b9e3d86e37310ed808d6f136ad384d4942f3e3105a3c4120e1229cd5f43974f241e7de2aea7177a1490433b07cbc44ce5f9b3c0ddc37dd9d2f33577c74b79a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4b61d49f31a2f241c04c010830e0b34ddf5b96e4b2518c5da7c01ab43b23aeb67159d7754075e2a21f79ca6cc8ae6ee085ff3553f6fa56043c5b74b8b93afbad32fd099c7a2ae0d2cb44b98523534d5da4331da346a4dabb1e440aa74875a0cb847;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc08ae90f4274ff841995de0e8719cd1a672969c1fbaa39ae52a02a5b05b4c2a4ab43a1c9eb6ef7691efbb622f987545e66479e0362b1394f13652963ab4e208a3cf9b309e3323cbdaee6c5e19e3a54a5a79387eb64850dad13a89ad09509cb31d873;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9954f0c5aacb75438ecad3379435c402a1e27afdde019cf3f4adc29745129590a8f085ae102858352dd25d42d398747305747fe29cb6c58b01a975ea403c187ca76024b26dec5f08711cb29c1ddcfe3a6e1467e074743f0e6cf61994af912e9edf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69be35c8fd7b38519e608016de1ffe8872ebdd952eead469f4f4d1194d1156f79e54d8a3dedeb94b0fdacfb5ccb4b0c0ba89b9e2082dc4ef5fa7e5b7dffd44869873bf529e9c4730211a1551e0638b76d09d069189a885b3b19b8c0a5a762a8c4222;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0d998e6f14e89919dd67f7d5e84e29269a77d6ab21750369eba4486395cace7348451f36e1d2ebb64c44be68c5eabb57c2181a141028b4e989d9b17e398e5a35f210d50921407431281f0df3646a1fa9d1388770823940c2fe7e4fe33b6d393769a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fec2b5eb23d04598e751d1ca7310999a7dbe6701bcfb01f77683504ab168d86cee3dd74188300080a05f0a8cc296f9603c64618abf9aa0482f9a79fedc58fb964d2bedaa6184efa021acc277ce67c3aebb4b670a530f7db6839698a779cb395933f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8179097f4b0d8f7825f12ee7b4db524c3f6b094dfb77771c8d98a4d74ad0898866fa7ba889c388400f6cda1f845e87fcca5740e0bc98b674ed37425079467dbfcee621d1bba8e4a5d2d9d62f22a38820bf00f36f80953aed15ad4012084fec60eccc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f23ad6942d1bad07b46aba885e7225fd6535f8e9268f73cd9cf11686b43b0fdc3a2b02d29d3186a03b33e6919ea906c98fabe66ec8f49876a2e07e05e43809902437dcf09d33c6544bce33a809dddee22ea84e026db2ec1ebd987daa1a36caf8acf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62dab68bd8f49d7fb80ce536e6a8ff2a19b87e9558ec50bff945d86a4ca538c74c92d5f026cb2ede3bac3f5909d4eed2c9125fb2cca5c4c8f92f846ec9b93ba633b660ad9f5c9a29092394b5c09eb1e7dd2659b4ce4f21b7501bad5b2f56e858641d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb42081d62930893e55a0176561ee6f7051fd22d5393c4065064074bc6019f7306156d5f292d0f7d74c7875052974bdcae4cf807784e7b31fbef458bbf6771ebf15e84c2e1423f49795782c9e76af90d212a3b289b5f62bc081e0d3cf7135babcff98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5970d128abe633ae5ba41e0a5b8b05a2531450fd37429abb87dcaca0696ae2e0c23588b6f7721f9c7092e7500d8c108b3346a38f3336dc2828d2731ca9dbd2e03f37f2c4483b8e02b8a3132b2c3c3eb3c8e80dd14b59d759e900d0ac846fedee82b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1998b58c540b1348de90ef05a89811b8de760ba273ff96e63e7e73ff4bebeda1f2e6d230d56bd3b38cedcc5c2924dcc2ed11ad6ff090e2f633f67a5e26b58b5696df07bb5bc3612ec105731b3b190bf66b50c146e5c121942c22d4d67827fc45953;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1c29e016a0a44f29ae2f74f4a56d52deba6cd71fb915aca87c2e013f10e87c5912065ce6e8d0ec9ca4e0ae6d4aa35d3aa579b0074ce618c23d5a7309e89870b892690a1e3b1c5d23a14eae727d26e4c98cc9078143320c64d358522ba52131591c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea5d788d652fddc486ad9bdc9db162ce8b4308ae98f8c419f55b3952f329c09230eca59d16111f09883c126d72db2f86f795b71128c6ebdad7e3bc48f68263e8832fa13ab895127afa0c70d2133f32ed9550a8e14abe3657a2da4df21a205b5703cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53852d55cbb5224a33c66e7d0b8707a5acc22da6eb94629ce486502281ebdba71c6191a2a47d7f1624b4587971999d49049ec99d80779404d0e690e41989494cb0b1052cbe7b7a810c88f8ad17a71b02de29e6053ad29b7c78d7a46c117ab025df94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39b1b1ed132c55b68b4080cb9149b0fe7c4fb2c0d7c13804ee5a53d6642e80d9444cc2a4ec0453cda10d07c532b6df4917ae49f585464a0d5bf996914556977f38e972e5d3dfd5c084e71b4fd7adf7d71717566402713d8e352c065d818719beab16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb184400f50325aa94049bca500f9ad2e20614075778376ec8a226cc0010ecea4c35bc867112daa30a7b321bf4f8f091582033af6059a09cf2744f644853f06459c7c120354c7014bf3fa2ebfa9995db94fac7cfd3d4b38a3026142aef81e0ccbc12a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30d285b3a25e43de14248a9a01ef9b55cbff7386e1bb1fd75e344ef7696f036ae4028f32cf57ff1c38643306ee1278216e1ea6054919ccd037385ed1eec00f7d862e86e1adc2324b9d16514b4cd4651a155ee516b6451642c3c900d9ec4085bff444;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2dfd28bb982abb1b988b963a6334c6236fe9004043164c86cc39b5e7712b6fb37ba3fe7731e1cd645e0b5bceb72d542ae62e9f146891fc68742a37438cd803cc05aaff22bb4920c6f38d8e030cffbff81195534f4514a063b4294ee29ff52c56835;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbcfdfe91278425b75571f6ac54dbc8beb0c9e307435c1dc665bc2ab1792cc7425948da69c426f777a1dde8ffb5a1cc71ae0eabc68d3461318046f56ad645735ac58b71220ce04df5dbc7e7fa2f4bf2d78262f3f9dc8a3c381877f55fc13fee243a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h416e04704c0b4b14fef0dc91bd11aeb4d1b133fbfa2c35132cfd21df2bd946e988e2738e65233bef202cc49c89526dea40ee0afd7885aa97c2127d3c2103595944b52fbfc66920e5140169a95dd375a8f75c8179eee91151b5ca30366382fb60c24a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec51ec01d5f0af2d6150e52bbc9fc2f1a15d8351befcafc13d99e3fc44ed287d5628a45e936b893f5f078b1dbf0691ff82611ae370e207e07735ef3148e1f0a6ac06a42edd1be15601ecff71e18ec096658dfbec2195d13fe2d64e4dadd1944fad56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59dae1fae4ac74d56eb12e3842386ae366d59a9d874bcdeed2a3e3a7ea4a0f8d58749227207aab4bb522c914d076003b47c687c681ce84ef2d8ab15c47034e87611db862133c3e6e2b557a3bf6077fad553af0379c068dead71575702c25be98dd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fe848bce793339e24a3f741e56149539e9dedf5c7a62abf380341f86ca0611b2a1e52f7c20c2a8765da58c3ac2e01b180f588d4c9f106166372152cc346647b9597dcb07cea331d55d33840b69ed7f28a532cd781a0ba8cb258a0b6ace366ff70f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf03e799377b085c3bed6c64801397e6602a68d5e68de5d085f0779fbef8ad3bec17763461304ef58b036b0fdaff8b2e2d716b803f994488437448af4f951f3325b907fb958fc5e9f1f3be12790bdc976f39c0649663222d7f1d2b77e4a42c996373;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb57d99ff5b1c26891379d5226cad767601cf18f7f14f542144a19429255556d876573088e49abe2aa520b6f595a439cda3fcf3cf62d2c3fafb6feea945745f18fcee331b1fc37ca4ede7d5b8eb4153e2de50dd5b476df9b39fad71bc1ea0e8f873a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5100a5cd78dc406ced1c540b036c5e749d2a219f2008885861fa5f641aa8c1d8f7d978404a0210621d20d887f421b15b856543c7d90edd7dac92b464e7c3a8b5db520b700fc55604b4ddff2cab1ad49603779432c7dde065024dd990dd5d352a1d7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3dcabd6756699a1a30a7574052ddce3184e1f5ceef662a318a75a78e12860b62c1807f8053b20d495579966434d54cb9999fb253bff274ee8d0e057ffd67fe744e772f5066b095939bc24d6c13d2f1c8e16caa2a3b0b3e52f31a72877eda9bb8485;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h636d3fffa3c6752b06cc55805a060319b82042ecb70f2af7f2fb951db8fe75ddee6385b4e79f12252ff81f2ca819ba4fd6b23c3e9e5bbfd458f88b1fa1e1a94c509df590035373cbbfd8e7ff026aa5ce441c60e0a48e99280a1e70ae87126d8eab8b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he40f61bac96f119c914e5a5bfa770cb92f17b9ec9235a5d2871b3d8288afe096853156000d1cb72dd9c512c02bc6823bbc1ae8f96e0f89ad441de926b6ec8fc2a770ab83accafa5a9685163f0cf11b94274c96ba0119cada002f5a4151aabcba8bb6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef54c4328e3809fd2fa7c5ba53bc13093aeca1a3ce2752440233f08c073439eac50cd72e8f5a80dfbf846632b3ae5ca1b1b783a8a8e551460720c08fb5aab73afd53f88ffb595cf3fb59ea7442157d9a5cbcb6d35d314e689bcad32edf5e4ce78ccc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30a55f28783f3e941fe65973136f79237808f5de8cea9d6caf2d98a4ab0d66426465782c798e63406b129cee4e4fc5e93a0bf4e76c927dd52ef51e5820ad6a170c8bd30868bcbee0a9d39c8fc454aa2e25cf03e6710a595fad77658dbd4da7461dd4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1626ca6aab7429a2debec7e8c6064f4e0cc124c3a6f8615af76ee751d55468f7c273e0347d309d40f19ce7fb0f37cbda69d212bb35c879bf05476df8f556cd9438c5bdb40974430a93112f32a66ebe81d94901461bc3ba91a04526769261a0d8b10b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e1593564cf22ee7273c4bc4e0cdb066d94f50f22af944cbc6188c1e91c87f16002a570b41f89913663a64060467e5e7c3f4626b7308422e795bad585fe6a520daca5d43a12a75fc8fefbb628b634918cf034c8bc89b2872f983f6ba7f30438edee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c00adb5cc419d9a6ff2b0574fd6e9b3d78c2ab18960f77bdc33c84142f3e69bd5d176062ba73b5590b528aef1992e04eed2040c914e5434952562e996e078d6ca22fe3eb56e440dedcf19f98a63f248acb486b3ca83266684b6df0fc199c58560c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee5b4ae297599ad0a364fdb72867cb0630d12bef0c1e439aff3695a4e5e63fe689337c5d9fd3b368e6b73fe40bc9fa613ad3cd8b53e34ced8270eba9f8bbe55067f5a78cc7f3e18a95b3b865fd0e7dd0563020543a30491b58dc7b698f308481de32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ef3f061235e5dd263d998ec2418982f4e19a1a7f569956c46bd87220be89fc3f3867c3c4a4b2dc8fc5adfe311eb5dcf583a1f27eff1dcefafd30ec38e8e6cbf70ef6821d2f3351f634557572beeb89173d54daec5d2fc2507ccec9c33cc40a3d47a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17c47b0282bc4ba86a56afb9e478b23aa7eb48fc790f8431af8f70bbe16ec8c7e6a81f40f407a0d6b2c9dbba7c0975ff3a6a9f7d15bdef17c946fc9bc330197e0cfd3e97d3b6c4fed6e79849c90a1d5aebdac895335d692a52e043f45f8d3dfcc7c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h788dfe151966fa45362ca155aceb98d5dd78d6a9aeb0ad12fab00f26f8bbf7b152b556a6553eb2100d497585332f677e4d74d9eb1ca5c7591348820a6a5fb7c8aa83bd4a8158d709d0f52a9ae62ee2272795dbc5643e5a26b85630b28a74ee75cf74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f7ea9cbcda08c1b3c992cf54beb95bb476bd9ecd98c2921b4b44b244b09e03a35d88613f0d6b373799aceee081dd0d24a6dd5917efaf860550979e26d05c63b9250fe4def800f3db9521862d3c180efb53aa1188275bea6b24b414f7ad3358a888c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ceaa8cc20b3efc0a66d42e2906ca55838a804de304f7b794d48726c15737aa2c97ac451a0879d151db9c8e57e9cb596f66868c6a0a99d8b9ddda08e46ea31ef22e7912179e124f1bf80d71363856b920035e45124f64a5e5a952a3bd3722704b246;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h369c0f2e3c4e1fb8e814dc5e4f1fb384ee86cd066efa2b3ac4feca50b333aff65195a66c03da10349fe1cd3f5971e0d8a7608440f0032ed396113b6d80d1d495f3756d727eab3473094dcb160e362ba6dfed3b430777f8106eaef4182b89783881e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc9432ad63be0bd2e6131aa618240f19ad90b0de33d7f160af3e17eb723a49cede86a554da459173dd4cbcf30fed47bc9f993c0232bbaecade62154aebb6708e4343239056e5431565cc6d54b201aeaedce6178c291a312c0d89876f3f91df37239b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4539f4a0564f18a9a3f537bcfdfc0fa2482d6b9af1ac6c0fbe614bb59be3b80f7b40e4f40128262fbf33aea1c71c6b512e7bdbb3def2d96f7fbf659d7876ef46cea7d9febc9f7c03e813145f3a7a8667bf7ae36bda86c4f7d37cf01ff237bfdb1d81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20c36094a0968798f97e886be7f817aaf6a53e7ac8fbd43a1020209104da1948518e58541422e7d2830e2b33e116f7e8f6a0242e43fd7cb9e7cb868d40f00555e6479223ccbd1c794245fd0564651e009bf018a443bb4454df08eab8521f731609aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6e956e264c202b38d157a0800ef701fa3d2d96894c8287d383e0e32acc50a95d5facdf2280cdeda85781dc7375970874f66db4e7b7398fd09baa49b69259112c83e377dd38d10c8c74dd1c61b48f0c4386ff36b3dac2ab72b14738c582c33352d63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d73ce8dfc4d76f77285af8cfa890224cc71cdc04f0e1b87b8051b86f92adf6d8220a1be14d07b089d9f5ba7966a6813d69b4595dee1cd603d48188381992035a34d81a62cdadbf84686d2cc51d13ba2123e23a31cd6b9e4f80ee1e2bc06aaa2748d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3168692ad3be85d9395bf32cd8405bf22f796354a73c3ffe9b70c91e1a284ede36c19d9b693e446c5fd936f874ae913ee80178de25333e8e61b596e46f025a9f5fbff6e7c751864599a740ff252bc180459772d5276b93b324333fdd985756d1eea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22e889ca89d0608beb5f52916957db5012b037d535630e13daa88a8a453ad369f2dfa5fcb75dd742357152e44cdc3939219b3e147f8f9ba412dbe28b7cb83043015f9417ad8ce786ea5ac1a6fd82635119af4cec4d8de6ccb806db265d6d6aff8bc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19800e0b6d1d620fb14a0479fb177674b227e91547c52fcb82fbebde7fd052cd8526a8dfd15da273df4680f716db6803b127063a6fcde75f645de3cf60b8a3a3a1118de168d84970f612a806f4f6eb17eb5e45f8268cc41bed2c9739db94051313e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef81159a4717cbe04597d17d7575e82226df505971377228813ea5358ec0b722b0d1450583348491854bcc8adc640f6d2a834d230b1330eba1a80e932d54374b11cec63728343884aa4cf6c816b5271c5fb1309910690094faa2f18fc13f5f3457f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c785495d870cf886ec974b48caba461e6d30e9290363a1842077aa6ff97b555aa9f6a42adcf088e49554260026b3b0f01866c628c7ac47d1e2e7a518c6d03ea554cdff3ca0e3028946f1e08e85d654c5002727f5ed0dba20b77f96e44d0792b853b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0ad267a02928ce5949da23f2b6805a951b19c6c0599b7f8e59d4ab0a6704dd2e527217e6e1be52ed0f119f78fee07bc14663661ea3d72b8e8c991d6f552b50eddd564a3054af95095118efae926e49b046ab2b52615ad41d19d28a5630259fa40ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b4166e58e9a6903a1b2404d66586e22a391d55b5c3d9fb36f5239d8032a5fa40053b9e458b4d11845889f5a95b55d1dd2e18240ff71d2120772b0c1dedc1f051110f6309ad3895af3b84ac927f3b587c03498f7d2bf1644662978e0612f653fbe5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86fa3e8c7e998dd5f770cd113ea820c9f1b74b769fa20737a4aa8ceb5fb51a631aa7ae057eb6cbea34e7e0899b8aa52c14c90898e972269765f5a6463c5b56b7005b9049cc32e228432ac75972f87ed4a64b55c98720f7bfb1a4f923e9a09df734a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99a098b6d3fb131121aa174d7d3b25d746dd3b9e0a0be3dcbfc0d6b67d371c2db8b92734993af2411381531df144f09c4414c1b687cfc82d3969b4f5aadd3f29803f7ef5a344e7f9170fa664b77feff54ae142968d2e1ffb7fcf52723197936840e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha91e030450783be0ec05593a6dc4c56f2c6d8a07f4cfb06375a98740fa0d45a32ac1501e8471909ae921a8fefacc57ebe792a5bf7bad90ce66665aa1d3df76be9353be9966f43b2965b5536947d88abd3a2d0cf092cbb5d74a79bb46267cbb66b47b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbbf13f302fb6ce631bddcc2cbf3f3beb31819c34d237022132fbeeac6273ba6b98599bf188a7636309ffcabc13b283935ef8f327591c574e44958481b6a82065eb60e884fd85eeec0a8fca7c57736bcaf9ecd11a6db2a029054d908a985c40cce81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf314b90641cbc3d21c6f45ff7668147c78160dbfa3f99a075f73c480440ea46c1266bba3ead9213f45dea791a5e2df8a56b13540f13e6ddb2ee59549a3f4d7eabec80d166d870b33c89f13298e97a744f91a56504d160190a1eeccee35ca15dfa39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f0743bdbb2f957af98eef4134cc59131f16388d30da24a006f17cf30e709f1960eef5360eddc37571ff4277dac153877bbc8db9847c4c62a78a8e257712d392c7616c61ff198112b0f741166ddcc2fb42bb47b1c2ff39a2f7a1937fc327cbcb32ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7235a1282358e1aff1491d98648ea3e0c141ccbed00b5b94ccb0e62905cf0f4a0fb95f424826ed354406b67fd90761f063568a6969ed12873e08afda23485a5772399903467d6bc33d3060f34622136fc5148b1318fd1b20ed19f7ead5d6ca00f104;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8a6d61817eee9af47e9c568a2f2c31859c5ded2591292f55194645998cae0c8c00cfb3f6e59c9ec791fc34e5791103d9db1f06fd89a8394b084a58ea65e89f1623b951d65f96adfd6fddda6b42b20deec21dbd213a9cdca57780957a9329dbd4422;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7458d5365639627c35bd18f55184ba413973b187437a1c1d7d7fad598ed9a5a6e1531dc650e0136c28460d00dd6e9f4eca3c0c100256f89f6bfd7c4663c7c0109bfff6e6ddfd2a0a153fa87210e1650d50712aff192ee1ca41e539ad76504bb0d8ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbdecda0475ce0e0455658d03b6dacb810f125f8a3c73f3f8ffbc6601e7dfc031a15de8dd56a3a3581d736de8396bb97dc35a7e83c02c893e36e149cc6ecc4ba2f83d35b57f7afbf082b75e6391077a88f4c1cdf82445dc4cdc8a14dab03df831c1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ebe91e970be02974eafac72d949e4d132645ae128714c2c4650d76e70788fde6a1b0004f1c60966347454fb1cb782da1528acf027f8cb0faee7c400be8e09b7962008f995262abd015eca2dc29968ce906b936a662e782c3f7ff284ad45226f683;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bda165af8dd30c28a29f37cb31f0437bf831b160dc5754ff2b1eabbfbc3bc99cd2189eff066e14574061a0d6b008e52482a95892a0accf3e0902f33aeba580fc1039f28abaf48c54f43df62e3e27acb3e1e8ddd4bfda408e13ab0908c786667ba76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89c588b3f03c80f01e93a268038f9f25bfeb1450040d1c2bc583db66b3ff213654dc9cec4125dedf6651dd415d14ad292f5dc4f3cae8e8e79e39734cc403a0f768fdb60cd8e51e454d50613937a2bfcc7a1d49425b7640d3e50b1f9c603273331ec6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5b63dc6ff7d1f59e091c265c45ebcc1c0ce06473707e1980b5d385e898eab116518ad20f1e5fba9cfb82b054a7d8110a345891048c9a37af16d2247f249041b1c6711db8699230ba074f8692962acd44c86ed8527bfee6f7858cae448864a8197f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92c9906b9943d79c7e59d8b94844b9b725bc8daab6a62a01bd2db2b07ae4fb89eef2f860d33794f16bc1a552d398b8aa198c46829c2eb093bfa12d160fa9ede638a7f524707bb1b180a19b7cb1fff79650f45a2a08a3016946736f6b6cbe29c7ff23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6d7fdfbf23e2d024e64fa445f71e8121f90f1c49ede57416f4a88e5aacb979df6d8ee73ca826fe1932a1260cdf5e94c1b22d0fa47abfbfd1300ea41fd6d5fb98488be53e9ff87f76a4ad3789a159b46edc3bea37cbda1dcb05cb640c98d518d9b31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf45056ac24c88b379de80f7745ee476ef9ebaebd36118b1559541dca90df2af8fc8379534ae1125353f504ab6fe1151f9f43d149f3ec63221c022a314b99664f16a64e1bdebf58db6adbd94fa8a241deaf76f6b4a5fe8e11f1e11364109b36612384;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde5f7e526d3c5a3be3f15b07c724339a6154771e2c019111eb2a9a84900a1789f62a4f50eb89333b40477f9ea833909b660033a3231fb12de22cfe88bfb919d587799948d84397c60a20bf2be253556e0e36905737e8b845a354cff2772ea27f2331;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35e0459e8aea516ad4e60751daeff6e23406f97dea44fee079b4670d91e2584469acf5fc57f65f61a0968c248d6650469690759277b580ff70261190171ae8867898905bb00ae5c0236d353e8655700962057a62daf7964b0f5fcc8b4a5952e48720;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha11ffcf964aaa4f9a31d9482122fee566d33cb030a29060e1ee1a5d8c0794b33326206b0caee81d015642669d76fdbd9223348edcd9fb44f3c3455af937e48a14426095ecfcbe85a45dcbdafdeb6c9f27b1cbe506516473a4c8df22b6494a8eb48bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38dd0ce78afc67c217adac5b190dc3dedd82f5521dfe4b89ec0e8c890845605918cce7b2737404d17cb1e045aab3c0ba1222f93b37fc3e6547e2c3ef592b373c20c9c18bbbe8332a9af544b7dfab2b545a953e3133808c6eb1751df54c4541fd2048;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0e3b4e1be8089ceff933d79b70024b9fd9e986d73381728f6970aa4006904b2d0a8bbcc4cd76f836a70e8f155035f572e4784b59016380bc3d9e4a36318723e1eabda2106f4828ea72048ac58381c5491e9a0ce93b49f9591bbe658336580335bf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb05a99e1f4cb2871da603d87b69d8e1fa3403c3c91465fe4dfa31a28c911f41a09fbb933b1eedfa98658922697fdfbdf63ce717a078130d12d6fa3516b4619b48dfda3e0bbd20b7990295f0208976740a0c4a40da6b214a2fba3537c4a306b5c42f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21e4b1efb689749c4b515779c8f1e6d5a1f866a1b05dc2821b5c3be9afe93a136b1e571d0e46a855d90b71772e0e081a2ead6d78be4851c7f797096bb10fd3a58bcd844680d5bcb0c0c8481e8efe68d6c65d4bb87ab435e13c233553f229edf8ae1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e0bc6bd060e34fed193e7278faf3015ded3f2032e5fdff1204e77b7b6b2047bf6b72f88729a256e6a7f90b3c5c516583f84d8174b9c189595cefb87378220201ee1a553ce486f654c11fdc2cd6c0098be6404d635de7a19d60996b40ed54e84f127;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4871e1617ed2e75a9b77f7c6320212257cdc81317ee6159fb8af1a4294ce1de2ff72a67ab9d9b5da1b30a1bb16ee3ca4586a60ed2437ee7975b17396a78577e3da1799b9e696c793abdbff7dac8d5dcb7f9a9a4854f87ff1c8e7f9291c7d12fb21f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a0d06da2c5278c364a3af407dfc1d8ccdc4994ce6dbbed88938d1fb01854274141d63b82f37ab533cc8fe582c85d0e3b025cf2ea0c62c108ffae76e68c3182581e314f6fa2289f8d2e5fca130dfb9242102bc153b76d6a9bfa40fefa52c16d706ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2423b7129f763765f31a40ad284045498b565bad0a0fd91c1793024d658b42b0ab7d62eeb96fa081904bf69ea26fe1f315e5e0c5d1b726dbc8b9dd2a60364da0fdf73cb5d4f36e3f678fc967c5b065a61c10b27fa25f121b5295084672cc752c509;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h466b452028932719d4e436f2c692429b76591be1da0b5de1567d8f493a4354bf8bc71582540e15cd3c97ed21237d6e743976f4ac3076795bf1f4295f19480ff4fb03df53d1bbb742bff60e54feee62e8b9db58b4c3e4f6229846db5c41249d7c8484;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc44bccbddf1a98de4ce19326002529ed4869a71e0cbd2e2ebd1cc6a7409f24774b026de78e14750f23d11ba37c93878be6841186887a8dc5014a375f6d46f3fbaa9888c7aae5bba7a918e63fd247f65aaf5e35982a7ee732af393b03a1e03b650a3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e378ca55100424bc0669b3497cf1190f28209364b653ae6811387b53df5dd1f47b3300b8abc0ace90795580ee34b6158c7b14e200974fbc634e6f460a30d137b9983853b79ccd23f84c5da13b89b928a7c0de0c90bfed30afd812370c6d5fc606b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dab4d8515a3ff3bc42d5b369c4b4dbdf7a4ba7e64997172fa7ed4ea799a80bf2e42e790620a7fdaea7abe46ae54eecaafb8670c4c6ed704781f288b8457715fd574f4317de509b39a8fc89e66877c4cbf423f787a86b461fa490a4efdaf3fb689d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h967e76f9804393f33c59ea3974e414c2fd34fa4c608d791879d08eead0723a14d880fcc40e308bb8bd66b3d0901075479d8cc4fc759c38db973bc5912270d7200dbefb3660795454185d080dded64ceb7d8963a85efdac7e114587b3a4339a8134eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h397d056f427dadf6f103ebd54f45d7f825a21384bec32b7576458599f5e0b87014c1a9abeea648b2c06f9fadc6b589b97560195625a1ec9ea5864f1f6287df0e20f4652b063e0203305829b694c26c7f36272fce7e1cb015c5d3931ca90200d74384;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h987ef33ffcdfb73a02ea44e2d518a508e292755c258eeba5c988594f9de3eafa6edc76c36a394a2d57c0418f60477e6025aa38e23c591aff979e63855759316827242170b0e4bf545fb219022d6671993604c337ea56bb3843d8ebfa8bfb42a6e887;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7623248778e129d039190b4ef91aef9ab0f431b5ec387cb29444d9d1ab3687743e314c755a608173635f583788f058067efb4ebdffffcf4174d7455abf87cbf5fd3a7c3e08447a1fd11b5b7ce3f4e899a6e21234b54fea4c08b1d51a875efccb8cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f5ce34e3a20bd6da70516c2e1d4a1b3f667143fd47b69588035575f13351dc0e5ae8592867c07c91557faa4e5a654b2ce52ca58297be5bb0915f86f560a0a19e852d51787b02c9f972889018a86cdeb0ac5d7001558587eb20be1c0c32d347a25cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43ca9a595fa995e7cec0b3402d426675d12fa07521a3a337c93f54dfdfef4560cc5ed1c23926a7f957af130d126ce20753e82248d9cedb24f6a8b5fc50ca5d8f20c4268f9816843409245d574dd327719d0ad2f35374b577e694fa8fd6182eb7f42b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd792a3faac58ac2d58c8bc43495d1d26b184b262b0fb36ed41700b52a0e3b7e5c672e7de71f734652f8bf9bdc8603c71a9231fb5f3454822110bcfc2337ee4de1faf2a26afe1e3be35a0d34f2eabc59dd31ef6732bf81e6e75855158731f1e8fe9e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa0cfc28235d2c9331c6e03ba2f03abdceb624ff7576faa7f79045f16b2fd37b1267f030c186dbf3f60e743c327feab49f923ce8b58dff373e8bf8fec22521b4fd23905f0d241d530e29c2664fa11b2d692857d811f9905dcead9660880ffb62f29a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h173ef1540c1a8c25db4f948c9e3f2a1775bdce4ae31bb3e7f1f1f631cdd07178f7f12fd4f237be63692ff32e77492e4c45586ae2ea406ee5beef480d35bdf6b41654baf4d5628b2e67d77a70cd325e069a4895bfdc0a4276b18ed0302bb35137c309;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4605631ff92b200ed07f4c0fac9c16beb3f09a908dfd917457a06cfbde125753417e3f33c17e2f1e346c15f6abfa90935f20974d2bb41610d95bac3e948967c3955777edb4d9ad7aca7f14c9fc30a590bf08f59352fae9ed619663f6791d2097d9fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94fe5b37a7f778f172a245a86293e6946540a4a5502773b99b595623764e9d7f0ce25f3bb0d7a942af3701f98141f83a7765421fa45e6f52902e437e42dcf8e4225b0928d6529d669171b5ba4f4e082f55baf94d94299faecd5efe8573693f5cb727;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea88f9cc326875718e19b78cd872e7de0ef5c2153f0bb3ec153de6395cf642847fb2f8ad4cd00e2599db9fab5a1a7b25f5f8f396e0a2a10ed9d67ae7d28fbadcda87229d043cd5fe7e50b084043188076f1bfc856578f92f7b2ab1716393a716a60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h291fdcb4c17f7d31a12b65da0397587faf5ef8b920be37fdc9e32bd4d3fc172d6be1f174c83423701395674bf712b95334d4b4c315c179a674eb41e05add99be7c7d5d9c92253dff398466f8a585b3d9c7b44b18684890708c36e9fed4f411ee1f35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h792064a86eba236d93599677f546156f79c5385e4ca6399e53f84b99a694f1dc086f5cf387ca301c448f03bb3a91ad317396613364e6096b514aed4ab5a61de093101711ef1d173c74ed425d3923086719e50e778cc9bf8141cda845fd57924eabef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1426d9477dd64561aa002f7ec363a42908fb9e2b39c932be82e3644d069f0c6a7cb3a8c7c5a23247f7edf0727738687f97a5eab5c296c817d653424c7e59c733915ffcd073b955b61eb9bea9196f8f4be480278c72e6e1dd3875b69deb85fedf2d96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec79de86f49728c9078c2aecfec5e5e0934123ef69bedf511850d0415ea2a193c146d050201e33988ffc6f5e6cdb0e8843566df9ceb859c9cf1c96606dc6102cc75855bb5142cd19818c2dc825f14fffd9d4d1289e3bc08a89a2864aaf8446533b1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b7d66357a2e0c3496c296a10b00f26f5a9d4794f8b9626cdfe521440bc177688316cd5e68580d432fd593684108d936546ffe24418f5e21b2293a4d60d3c0fff0d3c6d6aba1f541d9464a5e7d1f60891c3cf8f48de457101102af098320404e0db0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3104cb5e6c3d916d646ef88ab463fe4fb3a3fcde353ef3e7c7242f512e98e555d165a1eca9f5349411100c5e6831723919c5a37baa6db7d95ce81816b86a5aa2163e08736ea9486cc98d377946b06c359ae739963cc0dc5c6974e3edb93eddd28082;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf18c7ba67b152f114884f59c605d93161757dded5baa59a8f41a5a2e5cba41e796373040cfbdea08b627a1a96c8a4980df3cb56001b6e3583d2264cb1313e0e892c2a0a3ddf4d8cd56204b81f29bc1925d5c0c8c1e07ce9958e9ed63ff0d37a175c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fa73377dde7511355603054123ccbfc39a05456d010ae21e3a4847c70c2aded4857266ad2cf96aaa9fbd7415ac598029219452191a270534772145e8f180b8dfce89e15fdd402ac29e42038767ea598fd8058aa3c4e89641ded354501af2b45e9cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd794972214a599c39f7554ad3acd586db42f58b06eaa8f6563d352dbdde45cf532cf979aa9c1673e45c6077395a83c52ec29b0d3869096353aed8d98c93a91f50068a4169c1bd23047f70dc69fefa258723195ff248ff9d6bb1b3667889d83805f2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc0500fa7cd662d0dbaf087e3fe52c7680eeb716083152ae462f7f262a2f37803f0d02050952f4c9ff13f3ae22f40b3359fe50580acbdd69ddc23cd920a0b4d9311a830c30033bdd0b4f52bc22cf3a9faff7e15c0a4059ba6ed6131b54433e72a88e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53710fa1be964e339550ee39ccb8602d4cbf2f1794009092e51f1032679cf9ec086553282775e48dee1a50f2b1c669f86d22e62dc74131c89305a08c61639a5b1e1a7ea77fd3767154e83258c23257d15e702c072f6744bcc36961b1b5d4b5ddb8ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h857aa0eb1c530cce7b9b51df94a9b6bde837e4f71e82783755c2259832e507bede4e90564ba0e97ecc9e8830a390b26c2c10bd84bed1ef07df6b6e3df7cf45b9359124b83b6794cc0f7d1f5b1fc0904a27a44c445107cfff0e5f4b49d8dda73697cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd25b7981cc24da607baa9a92de68c12894bc5dc638fc4401753523d6e31625910bda94c674fb28901fe68dd66d1e0d003dc7974a82ac6037ee8017283e3a7d25936e2bfee34521a273e19f2454e12215e5972f2ef68e520a8b37374292e7b089df9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5eb5af0c569b25e55c5f7a1bd3204648946f8ea9fb45ca81d2382399c4255a5e0c174b022df5171462f9851945bf5bedf477153126be6689b6414e7c9491dd9fec298295c0d0dead30ff99699fac92848e7ffa527c0e46a6ff6e78682d2f33edf0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cbd1904b835f9cedd18e5cc841a85f748997495cd656eea438c1ae73a87aaea34a52f1fd21c534d58742278cfc067411e50e6ed4eb2cdb6f6b1ebb8d13b31418f6483291f97e20db82d31351e66c0a820509fcd32a8ec6da7877ff48b5473aa9893;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1787313c863980f3cf209f8173adfe18ecbb9426424d6234d10622cd365a12a413531526f177185a07882892b936eec8088258ee0dc84a5814806dcf7182acf7b0635fd6ce87a96d25c5b0606c2f4729f4bd037b52620ceb8195f960335c539d3f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb3b9b65a6a1e99a09ba30ad2c49d9acecd073c3c225daa4886ed6da7664825c1ebd0ce5d8badc94a188848fa17b9ec76a1f54811ddc519fe04d9d03badf76033f855080ded65f03c63d363842ef36739bce9c80b38fc7e6bc21760d42ac4252c48e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a27cc3d7bec60b7595105f886ebc02a799ac9bf4aee4e5aea7b5005176353f4a1c9b11a68100ba117b0c85f4fd9c1008181447843e5f8c40474f6288167694f5385a86a548be655f314f263effdc47d0726cb0602b9d55e6e48c99dabdf9fe14b48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb77b928f774e30667d1dcb2953b10a7b41a6016e0c2c86827387e8420e0f71d4cd72cd8d8e513916472548d1331d6834732129086b637b698a047a2392846047777419e0dddd835a0d329caa2dd2735da30bd764d6467154646202e0bc44a4b8aea2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf620a309d3baa048b54a470994a085de87c266e8085aa0ddb7f36231e85e8ba8ec76663ce08ae711bc6d31a46640c3024e07f1f005831753b9a3b831a2c99be5e4dd23873a2d1de28a0a86ff078d186e25474fe7dae31f7c42721fd402f4041687de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ebbe5733800b2d5592290840317ef38966ca3dbbfc293be8b6b58071605109ff0fdcb0d3090ce4b03302f7c7c2a339e477b98af20df581d317ebf9f64a1850b7f3ed8ffc359e7348275995b33af976b016e760ed814e4e10fb2a4bf219310625cc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48374a2b92982ed76c0afd98b7ae5d98e2a495db9bf808aba14d66308ac2fde12bcfdabf2b7150787735d729fd32d8f8b5056c2891b6c614671c981b5f41b0b8c891d6fe434bf1496e870db9395f48287f226c71f3fb77ec9279e27684fe240decff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89a0b1e56d5dca831a85d42a71683134432aa7d5dd7308b49407f6254422e67cc20afb16b7c59c4a6d520527f46a4b077cb0bb68fc7cd26bf078f2dc0cff809a8e212b503dacfe8e15c493cbeafaa2cc31a23c3e4994e09243ebaa66b81d621c0847;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9426711145ca84eaac4affd0b24eb641219160bdfd85e11ae41dae673d41ac41ec4d2270923e5d38b3d18afc33e23adb6c1a16dbab45b31688a1064f14fc96e4220403991b6d0f16133d3427d31d00feec696d6b6551fd79971430cac34279b05a7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4d0f7748c50661e6906681caff22c777ead2badf48029aa9cc83b7b4da95f87f034b93b3f1592380b775d5e473342ee1b069d7462dee4414061487af6f9e8c3545677b23d05b74639571987f79bccb27b525f3c78409dad8dadbef62231aa1ab715;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa21e0ee3693f838a47b7dc858e422c6b452a9506c9d44048d8ef1ab8e84a42b75b76d86f1c95f26a2c8a50944a26fa6f50bf5949fdd3293756711dbf95f86e64bf956349256236f438824686cbd4953ae436d6c8541e442ae40679f3f677dcf6d8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h878993d439f6e84d5273a4361c4df0ec52a2383dfbe4d15a9309ef0432c465340881be45d02c6c4ca2562c3b776083adb9fbb20d9742e4c2b2800fbe0718a4e09d1c42e8362aa2da83bddbdd0f4d79c42c5c78d59f023eb23b2920f0f66494dbfdd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h121d617856da36e038245f38b0e65713a13d833337230ea8703a996914a28f1ceb36481f7682989e9a1a4f9f326dde5e0dd55f34f052ca58172d8a75dc785e99b43ef1b0c6a6b3688e4d86c30fc5b071e5f0af8a7958d19dacc8b4dbedb7dc857cd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a8898d5aa0245fc38a3db9f5fffb1a5b3be0438b1c49540da3edc49de69649217460beac101ffd3cbcf5fba3f091d9cd1854aac152afb53b37228c4f11cc58fe742f3d338ed9aa83707fcb7ba4c466d87c35cab6e3ac70ab8ec95d9fcd4a33439d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc45312abd03b22443e19eff5e533cccb0fb36e5ba5a9288cd847fc52cb47ad8683efd6780a38527f19ef5c69eb4963247a44eb4741c20fde31f9d9639c915e4bb10ba4b818f234e8fa874574a0b783e102910f11c1fb070e354367427dd5f3a913dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8fa6382e4b268524651d40890586a32c27277c921f7ca320b213cb0ddbe38912369b95c5fc00df4a4e049fdf1a68767a256b7893913bb71b08c91b34fe19892504e03c0c2891f1e9b033078b246ae0013a5b75bf6de11031257f51af06f90307682;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd333d27faa1c431438521cacc0b4b2d650be6f779a3b3fcc2c4ea7e1329e2ad02da1f30853916a950e3f1ff2bfe3556fd295405d40f2bfa4d06126f14167489f2adb290371558320b57dd6f15bf12b59c4d6ae59413673f36ff945de65de46a6f87b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h182447f7e1788adcf95e408be26b8ec5985c0c48326073c43e86211432146f53c6771ccda8b8f8c0c08e6a3c42f68d68ca10f97bf482eb2243202d7558c15f966c71feb838694a04ec05db45763adbf4725409d276aa43942b74ff85f911c72e953f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2935dea8c9be5bd30c5b1dd2f83b4aeb10d7a546a3136f81ea96ae96a03d3190dc5471245bdc47a3bd01991a25bbd329c66b14fcbc59623b93694c5f757c613807073b86c4b239878d654e1d6cf41dae10f3f5af8f211988ba490324e66068e841;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf22521618c21c453b62999f098a4760ce5a5dd559d1da740bf0f09af6e1e213b33fc35e37029d7304ce5bd0a34f126038b5f817f3965a22bcedd8dc5799e006dcd135eff873fa3646dc77e08abc78f8226bcbcd448c5b2a9bcc6439e206065d52e87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h332235473c67134ae5c1202933cb7ab3375280c60c7a955ce81c3cadd00e482d648b83aaa37d4aa4773a1fcbf3649d5c696e1ea6490cd510b04310ade4f4f9f7edd8a4428353c45b55de871e9eb078dac85809f76c30ed0438781c3c7d5e9c78a8ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6eb76a672bbce9ef1a8ac0537d3d457b0ae3a2ea3466074ff01ef1b494cbd6079783ac8a4f461d39662a49836ba13a096fffb95882f6ca4742f3685ed64a28998a22dc8ae795dceb57898228421e2fa9532c114621ccc2bf358ba7dbef2fa1fe296d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc3b8aea12b55a9d808e5cf79e6ae244cddad82fc34be898e307677ecef517990b8490020bfdd7ee449ed6558eb867d6dbb7dee2bc6e8d784bb0db7219c372158eeebd9e68c5b7f49bcae6a3bdf7e2f7bc619dd1bf8863a9c633edca27a3b7ed179f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29fa4e4827818d6f25ec187a175ed77c0f30383c28dac47b39a08fa5fc8d0e605cdeae9355d5503f3a7f254aa2f69aa13854f39414f45d0a878b0964ca308a049b0e623ab3703b448dd6d59c65df27a9798a3d991af5c12637edc90b1f9b7426a3b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43ad6f9398c851b54780690df71fa49ba93b414a23b4f4dd53f564b476f4d5a7dcfe2ed8ccf503a494f030f008d0f5769d22e88626de6fb75a2ce2d11590549b3ceb53b466a9f8da570030dc62b12a7302bb5ffddea0061dad6dec6b49407bdea7c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1538c78c98325877a9bdb81e28b226c913be5bce4f9cce379b8ce1f5a74cce35e0e1698dfbe97708a2fca1d57b1a79f2932decec53d8fa13e13018e91f1aec56aa68f7a324df5b446a6c47367e85d3e5d6b720ab663e6ff80cb41a5c4af64fe8a8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d239cde626afe43dde761e74349f9766b9b05011ec5fb1abfbfb6fb4e27c16f26e6f92b65fbeb2a553d138f2f162d5dbd656d2acb14621fbb11a36120c240f0dfd94211ad63982c49ff5b6653b49b761d2a5706928d1661dcfabfe14bac57a40345;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h616608da9ea71a20555286876b01edad2861e81eeb00e84f658ecc6a76ecf0cbcd8832d62f185f8d3247c7a6127d1f18acef750f42b92bf8cddbfe76ee07f36a51c53c5eaa87ff6e98b2551dd0c734b5ac9663d04f09e9fe3549e32b28ae580a1bb7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a0cb24109db6ab9e91f601a62f2564319d12f748f76a300c4fa9f9ca105868a995e58b67a821936d56f05925c3650ed42f0edd19d34a0031cdca453ab0eb7d1756e5004f2ce2427656f48a19c0ce305083f23f6ed8bf51a7aee65fab61c329120a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcacd28cc5842ae977eb40e615c57cda7cac377ccfbb80052175fc85531e38de3a150a3450a8dc82bc32f1d5b78e0e8cb291a1c6df27c20f7dc9808e35bddb57f7e7badb29a67cfa70ba6196ccadde1a8412bc8cabfcf0ac5b4482e582d1ba74c99a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf11664724245dbd79438d1b350182980c2bd6b90cca821e37e071d6b32561f7b9584cc8073155bc4c8f2273ca737fbec193f87cd7c18870998ff21362b19cf49715a08e33bb04627b487e96c2da4a71ab2469bbcbb8b636dfeeddc759e6ef31122f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf98cad6e7585e8217216d2727ed0ebc25a299d9cca3858beb360836213156dfeecdae6682523b88dfc63ddf5dad1b1a46f303d75cc8a034ed0421825865f6c7932b339cd4812df7186c25738111851c275a4ba2f27149d615440cd94e9c5de8baf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1465d733ac93e22117c67ea0082370f22335118d7e9f4908bc1df7bd4a13ba552bfefbd6e3a63ca6b6f7e31ec75d30b77a7230d59701e574ce9820139ebd52951df814822bcdd653bef35a97e632d455b30fde836f69668390227d896329be2abcc7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h780ff1c9994c488c3aea700055feca398307c9752aedc4be5528d9387b1895fe95e078c961a384246eb3ba827125836f7a1080a563fcc3de0a63344e2d3b4f6cf4e92198e47ca72a74dc035cd73eaa853f83c0024714b20816c43d1d18153ff05440;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d53f9a6a33e112101d69a48ebc8af6fb78e2b4f7e0fd6bc11f6d0020ebc3a1856cae28478d839aefa28b70df54db0e629735f7d8485301f5d908fe5c1848e9e1f323d847b12c1c2c6ecf44b5274b60db89e1a89452e5fd9f8098c10d2e61c8210f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef5e224170231ed29e39d3670156f1514a77ae9db395f5b0e68a3d2105bd59561a0de706fc884423b8c5b571ef31568d730a7414f0dae3ba7c6b53ba5024c53f22c04e5ec5a302ab058e3cbbdf938559aaced0dadbd6dcfd7c802c7eb793023d94c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbddd1cabad882cb2d0004e9b24209fa52b840d06fcbe77ecb854ebeaef931ce174758f690454d6ee173339a7e5e52b0ce8fbe53b510f6b8dcb102c16fc4dcd5ae07c02b7b9ef7f0fd7d70d6572b5d4d42fbd5ae711855111538201a8feb64a489e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h478260daa0a0d6bc355246f86db0dbb916210276104cbab1ac6878bc6640bbf5d6104265d2669abe61f895752c4e581ab4dd8947f545f539ebb8b7dbe3c93abc7961aba3cce17ef211a72adde7d540d9c955766df9f1beef77a38e4fb8666f4e39f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ed10ec4c3d34bb5831bd889ccbb4d6e607488c78bc350541b2df9713c24d6a23c0fdb4e3d4b0123af5ac15b8177e3c279fbb24174316c8eb7316e6ac333d1e75e3a45239c2b9ff0bd76e15a4684834271ae36954992296f6c291dac4be00f83f868;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heca69b3c1c8a4bdefffeb164288b980c126e5a3d2b8f37a3a43df61576b774e2b9720c63e6e63f40f1817890313b5ee94d1415b6180b40fcb980ce221f3c42ebe152fdc7a917822a70dc8147fa9df8ee69a874847ab9d819d88aee1f517a72113800;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc09ff1b1025936fbe2867e0b1767f72bc4509fb9e474d1ad66b3655cba791dfedad59980f56e870472166d7355f367ce5ef34d02dbd7d1d032f75bd5916feca6aa2278e2e4027ad7f776c914dce6450636a3bca4829c6647817687f16080a00e3dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f0864394c6091e274eede33d58ed2ce8294675c716f759afc675026794965cd90a2d1ab0f7fe58db4293cce4fc4acaa8bfee597417b52aa064eaf263687d7960e7344d57e700a7f876a6fa96edc5b46a402610b0a076e21859ab353f585dc62ef1e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b4123cdea2ebe2357b6599def5508f64c0ee3b866210d114b8ba53317c1b853a1216600b3f614c4a1e861d2f745353ec8f64f030be2a621fbc590389edab508b2dc89d9c4ef35419d06aa7dcca7e4f5719a7fb788fc530bf8d9d8b9d2c8bd552ed1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9155f61d85d4e89f99accf2cd0310ebf84b3bc90a00cc43cf1ad6037cf9f86b36430198be838666bccccbb14fbbb00e682b00c9b7a0c72514b03564a4b8c2a259ad1eea5493628a7dd51052e73b4a260651e6ebd00ad29956df0138bbdbca2e2da35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h660a94a9f1ed2ad288a5d1e72c090bc8b6b6c74fead0aadf8cd6090501fc2bb5ad451813b0f0e2a8f060f885abdd3c91951662dea9722bcfb75cb3cf43306fa82f99621378f67f49eb97c1a7ff9001b949e9e082858a612b1250f1f12109ab767422;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cd6f23ebed08d53802f3f7c211660c9832bc3d6d13019ae8f2cacff81ba460d546f70feb0f0136999169e3f6db6c501ff163d7622a384339867a068a31237893e74c70b9b4662036e0686311858a38da622125e424dc0b90b6467b555f93c9fef48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9abb1b959452e60c543afe26834403df7cf242565d0073840c12dbda9d79a3605fdc77dca1c784731bbb17e88a4a9b8370fdfc8f00d9bad721cf4ae459544b90a91514e2171e34fad10829875c0dfeee715997c74ef87dfb1bd82f31beca9b60374f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc5714a64b3b1819a1f1b415d629a312c54c65e27bb17a52e5b85136b1ae451d73287744053ec85b67b84c94447fa0e9b05083b3af2c0654d87375203a36f49fc64c9dc913263135ec593670e006513f587073121133cd068cf891ae2e6b18cad3ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfed9d2083b2f97184ed4ea425d734a3cb37f8638cd996e705a3f49c89d48981645568f39a4987f2f1db8ecf9f605d88c8af575e60fd55050f0bef80ca6e4e385a128b9098a6bd3b5bec323c8c4b2067f5bb34c323366209cd7f3d9b5f8f5a94f0a6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17d38add4e12c7022a4824deee9766d54214ad0b5eca442734b1efe111f0703fda3944beeda9124c3b5f2091df2689add9490a79a307c701f5f8639c7ee48e7d4c22e9f81b5ae2a081e15dca5b1c39468b707c2f0666fb8c2da3a8e8505d26aaf885;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8907d80a2b1a5a2a37f058ec41d49cf03bcf058b2fb1eafdab3c590aa2f616a0b865440660cfe4335dfcbc1b052d5252983d227d15c7668306741ca96473d603523791ea1e51035a3db1c90bbe2f740e407d2a26b0bd2e00424f134d30885151a72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f10923cc0e73bcc4feb38e0f437a3f4f3958eb2df360d462c749054028822772bd2c7d5b5f4f76a7eba8f5f2c4bb7986fdb7503e726437464e7294bc1f66d2a9529595bbf9b85817312d8c4bebe7601532f526bb3594276a9a2c1373380d72cdd2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2569145b23eafbe98d49b4b56cc28a68030bd50d963cd460061cd113ce22e60b706d37da88b8bea10b24876087f1c5b89384621130b3f7ace46731130c7d538b190c426fb8cf50d11eb041518e4f57a972b204611120f9acbe25b410da6dc6716e6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80762edea6ecddae90fb61d20586ecf8713888d72d4683f5ed2d35b8a305d5d813c844cc55934d69a6b11efe2ac4159d28595b414c898333681cdaf7b7406dff85a4e93d6f0fcebae70e3792f958731a05153def8d1cdab29e801eb9f3985f8f7c74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a9748a3fee69927e42d940aba592fb8e9317c6ae1a231ddeb064f01cd3553f15a921f1da25522685d22117d5b3cdd1d0df3a5fd8dd3c013c5bb8a28c967d61b0e2f7c992eebe8582414385cd64c444b97ed72a0f3ac6fd356cea4acfb41400d04ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8b60cd13aa3dfdcbaced1bc324e451d670016b28efd751982dfe1ac7c46b67330e5ebe58ca54a2cff98d89429842b9ef73100e1e59531c49c4003846b070040290db0676b4a0f45716a72ec651f506949a44d50acb12ee09cd1cd0329641addfc1f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd33fef94ceecd6199232c7d40895eefb5baaa5608c781f1ef1d352f52d82768b0ce2c20f7215bd3a69984b53ffe10fbb7d096e412bf2def92d800678911271b380028a3bebc8e9798d13f46a36697431222b27aff4898b5ebd7b794a9eff8222f80;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff912fe2ca0ad21cd611fa9360556a0ed732f4ab89deb7f42cfdf388f75d2f247c76684bd42c813993d5af8eb6bc98d6f1fea0a0c9e342855d2064b38fbbb825255e6c94b13c7bd299675ff054f9590928afad2398e1045e5a0e1e2fc0bd1a9f749f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbf27ae2362c36446cd1450eea3d8b828f10fdeacf93f7457a1ec618b0bec40b07ebe351a5b3f20800c4ba10bf05ad83ff3c6750224c23d009af57adbb6d9ac335007df5fda7b90ab133b715d4d997a1d0f2c916779d3709bb1d70eb6e77e6001519;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0bef290b914c5d14a6720bef4182080876aa756dc8116fc7543b411d396f8d11e3a09eccc63b05726e7bfffc9aae586dc4ec714be3b100f2c3f88316ab09448b39ff44eec5a96a89395fc8b4652f4619216ec666ed88763c61c98e4eaf0e88841e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cb878fd199eb5f8261a8f3b40996c2ac43881e3f11da93d77fd815194f4a26172bf7e0c53c159da8f34868b41d2c8b5f8561b990588143e531027a80a70bb530e5851a6d9af79bfc7036c057f2e3b2c69a271776e26ff9df00a4ddfcf1cd8175632;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he13b12be84fd463de5211364b5abbf4d89f2ced4b5e02d71856fd85d4cf166f6700db2b760b96e155dc592b918c57b207bf80b4429da8e97265f990aa730c272f64fc8a4eb5f4ddc879da6521b4bfa207f842ec9099d36a84b8070231ae22957142d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e2b8d23716aa85e943228acd394bc06603dd156f7d83250c89217bd61128bc3594ee56f95b37511814a5c67a4a2580c6d5e589d69aff10d403cf962cd43b654e172b4a15031c484942207847f1956e5c0ab955968d49c5b185da6fdc2a31fdf0841;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e2a61e49cd73bf9e01f557a4175b1c188e8c5bd2dcf267cd8157c7272964068f02768f55841da79e661b392de7846a73550d2ad28fa753e899d5269541f7eeb062f05f9e893eff04a3c6245b5bfcdb51cd81acc3c3b31ab66a041b623623849f002;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb73a86c3353c2c015babdb8e60bce2eb1472860b2a844d69c90305a74b02afb57a93c1557343a914d74b26e2db846d0c92fb4ae23872d1123bcb0fd8d54f85a1255a2183a5b877bc226efc8975670d20c7cce292db1ac835c0eb626ddec61a8cff9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49b21d476ecbe623d2b58de1f3f4b96a25d0ada429a02a5a63303945554a717a59233e276fae4936805b45dfb56c62ce415df9c8337f8c00e63d3c6b58c67c86f4b86bb7bacdfb5c7d3d40310519c6b11d3e9a8790c5f323c88d1914eebb380987e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dfbe8d314871ce7b8856796a9fc181032f3b22576d1331ce86de4696b205609058c942e4ebd3e5150fcdaed982a5abfb802cc24dc050c071784382b640a1c50c4e0b2b4df171b90d1460d7b5f9ea7ef22d341c2e52b7df20bc6fb341ec9ecf38fdd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a4b191d7da2fdc748de21d3572a8f36526b8f0ca73ceba60cf3d650486818081e8708f9e04a20184a831404356d93ef3348bbfd3d54f17af1e60d52b4fd020af030c1fb4ed2ba80cb2b1936d30b51e132868de1a509cf9b3b88c9d7dfc05a148d9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2644a9f01d92ad0ab3e2421cd1ee2dd6b524bc71a774a70c54948db7bfcb34a88b3564c1856e3c26fc58975c20c96647fd72ca12d75547acb30b5564721bcdf32293d40d5f945e368868970aae6ed8248f12da6c22d11c2d2eb4edc6056c3fd350;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23eb4c378217465847c5e9362d3297b57e364dc73f6bc6bb9f01d10a4567fd79579983ee0f91d0ebcb9db830ee59aac2b83277e0f02e0d8de93d508b99dfcc533f5c1e15834bbf6d1b349fe6b50be98f1ac5699c9cf8dabc9ce8a004f2cc3eda179d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca92170f25b6f0a852d7aac2d5f18f9e6ebbe6eca35e39fdbfc8c205e4d234db4a391e6e50be3a2e369031b4a09be1a4177557b1bd12de4a1d0aaedf8bd718add38233893590dd1df09e5e9d0f2b92a8e8015fa35167d33b2163af2dacda4e0ac9a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha31252cd3611fa09178fe59f5730c76f7b8f50e20cc163d18ec5f3d92733d6511a93dc9ef051e9129262d5461372a2ae24d842fbc87f97864d14b15d783cba8ed0a25e1ac58acb4622dcf83399dca3c1ae23e9294897ca11777c221d102491987e75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h584126c165ab8cd67d275a5b065a3b5012935852ecf53bd070bc71ee797d65d2f7aa32c87cb30f8fbfb640412e7be4a7b49d88542d61fda570f8ab10b823e815feecbaad967bbb3240254a9954fc4392ba3a118edab960e14c857b5abcd8ab5639d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc84b7086d9df70d236b69d795241e374e175a7afc63a2d781eaa770ba36908cb73d419b83ace5c62988dde1a9bd956d682faf3fe1b30e254009a5f726aa36e52879306dd2d07fc8ff18211f056dbd9c64c7a1f5051cb61bf297d51e797f8055e1863;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed4849cc3d59db4ea789df9977a5fd6e664c154079e3689e018f65ae25afa0da0143a35f0b5c85613b4804b3bc34290bb46bfcb08dd927bb84602b4afde75070e92a8d2186b0419841fd8a2b03557846cf37363891ea290b40d45f39ba8ebbcafc5f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcaaea8a2d6e80727f3be0bda54665c59f9925bf881d078850cbf9b4413ad9eb369bc71236a346de9ee156d0f4082c655893ec2401aa680f43f8b99c237bffc146805db2c5a170276209b39a56f12ccfe8fd957e3c9663b4c96ccd0812b1cf1f4ae2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h278b03b20a436eba70461bfb07faaec6fa931af3b8a9c237ce4ddb5a87707a46c7c5474f95aa2a1d11400a92dfa197fb9353106db30ab954eb8d9aa7d52e560486651b3a84c86a5b9a5b76ad0cb8f9cf49ee562bdb0c0274a60975a562a75570d4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69b63e3cd69ce55f5e46ec858679dd8312358b43d71c7212ecde475891154b377ccaa6f6423e62b2e2dcf1ab1b1db30832a096741c1a1927aede2e10534bf04a55955dc0c3e459c5b4e41cc81790fb741797032b1877790ce8391fba83b3ce92cb07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeec1217b381c219e24854293ed56107894db274682b4054fc3d2b73f21849df34a8e1ed63fff05fc202b812e770b4495d1e6ecac31bdf97d7c21e914a8a3969c91c7e9fc1d078c1394605a5f973f8fbf4f43f464ae6364c9a07825f4d0919103582;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2350557e96afa896f76859b05433572460d4498d49b2dff56bf364a1ab62f83db540d4149eb31ddaacb0e662f0d57dd335c9c0ea1443d5d0773f6c00e9c2de760a29c71c58d69cff218cbc0764705ae23ead3972a22fc338ff1b424e1ee6f312a004;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d374af658b03c8cd9a0a31c93bf7ab00dc6334a63090e5d8921e5e773b36533a8499ec0da55a39c323946a540258c4ea83c547cce956bd6f86a00ba8c92b9a7cbfcf391727a98b4fec63feabd97cd0970a53db4550a4d576be72e150f0168c55dbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fb60883b96bbd562de1c309ede05895ae962e30c31eb1d1bad605f2d738a2af8471cd5821702c92b01b31028588e1c7af31112ab32bcf7986064845682d2c51d9701f763b4ffd3f91da906e62b358aebbb51fdda9cb4f5bba3b6774af04f0e6c3eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfad3ea5a422abd4178545714ff604b66acc090c159b24a17e42837f6accaa1a8af79ee945915c37c3e0baadc7963a6f150b1d347b0ca083ef5433ef26719affbfe5e720012dcb01d06436791ad9be664a0f84749af362b7d7c290867d6ae93f38e33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b75efee2e3baa8815a3357791fa8f53d8ad542041b44afc0c070a25ff8434acf8b2ddb8874b34f8476b4c6ef5283af380aff3f9c691e0f861dccea77f25e45032561f0d488709085ba2833506c93d44fff1721dfb198d51a5450c46be14b1462e27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7de2be256d65067ba69ef9e6b5a10dfa3a93cf426b12a5bc1b544e672d2722bc2a9874f20e4fd2a1d4f6ec50e6856f7e01354812c737b70c30c78a849919f32822287f9fce3acb5d0754e6b1415ea86b870e43943826fead219a387bc0156109247;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d026706ea17f63fc28a9ffac12264a9b04880f64d2bd2d2a97f8bc1bfb961918cefa209337ff7a6f9c47b1c0497cc28e171a42c34b05eab13545fb357356a981aa0902fcaaf28a021ca1a2d75ec44bfde22be93af73382ad89028b326e4b2ed16f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61c42f4395cbf3c94b9e300acc4ac08e0bbae549221da258a462aa87ed72b68b09f86b9da37e1796a6dfe4124526e2e28d470d702296143d33e466a29376095d8fe681170b7de8cf0edc70f3705b502f0dc6a3c66dad916f750f6e7b400a6f128a1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h427617912cbf4d950e06276857fa76d8b05e19d1b69175de2868030ba2981e8302f3613ddf74affe789b6ca2f9d1bde3ede5ceb1be26af2bdc0fb290766628180d78aa5c5e273a5fcce0797d0727394f44e49d7718fa0548e8238f64ec0f00e7cb37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18afa8f926f3a3f213561c21f103a32c10c050ab2aaa6ac351f7d674b9d69fa9780555c14a50e260c14f187ddb43cd537523aeebae04f6183271b4757a93ae73a46c991478400ee418f7bf2cfcf991d774c4fd2e53c9a661c72656d4e600381cfe49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h457a4198c91058b21073d6d7ed04239409b46af444866c9fc2dae0951a8db1f16df7a4f54b95d7341e7d03ccb5a9335ee326f205f02ef7e95f796925832f642e750deb60522b47e7777d5bd1d7c4aa19fa694869dae666ef775719e2c9be857f3d00;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5339f01c6573ee242c884a714323aaa71efd08b2bb6ef6ec457ffa3a6b8bf6065fd6e8342474eb530d3d3c37748c69b1ff71742d214b3e702db5b87e1afd35b91233b23b367804c82177e6245675a970541399f21fdae581057f639a40b2b5dafb20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe0bc82565dae6be04ac184c964605f667ac9092ad2e5114f8ea7eb6833d84da0c172956894dde21d73c3a2d199fc947ac784117a523912e2c8e44ac8d9f37b444849ff0481bb2addc4c26ca66695887e0d058582a22bd611da318120701a60085af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h195c51f53980993f50273b3785d3cc750d90dc1b16171fee1b3bba30cfb91f6a9b903b1e8913262e0a7d6db3828aaa9918a58cf6fd6868a283ac62849e078acac4f0bca2d03efaf6a40e942136707b6613c0499acae083efab6127f2e700440b7a72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5df69e178c406d75e3f0c5bc7b4777c5b7059a479695a000dc600ae7c02ca2b85cdf69275d6a6a9eb84700ede3296176eb6cdcd28de797b9aa5bd13e8d493209eecb2a7cfac5ad066a440fd05d52836c4b7c6bdb7a10981375c39a0ca101f74bb8b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58f60e1fef124f23c36354f96b1f202126eb151d71dc1c348c536a729b6a34f96bc78e57cb236f108589ee8ab74b267ad93ad1f5ba3244346eb24e4d670924de66727d2dd9e43a153230d33f90373722d150be1af05d81655849f71843783a3eeadd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1563144bd3aad0aaf3828f7af3676057d9f94700e399a73741316daab8f0cab34f5e9b783935be9c3849e40cb60e5f5c3ecf10f8ecbcdaddd93b457c782d551795ec7cf565ae382b0fe244fe014540db0a3499dd2eb2cc1e6425bd01272e69dd8916;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66d87007436e86fe579c8d3925c8677bce26094ac679bbd004f132c82be9ac7e70f143a73573046ef4c938843d2fe23944018355ad969d78524bb7bc3a9040df452509097627bdb1dc4b12de82b61e14f0fad9b9cfdc6ec425e9a5322c87c2025b62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8469fea98227d6a0bc55c6e2b5921fa59c75a1b0b21b2d6556190f1bec01a88fbc7a8e7fdf08ff080179ebc7a416bf2b40b2da353cd3def04dcf9bf523c27f2cf51ea797fedf8bba1bbf990ca0a2a6ca9d779685d8ab8d2703ac98ff5fa278629d11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe108c7bf8169c185f2ebf946ba22e44ebbb3cc47756e08b31694d010dbef7f12e7130ddf61c769f0097b9d6549a031bd4b9c6fa97b9dc6227296b7a8d5412662ebb88cd178f78b89bfddacd94a424f6e8cd75130ae466e7c47e121cdb4ec4ee29a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf39ddde06730c09b71b1487d7d619b6c45f9b9cf33767bfbc8a6cb98074be5376569746fae7674e474fd02abbcdc7c7aeb74fa40093af9a424a871483dfac8ada57b8b0a99be94e8294b9a34622c609ccb22e375b0476bab12e0f7a8431057593fd4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h155e2452511c1a3e5320c3e28f8942518aa6870990d500bfb72f48bf4c69d84af240cb884f822bddf25d252d537290082233d3ed91c6a81d706044f4c37e08fec527353c52ea809ca4e67447a6af9bf848c3eb0a5988f9592f4d0e15d6188c00ae87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h371aaf474dfd5bd8bf4dd976cbefe0bd9f61ea5813d726f7ada99bd33ccb860ba6ff7df8103ac4a69c521714ac55ff1e1b91a7634e514635ea1f82083078c598dce0b6954ac01b19d4619750db222e08e795b811152cf86feee3e10090e6f3be78e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68570c6debc5811ae3cd8bc45f98833e2fa6b5187e4e433e61f2d5d17babd796ea36a07b6757702b79520a3f4c67411a4a5ebbc9e6bd0639f9ce27c1439d0625b82d8edbdf538a456f8eb5bb1dbb1df7b9f7309884359ec9ca035c2d8c3b4f4ba6bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfae523715b53797a25b370a1fe04a47681041c8b4fe50eefadfe22536ab5e9aaf970a96efc65f91261b7e2d8dfd9242e1bd9cf5bdcf44323b5854e682bd53c43c30aec751ce6c04cbfe21ffee15631ace5d2103b19d97c86d21bc4b1acf1bbbd535c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha54bcdddeb598b01054ef2f0aa50adc495c34945ec97c21669c66f46626ed24e595336bfd95ef5946dffa759fa503f68019ba9a65f73c22f571b26ec1d912dfbcc00d0a827e7f28fd96043238018c1fef95ffff3f34fc33bc0521cc0cda2475e359b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e3a01a163a677a960256f152a8bdae102e9056abfb1ac415c110f7510d5ef8a53a9e5bdba2bc03929939cf11418080e6bf018d2a245f82db52a820fa7dd9d2d8d8c6019cf82f4c2b1a14dc0b6d217d4f3ea4e739289aa8c585401e3d84e68f6fa3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d41c5cbb02283d5d1f8e080a637cf7831303dec0ac3e7ea80e1fc966887ac855b4b5dc721ba16b9a91507d2a8d428e9bfca97bd489ff483502eea5dd2894a8f4e4d9a27c733a03f1b29eb091f7469ee35ca7e4b2b516b01be254cec0a3a68b64cc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2406364aa2cf7a89b72610245074f8ef046fd175d709a4f6da5087586fe09587f611dde39950996ae2d1b707b20ac2a84cf57fcbd243037606fd90639b157e3f2283ca170a093047888782269919b06444cbe7fffe0d5816f873208dcc49ee5f90b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3464ea3dfc38587a62d4a732e4ee0845dd9407fce28042ce6ec91422d9934676c4c9e0e349623d6fad553c78f52e835f3cc62498534a423989ceef8d63465a2bf18b684a29ff2fd1c5b87b3f1077c17d23317cb60f86d78ed3fdbbb51ab0801deed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca5b523e9c63342d6dd36216e29c9fcf2bf338f895e27f0dad98c33636e0dd74782089e6a5e1c2fb5ae7830c76f8d5c4d7db67f2b0589e63ea2f23b5026f28f3bf86a0948e631d31fc5d17ec6950766391c10ca9a219c07a1043bc4406edd96b1324;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h292defd302d2c41c894edd3cf6093dde39f267f46aa5a002424a56d4e3c401c843f2b16587377db6255133aaa5c23f8851e2a4f1ca2596f1a971f605653edde8812bb62e8d26a5ef441a2a5382e258d97ac7c1b597051b89ce80bc27db2d81f36003;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h136b240395665d96d858d00dcb8bb312c270158aeeccc7ad26328daa12fc73b8e5891627b851833db363d2d6316c8284c2469618643802cbb48454aaaa921a90d3d825a22cb5c892e412fb4139f018861430086555c2d16e10b98a281faba4082bf2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bb04a94030c7e74aa6045c6de218f18b3bcef80836763c90a1b0e85c58bf495622eb51cd96618eed98493825aa8734d1b6fd3fb0aaf0eb8c4b31ddc8025be023fe5af34cbbc2e30919b65c56d58c7508d828be68385933b40f8cd0d1860612c0570;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70131bb96145da5dd2ecab60df4522911b8edc34ad452543538759661d3d44e9106e06959542f0bbca22713812a8f49f7a088d2f74389b61d525c90573fc57292920273c10889cb74b52aa18b865f763082a045c4e4380906ed3790fbd514f4720e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71d82236d1a297b4fc4c66918da6b26bf971db86d38eb8afd00712829e4d349e3057d0b5710f45fc4980fed1706de24b8c6c2b17671ab224363410d50f8f5f8b79d3529f31e31f27e69e6404c63de9da54258a0124da4ddf11984b81766d63d4ce5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ad012c3030b8eaa200b0fccb555cc73284d8922088d5767a59a7ccec2349f891916ecb35eac0809b85b8caa30ffee289faa86fd4089cfc6298e759c4d1990090a0b83e6c6290bfefd48437ae1d4f65e392386f97f2b323fb37b100eac2b23b6403f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41a95603f3963ef668c14e1a7478035f4b9888ab47e6e9cd0607daf9f4545e33ad27473d0a484202a0e020d9e9829b704cbd7eb8d865956c6f4f5b36b6ce8d56775d8927e30027d0d0d7d54b7508437bcebaf05f45193a4564627c17aa8122443ae5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfaf4029a6abfa8719097440e3168e60c159ed666401ee57d249b226b667966d8bacfb6fbf46224721309de17c3ebcd5cf94e45152331e39598b1ae82fa78b837037af0503c2deec178756174f537e5ae736e4c8d6e69bc1c8fd86e1d01885b607222;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he794a2d295db48e4a3b735da7ce608cae4e2f081778f20c6bb08502e568dd200d7e9803f60775f6bfcae7661621270320d1e0c8522a9a92f4ce43677bfc06e89780847395670cb4418aab31ea856e181306892322c23dc1e902b2edc9faa65a29fc8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfce70d29b1186cf18d7f4af35ce71fdfa5687780ca3d11b23ac0f1a3b95ee508d4ee5c05177e6a54f08a7fa055f63299f048827145210bd1a4c30ce44c92ccc81a1ad2d5223e04e0e17a068d5eacb2441ed3ad0ca518d19c4d93c96da39e497ef95c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ab49d976971afdb551b87490307326f40aecd58d87c843d211c4d39421fc620398f335382826ccc2ae65b8659a101fa83eea726395d4cb6249bd7de5d4c6aed5da873dc24907d784873877bab23b5ffb0ebcf1d60c9b78372ca22d4d097e2c88999;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cc3196a17c34066ea9471e4aec10a97316a825618fa81425b35160e7b99f653c75083b3d7fba0692bcd2a910d85beacb0afab11197f2650caaa46cd5bb3a169656e8c50d32ddb50feb0421afa00d7daa60858bce8ae5cc09f5182432b6bf8ef082;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85effc5c997dd71fd93afda23da672864e696044ac048cd901d1757ca5c554180ff557ee189d4455ac3b69a0f3e2c4125264c70cb7b57881cd41eb81b9a7879b1682c46f1ac24e8c4e892e9adceb1d7e651241a35816b6246cb2b538dc208cf3b7ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9af9d3efc318e591b3574af47cbbe061d977136526b0e1a4f1705c2d527e5bc72b0a759b151d87fb2326702656ea7676a2802aa0cba763a8a15368c68797a38c2ccc1af366d282ebfb512e45c08285fb1d611b76407f7def6a724fd75583e3551bb6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2f61936383a85a106cbd4ec6aaa6536e317b43af3ccbb9fbd46ae2a7bb31a07e502e1c6b93f451e5412ce1a643f789e974edb0e99b8b36eecc06c4d4312ffa3d9fa1075e8479ba6ca3c585f4748f855450c160dfe00e6af2be4fd097a7ca8509ae8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h803f0b92a537cf2f7e48d17836911008664b1f2887cca49d191afdcc507dbe7c71eaf60528b1a7d2bbe8c25e88035a7be7e4ce496255644b4450d5077960c504ef3a46c314618f72946e76b265faac0d286a2b91d56dc6cdc67810b2f53c55b8f247;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96695c235ccad781d91f8bdeea152c325235317f7c4ec9632abeff3ef18fae4eb8ecd5ff58bfc030599b3f892274c9b03c298e512c040d9c6e14f5691623ee91bdc101c0f4540e337f58e90cfa7d3934b2707da45c8e5ffa2210095f60e3ceaf5944;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h186a06ae3070cfd66bd502c9e5765d50f7ec8587d9d3f77ee8960518076451108335853baa0915c372ce68ac93f19658340ec2510656772379e695ae20fd182cbdbf60952a7958f5129b6d921a295912b5e93356ef47f724883bd42d9327181e09e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f8567b94062fc51751e9f1f5f2a5ed675ff26a911fe416e9c80b932de0a50c46bd4ad5eabdf8c69aa4806bc3c64a5f2f8f53b7af5b22b47abaf5f2551ce94113af980dbef9449981443f39d8111361337c2ac961b9c80486bf60ffb1ce19a4b425;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14e80fa6bf3faba212688feab3c6179b7673c8728b0cc05d9d515c248048882fe8a481bb54e248e32a052f38c8307393fc8b48d546a2ba1831401e1ec7b1b92a313f8b898f9518d379dabbfb61cee8f6ebe82c6d3d6f0c9e755a1489abc8492fbf58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d8cccd5e6a4a5758b6ec57704465f7e39775430558a28a59c9e13e6b110c5a97082f4983be78cdf2d79de9169d0f3f9dd5642b6e0fd83235c8b660f0108c568cb279c92497c037cffe6a2c395ee4fb313f6222060e328ebd93194c4bc29d4ca3f0a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b17270f47d64798e5ef564475326501e260c8bec6bda128c99f8d634684640d979c46903a59e5074d5c5a5c345b4f7729342c4771427872ce6ddca547b6517250e5feb0a806de4811603af54f6dd47491904772f0a1b58b1ea91beaf75b1322074f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb84b7e34dda81ec680051fdc5a2887147cfea7d4402a924877de6462578705424675186aa46a1865de352c99a65eb74b6e128671e0fec4d9df6d00253c37393f2239f013bb39a26a880f52a12159d4b4f557eed421bfccd194b57988f6d6fa3ba3b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b4f594cc76dad79c686b270e44a28dc004c85259f1c4dd13e51e0407552eced9482873fb424db17f2f3f5a6520f03adb064cd7ba5ce56f67be0bec3f224a523d940a99f31434e348fe8bff9ef75bb853769c58386063afa76ccffb9be685151ca01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73640c9cdb591d507322ec5655e54ded917cc6426b3dfccfc9bc0a4cee1160dcbae93a9a33e035f53a25295310dd52fa1fcfd63f18b105f3dcf576e463b0b7dd26eb291ced099ffb4c886304fa44e635df604e5fea89b5331f88fa1983e145d54396;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a9a80b2a122c64337728793de808cb41f0d4af6f9f3329fe1f562c00b05872768865a37d2d853c38f41bc1410adaa16653b6bf1a6167b9c613028917ba900a26c727e5d058dea94c9ea42ee1627e5ee57cd0b5043636c3f22d022b399d4ade49322;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2087d659ad7bf24e197c7e7817a848b67a8c617dc3eddffc4af32e5f0eee8cbd3b23f6700d1fdc863a49e2cc89859d5c7e6036421b52e48446a7a9ab261e9249344c938c978987e4f0139b8746f5edd36abcae7e47de2bdb91c1e4ddbbf7ee7a96ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e7e758e6ce9db4e39bb44e9cf40fa229648ce5963d14cd59ef0d98f4fe8f4456ea551e6e7897a043bd9518abb01986acd4e3a95026b55f186b130713cfff98385e005edd90f2af7c815e1b991a9826040cf40b7469ad8fc3c616630d56eaaddbb49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae2ec8e10a999d38e33283643f7ee5f683e88d4b5b4e921bead4c3c83bf61b91de04c715960e3d468eac326a75058a9879910c5bd7d0852ce2ba6ab5499ed52f500b788ed9c8ffb40109deeb514eb3763e693653b1209c8ed49b9fd0cdc13170988d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h217d9229ee82a5bc68ec52ae6301550ee2d0bf5167b61b42b48887adf5659125b782b7b3cd05ce9b6184d8b7e1e8917f26302c244403ab3726f62daac2e907ab576183fb9f5973323208cf1beb922a3feceaf805a3f73af4822605e688057f2db040;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33299f1b218d98d3ad53cdfa7bc6f4db48a537674378d0117e7d171516bc5b88770ba0cc25f52becae8077a707a94f75a604b7ef0a24ad2450f119f666081d838c849e65f40a451316726c148a77f42fe3ac51466f1909d281eb37678312c19da9f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca5f4652a17bef9ee18754f40d7c73df408130e2daf814f56a07367601c1139530178e672b73b5cc295ce31d82a39284a8427cbdbf845836b088cd6e811c40ca4545b0d7a165fd9a2e6790de4bc1c560288ea007b0581545e0bf4eac3f5b4e5826b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5911c6881c5d19c12e50b4a9f72a47fd504b4470bf1522ddb84540a692146e75ee6b1cdcc0a96363101cecf9b1403f9eb9bb1486a1c08d487af76882fc8efe9cdfbb0ec4ce9f7feb7aa27c93469b021c6806edb8f93c81ad9f94dadc096284d90db2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f82099755e44b2d8624772f496ac57770d9ba4cca56c77db7dd66cc6391cef559b3b5e7c90194ee097e378b1f9831ffb3243fcadc01c45c5462ff4f792943a63ab3c42ddff312df571ab800371e5f9bde4a7ea2757b4a0f648320c9e2a829c013e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53bec0bd6868a8d426a9f5f8d1d0f20dfdc27d8198e087c01c29e50dce28b60106844e6ac794e09e703782749393a24ea6eb581a5b6b9d02ab4750f71bc1c1bad7287670e9f8faf011e6ed5d565c52d0489ef12f0b189aa47bf056ae7d0c0c29993d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58a859bdb9711b646ec1c71fe0ab7550a08350b2ddf1f479ec073aacab171a9ed0fb40cc48e39be1219c86956f7fc9fc55c0050847e450a4631368ff1514ef832f83c3c339449fc896bf317b6e5cae2dda65971619f3289a3a6674fc6e3f323623a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb90f77e26f9e78b10e84440253878b2c68785ba8fa78f44196d5a1795c5829194127f584386ec67b4c8e5028880f81fa3e014e9011b6d4bbbcc7948d3334ffaef498a5ffbe1ba95c5d3008bbe8d0c3495db24e8106f7079c4656e438bb2df746e8ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1c575ee2a48bbee28554586b799cbea3ce70dc033bab5095b90888156a5f7ed5cb8207328906a428aa9b165d7912ff151f1c3202c8514438e822a07881bb01d11bc9b94619d4ac773e5aa140103c1a9de76f6467ea5acb9f5432ecddcc1e17d8f49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b6fef403787586256c15c01221607d6a15ac3d495b54212af2f13e8c25b8402a8f8cc57ede2addbaeb772e7b6b5cab1849b29cb87fd638209462e7bab16b8667b334068fd10787c443304e5b12c8a0d06a6bb84243632a385a35f66f1f7042ccdd6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h839f4698508ba72720be1fd062bee28ad1d061925ef8e34a6d4019322aa26ab70f1ac143c55abb4fa51586025d55a18098a9c7ccf33058a071715ada7697ae9694e44b0ffd5ffb237306159aaf9e71a76550acf86456383a05211eb7985bc0810129;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69532412ec0cea137c24de402a86ec01a59fa3101e5838375f005affa05ba226b5179e4f26452149dd3e3ec5f1962213fb680436a1c0464883b6026697472eef74d2c14bc11611c4cb4fb8650863550d2aa45e2e97e0bb09d770cb441d95c4df16ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e6ca64a5ec89938ef3dee860af157b3d579f231bc3efe76ee6f846546e083b783cc6000f68e0a7b60d93e01012aab3bf39fc9b9ebe9c86d276ade84014851f673e9386cae1ed302f245ab131b26dd4a982b66be71fbda22de0f0926cbdbb4cd2e5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1d5201c9fbdaeaec6a4a4e6b115b657c215b986fd66c9841fff67f0d2b7d8818b9bdd94561670d6fe6f4d5a4cfc5dbb8a4e6fc252297995c10ae9f46e86ef0e5bb7ff0749b39074999d1203a396017c3b14f3ce2b1e9870188025ea38f4f20a38e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2412591a24b8389c33cffb05ea2cb349b88963c8cb7078c8e37114b43cbdb9b709b50b55670221994499fb66083a1233d2c06c567a23f94f8ecf30a80670f5f0e4f308052485627e187d1b718016753e5dc057f028a9319221c46b6304b7d73703;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31f51a8446ed4430b5df2a3585eaddd6e4693f5974ab44412f9de92a767b7ae2a4e479f4917ad288ff0ce47579d208c40488b46a855c39f702814f31c5c01054bdf32815e6c672c3aac81ce99e59f19dcc81a40848dd1293949fc356cf46ac732b9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ff2a073fe383a1131d55993a5795045d91919da8c2f71582207a4ca0c46ffaccff30286fe9f03833d7b73c54b6e092f3420a6b4dc38772ce10a55b10badf56e575dd8272eeedaff6905898279c262adb473ed0190455b4bb8431703499f2482d9fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5126b97789b33629d833ef3c86dbb32e3e351fbf5024fc143b11fb55a65d8ae7c1190923d45049c259eec4cc4dbc9692a2a7dab1696b1c2795175a03a3d80a10eea637a5a80071726bb3269fabfb673985df5a5e79116f464b99da52cfd10486620c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aa46d88647ff359a0edbd6cc66fb606590a9588ccc7797dd8e9b026d8993ee2a0ae3497f0bcf320191693d9367c7fd26f52188ba689f16b15339b2a73f03e875406d70e6604cdbbfd2a8cfeb9ac98951fd0810a2fe8ade46e4338068656a8cd7207;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90cd3fbd1850b378d6119f10a54dc3dbc7fd9e40a7fd36da4c78f794183dbe39984f87c649e0fcd9662153a89cbd262b5002cfb1a49a3ac74b3fd08694324158ae05775cc171ac739e3f12a9d954cf31e7d24c917888dc465f5ec2ea53fd96160833;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccaa0b6f7800ac59525fc042d76644e71da7c4bf436fdb9998badab4c2d0b154b38e51fcc17169d9d3ed6440b006571a0c5b6266321d04afa0a2dad0cf3a74aa229a8982478feed69494cc21eb214ea925bca05c01c0b98c1809a1017d250e46545b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf16b3abf73f9aeed73768cd43c5ca787880113e48c0380ce448495990f8ad90a2b2c7b81305c139ce4416468c975ab5a972ea617dd0d52481ffd160439eea9223cf5ca9f27e317442768d39eb3219ad6dcabc2f1aa5df761c99e4168d7da04e6f91b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9ef642bd2440eb4a5da25ce255c82ce6d41a085308b2d32aa2672017b7af566ddded973be5afff3bf2851aa97bc568c617cb2aa57ef86b82ef310bee1ae055dd44dfb15cfb9989df23894ba32775761d6c32247eed955b794063c90e9bd70b0feb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he27630ac5acc42b96e2598501ad8a8b2680dc4cc675f235c8802e4215d737b6b1cd1a70ac8b974b919d2feb51a1421ce926073725883b2ebd9322d2d6edd4fc1c4c33c0f15bad5f65fa9d664538af3fd17d9f6e77ab1dc4b39eaad719e5dc9bc6bcf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d0726798147d17ad20c85769c7c27a70c61d842dff3d00e8c97801c5d728b5e9aaafef31eae02064a2f9d10dcb82ba6bfec33f1f3e50d354eeffa369f578467ec0134dff419ed3e8f7755a16cc7f341b3cdeb90db502eb1242b5da96698576b0958;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had93f2a0c64267de1442ced90db12a0558f7da9e1ebb1b4b1fc374a69deb1fc6d4edb056ff123e7d0869db6f22a99ae557f148e7bd57a0ef86fddcd7daff32dd6791e9ce9e1ca3cd2729c76d80f8491095f24bc3fbfb5d86e9e0d56c482a8cc3151f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48f0dc7d3ed3691674ec8f3c09e1200cf770ec6617e86db6e42ceb5959d76bf686a67f447e757240430010708a3247ba784c3928e8510f4a8377e9878a3b17074485fd5c1661190bd7e4dcccad903822a57c0e71bff196c2d45643e8849cb97cae44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5ea1e17e00defd9c8e2e1f61d052bcb82217de0bc5d88486f54fb86916616a47b4818122d2304f2cc485e0c33bdaf0c2402cc19eaa10ead65acd79df9036c2aab7d44fa268259a1f54004a33b3ac940f347f69cfeb2870ed5794147db4b4d8419d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2a9b8a3e78bdb3f446ff805affe7aa52518cc0d55db79381cc663718d9fc1ba6c4dace643dce76d3bc243b9c715ecc1c3e62c527001dc2fd5bdeb43284d87c359a1302e3690c1970783604e1c4cb75579f84e479d3d2658f488b4a3a32c04ffba86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h180fa970c2347a1d828a2e8794d2bbb0376f03fb36c8653df031619cc8fc99b8ceb7a4acbaabbe016f7672f776f6323efccb4281d988463642f7d5e9c7242c4195d9886b66d058257b38e167bc9e439a40c1a4c7de2040fc341415b5e0a8a4079a90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3efe4c6802cdc54e1c7d80d1c46b916401121aaed7065db5e666187cb4ebaf95093ccc51a4d7f79106cdf7c6c41198d4332e09fd5a24140321b8192c7592594994814b23814a0a7221785baa4b8985dad55c4b518fd7455702e0adfaa6e796539cd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfb396397a266faaefd6fa1b13319380db88991b65859cd1e18d0ce6f8efcc1bbf24dae125cfe4129d94e0e7659ed526a89fbbeb4058a57e4354c34b311ea3c541881946223d677223f135cead1e1bd06857d18743417e1f11806667e69d5ae2c98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a441aa099b51704204564f49b56254bb6df57805be1603b2aa457793dfc477a1122df481aade01ed09f1dc24712487e29dfa3c2fabd63fb85d0d172bb59ed3bf81b0bc03d7fadf5071326196a392e51426b068eb8fcb861f27f5f4a02d15eddee40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf36fbc4033484cda14f048f2ca9d44e35522e329d830059fcdda5060de923fc40da1848672e05576ac51237eaf6fbaedd044cbc0e43f6ef38fee0da72079536b35d34c46a5cf3da606f899d0df38459bfdcc63a878accd6a6def9fe90e26342c7489;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39168ff1c9588100c365323017188212ced3e60ed5d991e41d7131c08b68ca4799397a492912412dd31ac096ba6d1b45a70cebbbe58a263856f293499ae31e0a85f518221f2dd43ed85d6b8f33c9ba8fab339bdcb16787f420e86aa3353c0b87fbbd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha824891b471e085e4f31f1b9f562dc6d8bc9f7ce8015036d69e6888e1aabf0d4d57168a4c8b84ad55be0a377896945ba62baba5311cdf1c977b808310bd7f6fa766edbf84b0f4abf1bb91655c0ece8a23ec4215c6776a6baf48f618274d37515c207;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71dbd812064a89c8b325f68987460337e2c283c307a9afba595c8afe609e533a301cc85b3c78a420352f21fb2f8fff7dfc767e5901b5f59688d564e31fa729817d28e0868e567f13697fa8b43e6d0f46fc14a77ac4e267b64ffcf8f90738dd70ebf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he24f66e079a498fe8dacf129e2a306555251854c5c64f6094a33aca1fbd7a7116af6d95de7ab31280c52354d0b03bdc61a3a943745a0228c36546a5e145d74c36aa6aae30190bb0b2c0beeeaf87f453fc5790ed53be84a3a37c15cc3fbe6664c6bfe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf1558732145489bc8b0d8637e683e35e5ef366927a7908f12f99eb24767e9f148934ed0c1e770c700ac659ec7ec68cc5001812d71aba46d0d761e984b0be52fba0fcf00e6f45411717526d61d1728f0b9c6910b093c18d468bfbbd9d4a69b5dcf39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92b9b97b839f4d92bcf70edcfba4122d262ccc26600bfa83635f72f30a6a8a715648fa6b3a86147b8f0dc591067e058ab4d306d54b9ee7074ffc4c68e0dc2684331df763ab8d999fde988142248664b5e228fd4ce3b1db5f12876ffa021a55d1752c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c18bcfa81daab01a80e6c1e2797e9ede81c4e038b02069d5030bb211d6826b372e772c2fe338576d559ece7587c6b8f48ff255f23a02f90d7b2fac6240da1bfb312aba1397c93f58006f98e27ddc1c4925d581c5d0bfb987616430e3b4237c07ccd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2198e4e18be2abd459ae6d285867465bd6a40ee042a59cd0b9a8d030e6cf5b79c311fddf0b6988e8c4d16325bc19f8f3e42b5ac685e52b201d1e0f39c52afcb419d4f01818056c0c1dde37197fd10dde592c677d8da0527cba0318eca06a653a3c76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5d1df66070641d0607b24eb4f3328bad3b2630fcb71fdd4d4d2ad77badc0bb16207530ca6c59a99d9f118f4ab54499f7eb89cb63b2c2981e006e2ed94520dd6123935c02034b0da40e88ede9c2c88c89660fc3cc3b5d6ce08c70ae86f679ece7d7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha954d28e4973a4b38d903ef6b2867bdfa054a540d549b3625316637c9eaa5e206f63c0e7e8c2b559937ace82a9de09aff9627161cc4ad2eae1686e55ae4c7aa4e48991760cbec0ac5ec1219f9227db489e8edef121b8400acee147aebd9ada3a0331;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5633ec8bf6ef8a705049ba0df1b7d2377dba28ec3c7bb2342750a4da9e125e69b852de5d1604ee2c891eddf81c1a15389c8ee38d82c721bfc81b3a7110bb5ebda5e0c976db4ba29230cd6352ac52f0878ce7e378a36459b39a41f2af404007bf0b13;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb4524eef31d8f678aeac8c6325dcee643cf81f840e499f8543a1b1ab96bb1094ab36767b884cdda1bd4bd27a60cc0564761847409869846c7f44e156c03d90ae4ed91c624176b1ee454effe212f202657cfe769090377e5b6640f64289881de929;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb3c3ff387cdf42a11c91c5c70e2cd5bba7d574733d2d61505f2e77a7f48442f88db494b294512b1d1f7cb36881a93b8903b3877396e627c527a354446500ce20dade1d26929418c6a5a60455e171cd3cb4265ebd28458d9f45a0b77c2febf411679;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6d6e6da24a119cbc7496a69b734f772f2d3b3c0634b6757afb14e47ddae0cb57414d90f2a8e445d8fbaa3bd545ddeb1164daf84d5f163be877acebb1ae307be5accfe03da7c37b778d5e6dc7552ee84ff6a9cc125a7f295f41038db5cb57b9928e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he12ed72e62ed0fd4c0d748529f1975177f53e267458cb0010c0eed2953e0f9d3ac68418275265aaf2ad588efe117ebcba5229cb21848ca52f49811fec18391b7a61b6e1a7addb3c7e70b477bc819cc9ba692737666ca65efc277235ca4f3dfa4eff8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fd2f902bc9823c33407c77714158e87bbe86d5e6d1daf06ad27cedc2aeb29c2896bf525c4b9af56f59ff0a797864289d792bb154435293efb4d990f1487d0ea636bd844f83db755dd26f1a46c572acb048c4b73e958f806d16ac8c197dfbae6583d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc496ef60b8503475ad57ee545f7e926bc64eda89aed831b424ba608d9855be553eb96dfb89c2bd9b0988ce4f04e30147e1739d40bec15a3ce279dbeca7f0d0f27580eb510ac308e8b94d18546f87553dac93385bbbe7f7733684d0d1f60daaec0f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e3fb642ef2524d2eee791dd97731d16b750aebe24fd1637670df5ff3deb7caa0c9ddde6825ede23acfd59596428972d8420bfa640df1e5ed3c3688e1d0bebddc5577b8c577384738f93ec1b95a5e55bdf3346509fcb70b591ad44121bf20babebe7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6cbe3415b4f944b492df6eee091f475e3b022edfc9b80fb58852b4fad2e805cfff2083b6c26cad8769e39871ec6a18006fe77b6cc4f5bbc24a9199cc5e9c5960acf375000ed58aeffd93802411b72c0697e5d55e06597881f511e903f49a5c8623f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35171463e72a90442eb988ffeb2480cf501779d85dc918cae99848c467fde97c82849639e7d70facad6079abb23d42eabbaf053ff70f39f743c6c4bc8c4fa42e1f2470a158aee2f9cc2bbbcdd20e411aec05f68758c9b7e0873598033a675830690c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60cee2147ea838bd1d1896408b02192738741bd48f78a8dbc6d853cef0549507e3248f47404f86e170fc4e146c9342d2aa208c630be574980394c08578cbc8ff40ec15ac1974f63132e72c5b135d2d7747bde22736724afa83ed111db69b21cc472d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3690ae26c6b33684a25c74b3084e4f68ab47b112fba1a58b1e6d79d84f82cedb67040bbbe0711eae8efdcee2b5ecb1137ea86ad96e043130ec4fd1373196f0366d049128fe4feba69256921483af59094d56b60b59e3aca0e9ad04aba64d313d53d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16d6dda2e0a498d6744321e31c0e545a49e47f1ac6ff3aadf17d3e822be6d0d935bc4f39fc83a0e44344bafe2fe604de6bfba709e80aa32c9bb9be442d7560105b0e20e107872b61203c8d3cc62fbc2e2f2c321f21238e44bb5ea9d1c34cc955903b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h169955046002279691d8de2c6be5936266c1b4a051d9d24ca67137fc1f84ed7277b5c527f763e16d79cb60e6b57cb8d0cc3eb66dbe89e8f1af194e31ad3320678fbbd7794baa71f69d0dbd322d952fb89d424a8a3d4271d7a06c8c78c3aad388809a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75c5eb12dfc06a43618fcbc13e9fcd3057d41219066a0025c45ef6c8205ac32aacedfbbe24415798a820674083998db8764af6d0ec0bb4d21f0e26fd7366d3b75e54e91ef8bc744eb6a8720cee2b430a01b61faefe57508d0e61587bb1109f08b0d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf92f1d164e83570eb703ec56c0216e206ce0703936d8d91de64e201877c0de0a7a9bba1d192740c28880059882ebb1cccd516f898ff014c989c5bcd79221b0a3b7c437e75388f7cf6d31ef4b1ff748c79b3c0e834ed70bf75e8f2b04566452ed23a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4688eb95cb7cccdad8042ad2143a4a084d5956f0af84dc8c2a566c8b95b2ce7fb0edb38bb6497c351d9b367b859429890f930cb93c3a42f561eaa7daad38feea5dce6c7c561bc9b836f8a6f02db14a1664d1536b451a9389d215a6f90cd3572dd3b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c156487977205ac9b1d269870ba6ca36745b989e8c0dc28cae4c7d920575229d04de29f6050e3cb7773ff9d7ed77b7dd20803434b6a3760e14af945b896860633646a9d82ecfedf6078590e55f1fc259636035ecc70ceff1b4ed918c5caffcf581e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha36a70b785849ec240666125390ed2193f9809662286f66e70e299083f7209c7726a6338fccedb263c9bc066e5569cfac818af311591173357407b7720c9cc391f7ab2dc4d6d65ad4431924a3742b4cb7953c2e7f8851b0d6d7072f69ffa85963a05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dc229718e3b257f56b76aa288406903ff28738dc7773b1ee9eec28d135ef605f50b2438cae25a715bc0241e3636a0fedba41ef8609b9cbfa0d87b53b8f0e0b5d6a6d81be1f2284f9bd991c5233b8277fc296e00ddd322428008b5442b1c06ed0c5b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc754e8e1b05109a171bd64335b0308ff0ba642ab0c47e774ca51df870cc9dd710eb03e255eceba9174ffcf3ee3da9efafdda9f2ea7c234c8d160b4749e6aa970a3c5ea18630778ce02f147b498818d101057f81f87002d3f56c3d3ef7f7a0eca5b5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haec9f5a623b15f1e69d56b0effc8e47e2f07a22e3948744d1519f85aa3de2054956504b1281a22e6bf422fa4bf07e60aa61ab33e483300c7d9c3f32cdaaca64b2c14fd00ef9cc8a5b4d7564dffe430520f60b7d46bc04296ba993034b284b22a4816;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ad12c303aa095006ff5e09dfdcee901e3cc530d98f55f314b5dcb303d8b91c34a657e1a11e0ede3232aebb411b4f39a57ffe9596c2834aa0b87a0f2ea45c5fa232183eecb6fec5a907502c54d3e453bf6af4d00059c782d5baacc52262fbe8de8fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c202636919e23a3842ab2d8e3993bfb2add591af4ccb5f15777218150b4fb5b08579a744dccfe14230f833967d7c3bd32fc717bfa98203020240301f547b787dfa4a2567dda574b5b64cdd2a7b57d1fc7c425344e0abd9c9d415dff9a8b4fd8c21b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aa30242b68dbff18577670cc3bf88efaacc3c07c2730f620715c91862296eb18f83cc11857420a6c19e011f9a85e208d33dff43a36a9cd14c8e9e0f1af29f80f95b0a654a73c952deff613050e679872462752a15fbb24cc623b75d55d2732bb9a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b67508ceafe3831d6cbaf1e0986573410c1fd7ec829377f53aaaa136e8dc30e859ac06d27488464d9521d1a476d9a50d005e0217642928e42b74ba23262b79f6bcdd20577daaea8448b0d8f38eb937797fc39ad34ff7f2a2eec3aedddf27b63848b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe4705cade0d2fc548ec90ee6b4c253808cb1494ea1dc4b1a79231528441bfedba05c1e1af2feaf09e9af53e75ac58c5f56edabd741f3aa6a53ffb688ecf3a4eaf17a2b27e3217f3f9a9a5b76ab357dfefcf9ce1e891dbbeaffe77ee6dfee315bbd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b27a9e89cb15ee8b141274b8d24c3070232310612b850f598b178922ab4b743addf5730e3eaade97d00f9a03b303d4fb71be8c32070020580743ab198075f9823d75b65303400d4c117d4408a7ae91fcd41655eab19857a1f6b0a4b5635d0f2d269;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76e737d25771d1ab189aedf64ef3f7f883f88f7099283ea269bef277bdca2380452cacf16763cde9458e07a4dc74294a0c84765e0428dbdba404c96d1ed3b1b8351099298131ad387e063f6be4ae2b5507b803e289097df2b6d8e479554ddf1b9dea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f9e24127ba76e581321ce3095274efb0ba08147507230daac293cacc89eee424c6e8e07f67b167f6fc3cf8d0fa90f44a125c5780ab350116c3d4582f855d807042f28bbabac4cf3fe6e94a75bd00c351d4f597cb8fe2b8e02c0ad9d0b965f2d8d86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha97a30808337a3aa218435d6de6c7b6c1e01e7759fd2b64e54f1b46e7067e630a654a47e24516027c9a9f028291f2d75ca8676244e3de04e22c49a972e5176fc464dbcb06f90855989060c0903baad1b9c5a60b4eb6c7895bf37a51fb37076e55442;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2fc413d74817b06791dd753fa1b47c889fe0e4ebf070e1adcf74b4ea0e4ba9e3ec6ece7b2af52619fd85f4e709729522e0aefcf4501c82c1793962bec97e687f9a5282b21692be631f8aaac755755f7e640c46cd5a6e76eb00b4ae688eafcd226ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bbf5e2821228a7f46d6a1db1eb2b4184d20e5dd586916924527d25980cfe05276a8417615d8095b8aa1360f1be9c30329d8701c12af9b5e66d4acddb8d7d5ce8ef87d0f84529ba9d1604ff7187a4b70c741bc2db35304b94f7b9324d483ad6ae527;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc94cb75a1c5e2723bff1dece29d84f8288a52e293069b10bec48b98f7cee5dd01ec18b6f892550bb55fbbe0ffdc670e416625ba15b8cf4f3758e5e47d31c62cc47ede2b68ea5527d251d040d4d7104ba50b214688e4edd1636d94f8d5007f9fe1446;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h101de519af02f621ba41875986cb924417276db8b3b7f40039838f5c2b6e242d85c848c3292b316814ab5d1f855502b9202e4e7cdf309572dc87953dfa3972784b6b5fd190df449c48cb3ea86e0ca7e0644d0d15003e1b5ce54228a79ebfa6998346;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bf27531367c523ad2d0ed81b28727662acb5e192e2164ebd131f972cd449893ca3485b8a820d786cb232ebd8d7c4a23de29f4d5bc91d5e7fef43f4408c5267108b05ae7cb8eb8c4455fb659938d359ae5fc4a8de3df83bc0dcf78394dfd258f111f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12b15c020ac86c3b293498f3256e68234ea735acc0c2d710f0449d808f7ec54f7d3b54e717dea5353aa33d847e5616a3aeed51f6c90375e063bdbfe7ebb8d9519da00912ccc2149fe78ea0f9c1fa99ef7eaf7e2e9474ac2878b8b83ad85fd09a007b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0aa5a813c00a2356c7f2308a83c5849d19c2fc6fc98c84e3ccf37dee03d38b6656a67ca2f8373a16b0d3d27d9eb24d8f223fffccea98ecb9b1d3b3d6b0897de4214c5bd7ec77cbf0a84a9d0668a2e54467a5f790b0804d8b7b67d85f0541a449025;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e9afde7820b5a2cb563b760e21f1783145d5d044f704ba61da3b3866109aae99d2aea7040fbf1ff417f8115ffff97a885f034f4046a04eac303751021585b57608425ee50a3889372cd1b1b07915a57a102ea30b74a31165da3f494f49b83ee3628;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he90cb55bb0daca734399c59c756c55474dcb77b6e2e7d098be57dba6085bd466bb2340a48a896e866ed9b261fd35931488ea74b9cfc8d57de117703023ba63f6b0d037eba41164f5afbafee373a0fbe578b92b2279592f1285b75e7b72f32797b35c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hada57b977d647d15fa91169bb0e36a49d56bb7bd92d13a907be15d4dace5c3d7da484f4fb8381951c5d57a09fa5f0c7d64e983035399f410e6f0d8c856b08801ad1a6f404a3286291584498580a8b5dd50d0a1206613713a7e8e0333ecbb127e5b1f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14e748d79d8bed38c6633d2d60a481e7e034d77bb255c098fd670528d484fefa14d9ac9e0d36b512babbed6498d484fc563e9dc711fffc77ec870b3cddf5a31041631d291ba6115e7820e33ee032af9dd651ae0ebe3384c07accdcc4c7a1f833274c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf93eed9fd2e98812675a6ebccd63226a7d87d3cbb7e920b4745b9ae7fa27610cfeeb7ab880e04a8bf52a04fb016a3abf73961efd8da630a7c88ad83a7e2bc479ed048c68563399de3f2bce2a40784fbebda2c2aac170dab8c5009a6c200cb70be63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeca909f695f64eba56f6d4495fe0ed37f6a2115e86632656fab82241bb318c1b07e434ada9548b933a7905b147b7ab8657400d33b5a8eb6c0cdafdf3ea3b02f885916eb8ea9d11fd977b132071f34bdcdc6b049b61020b11d44d4322b03e046894c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8b02eaea3da49d004aa4431621c907c84cd37e1df7e572d338e036db7fde0754d4ac8daf04a7a0eaa32465484287ee470466c9f586147cbfcc62b0cb7f6d5c56164029a209a8106dcc7d0fbc111c488a5a7b6b1d3204062904aeb377e2028b9fda6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83e3efc01434744d47d83128e7c4137cf0a0dc8ee878c4e2410ac9e9f494b328cdc452c7518c3bd9c4b78cfe1debf7f81b447692ffcaad5c0b916d8effa049aac79cbe0dcfcf1c46fffda6d26c8d3591ec55b65feb80ed7fbb2b0ecc51e4c7cf7225;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf64a34617e4d1aff88d50a43b368309f4792790970b2f0962457c7ca8b8293424ed3980f67824ec6d09717be01c91d36b926373ecddcb3000e9641d515700ecfb8b7165460e5f6888e4dfa41663cc3eff0a91e30570e3ebe394b94de9ad618065be6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59e2fb1d37be675990f2b2d21c07735613aceac58460fa05d1a8044b2967a491d55c3a9e56e98bc276829680f06362fa9efa18ff9807703238dfe3539a156e2948fb4c855e3c459b2e1803693f70fe60282a132b525d04b253d791bbd78c8b48cf5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bdbbd35e60edb3704d41bb83cef3075fc8b38b583d97e9eddb2db0f69e1e6d11abc54db2d470c7b7b2c62fb0fd49f2cd49306bcd972d5dcf42ce486dda52b78cfc33d4443700b2b61d0a8d11b63eddc7be9599884730681db675bd0c3fd291d53e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3371e5e60e1e8824e23f0f09263ad71c5f371e385c8ab2b34df5825f0be51584334b7539f8875824b7a9244d366422ea1b57f6ea20fbcb7420a38a5b33f469d99002c06cf9fb34216f09fad2c54453f65b800132ff4b931d34a9249e1bed39aeb504;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha886b8919b897173d148751cf18e9307c00e652995192b2ea556e08b79fb7c405e5ae1df62a5225e0934fdd22edde365e40fa619afdec87fdd964ce6d26b7359e26536519b7f2fc844c80dfede58f34fba038f11bc07a2773e3889b2cd352035a3f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32a5fe5fe003c39c62bcfabe71fe1915bbcf95207396abab6d2e72b803b6de1cfd5eaaee9a6a9e8e59f91e9a14abf6156d9f5b42533f5f7a8ad4821f753f90940ba175653232a6916852d8eb30dc8eefeac7eb71101aabd5306820224fc6a3356daf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3a9cde402837fb710cc4396e2077221c94b1a7d62c3ee83c9ce223166b1931d4a15b7b9f4aaaf1561a7a7f813227498ca4284aa0061800ebedef95ec8b1c5d4df2222a6cfaa6db8f3aa493f372c707e106a194f772dd29cfe5299e697cd7b6aa515;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf712d5a9ab174344cb7343415bcf17e4ca4768d0251203e5605beeeaca7989a2c3e809b56b60051dac2477c2e513b49a54dab6edd4e237cd9d2029a9a1d88d954efa0ee5385ff47be62728095fa12c397b6819ab1425c15c9292ae779b8e9f0058fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2cdedf1ccc31d6306198df69d089043753c2dbb43849f5f3089dc96a9cdbe9192b78cb1fb19298933e00982869876d1e6e4ccc34e896f19fbb20b941cfe64454dadece16c3b5077dde69d46c38e3717b5c2c778a0b2a16449348c0973ecfa1d60f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h398027b75a5ec56f02dbbc8f09d745002ce4f1df39c3de3148a8683b20f44cd3777204ab8a00f92a50ee32174f23af59bc56f6cae792a574df2c5a1c0519f4a7fff9395f85986ef9eab064fc3b2bcdd9d14cf616f18e6fadc48f437aa56207b25ee9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbc34c3446ddd570d0dcfa48f9484162fd6843f020efb30863f73cd9ad130735337ad8e7b2e98e7b6d1788ee338c026f73b848b983bd18deecc3173cfd359e8efa33a3b7692719be76b808e6d3b8b9c99bc13b269cc6c24c28f0b2d137df42a60c80;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21c89b30616d78c6672eae99013f0e38794b16b1a0f11739b1a5082163f6b9c306577e635259f05bd4d31547da4cc68c3c4ed37a1df7200ed9409091d88ed1173c481c34e6aa98d4460821d350a159e3331c7c719b4300f6d1fe07ccf6ddfabaaec5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3e2733961d332229bb6daee591c93d986f2a280b6851283a91cbfb7f8c57b5f4cdab601cd2f0aa820f8d39f726a017c8de810cfba876a99d89b8daa259d7b667b4028bf0e711379bde84ababa3bf34949fb88974a26ea76b59e1e46e8022248e626;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c4285153d6aa3cc5991559521a895863b53972b0ce6f2f3ff6bb051a01c3b9bda8f56dee37ea54e49c6c4990ee1234fb1c9c431c27129f5bf924c66e2a75dc6ded4fbd1f12a6267778b1c2ad1d53f1ae349bf1275d2623890fefaa0c4558fa08a92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6c8c9bae7462964d537085c199ef4f0edb50006d33428f700b930a4f71cbc997f2ea821803b3cfb35a33e813923afee9f4dc04640af3c7824ea1d417f2ae7c84c5c24722b58143ecf2c3969262823a936aee2c080b038c2c6d488a048045a41965a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82fd41338a7d3f2307a03e0e8c5b94294839fc4b3784b797e30c1cd33de5056c944912a37d193d3e4c9dea01f8f36c82221ed032d4e8f11cc4222d11b43e968be7975d9511ba21a281469a781e31e13be51b0a500b1c669c424da6aa1ee3bf9452d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f4687159c1882a38798be380d71e56a4551358434dace0cb05f861e382d4d998355b66200a308406558a706cccc633d7a930e01b7f42438461355b14414162bfe1200fb85b290f39bc555ada942a7382b3cc13107863d7e1c4774cbc38af24baf6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a941fdcbe65137abd61eb5194b040d0cdefa8a8aa167b2aaf5e19a06dae3a88e896aef9c768b4c63a38da49528f787f6b4cfecf5699140b27af4b9a9d4be827f9f038cd0b637dc90a644d73112c253d7c6096b863eb8a3b10f2e4ff6e28d0827463;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb079d93d5a6af007aa4aa3aada478d5cbc65efa11262d6f37a4df11803a45b0ef6af8f68243cf4d8ba180b63b00eff6741456b382b050f21ad4ea24b4c4ab4af3902c9035149fe67194ecf7992c4d6b3831ee872d0fcdbe17e91dd7f33e2fbfe1ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf224669da85f7166912fa34ed700706b6aa2041ab1ad5b9a6eaba987737611087e2b0817143c02114ef21a0f2ba2c8a975d8b711825631b8d1c28ddd64b8c50035e4cd991fe0f2e3fc38bb1ac5475271a2f3d2c6eeed706236e9215804f403382215;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h432eeb8190568a00a2b3c589b3624253ed93fdfd1af6669673eac8e41d4b5ee7c339adfe5028bb5ee86117778a16af68deeee2c402e014dfc572d8e58f6dd4fe20471384d7ba2e768a3b5836437e59a449a8261586f1ea36a84ef0b4edeecbe8aef0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4425d72d286fb35ddb40225beed44330650a736fd32e772188f52907fe7fe379302a3b92041fecdac15ead661cfae43a184d4feb2cfdfc73a060d48f6859d5e26d49c6ffd8665a8dc194d209b599f72d900dbd56db138624f9c92dca2ba9179b53dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ce4ef70079e32eb09ad02f15b14f0b23cf10682299c178412a7994523a1659a6a556dd924fed9e348268a48eaf9d4b4bccc1f1dcd10f6842dd7f5547fca740cca7fa07c5ac9f52deae7209173b80a8b1050e434030428f50fb2973e6a77d80be41c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42faafb610e50a546327d9013ddde99a99321dc07bdb738fc04f1355d4ca5e4d4a401c149b4a6080f9e89d20b80a858ca4cad49f2ad8c6d8231e2ed582ecd9bebe4ac7ab736788fc5dd8551c562ec5192e91ed8b91bcdab535be025e9ebe86f67dd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf06ed644516ed94fdfea9867018c31c9f11ac697164b11e11ef6e2b51243211ab5a958d26a892d34d9c66a4873ee655bb2d4515682133aed223b3bd5d77517d3e871aa9471007b208a946e606c75eaea27d75f0ad85c2fafd489aae5455832c2e1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97a0dca8685e1812a5367e6ee1dc5c6a7b4a9d607639b3b5fd26798d03668e805ec8bc1c0358124679e3f69dfe6195cfe09fb39b37b4f20722e26de3ef30f288a413c40e7acb6434e509ba8f36789aed2563f6f9683edd44798fe593bc2b19cb4582;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7023699218d662192e99059d0700cecc3044f6298d60b30c374f7f39841f13cc666407cd322c381d3ad97272263d469398c804c8703e59938b71f7e1acf6be720054a18bde5ca47a7964f7a1174e893818a84bf2a47d1f5a96ac8c50a33d6e508e0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf040a889d61e41c1ccf242468d2a536d889889e6c39971b676f9a2155c32476308db004adf3792e7b069eec7a0ee71b403669aba95f6b869da1cf1c915cd3bf9258b8be7c34b95f3a3d3f01afeced55755e622a3b15a56b690e0d07500b92118fc54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h545d8e77ab7c141e046bacbfc0f0597d291a2001b28416f6db32f48f7d59696727fb7bd1f96c0b9e52de73c0250325c4ae3416f214a4c3280eeab0447b7af9f1569d60441a59d95bb6a72a60bba5466487143d0d56907975809410c57bdf367df98d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdaed8247ede10f29b63e47bfa818399eb8a089d5827bdab9c7795146897888492d795a54b8de82290c6feb2579fbeba0b97e18e37e509908c15409c2f18a919bd2f4fe7390bd9235afc65ef2b811e992faa2ccb86bd6f9eda4db1e39350fde2642;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda99a046f44cfeb3859fcbd9c3897a927ab9cd229bcfea9be79794425631055eaf873168072936d01d3ab8d1a8474a25ec9559f77d63af59fba9ecd4fd19bbf64d213aee66eaf7b4e1946ec8f50e43281892cb776d03f0d9ec47e65b609178f99942;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29e381b9d89eec3e430cfb70c3941a271daf52e86b187ec265c3ae83d3c905b716028885ca48f6808961712eecac4fa92755d4017869b3b0782dc11b5f7a09a76efb0c3bb7a0a90076d205727eff51cc83483db2ce8049e8de541d9511b8fb1e2601;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2efd4b1705a83d159d64d6097a2b076a9f0bc42a79c8be2630c76ca265a9c8867cb239692800143eea89be09ff251e0326494eaf6dfeb084fbc5564115ad74842239d4898962c767fe72b98214686d1d55d27a28820a4b4df37f9c7f483d0a39421;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d074794bb72d8de4f26b9ac733d4a92a769ddc541e35009b78a7cf1421e2da429c7b9bee003e1d0f302a94af7be77f746e97588cc51d3abe92380fd097d59c5043ec366a690558456fd2fecf2845bc9db2926220762ffb06c9d8160e39d9ced3395;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h127c45bf4dd969a3eb1376e1b8a45fb0dda6a73236b66b096bc5ecd1aa2a4ea332ad299d469a53859ccb00dd1c27c37215bc125f76ef27f49f2f1b4875c1f665222a7abda986527a46f9dfdb710674feb0d8e24749ab4d34de2ef2e519ac2ed0550e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17fc4b543ee3d4dfb3a585cfe9c1620383d7a1f3a54a5497aaccf30edb419f51dfdc1731008277839524cf1a0eb6cde8ca78b78df195bfc2207ee416869589dfbbceb837babbae0e767bb16785b79043209073cf325be0917a12bb7ebc5cde18e81e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8cf5c8e655424ec9076e108bef1ee3520cf581255e2eba948e3234dae11429c4ae6682f66a62034d295e5a0af3a87299dfa86592e7a1edd42aefcd7e5d80585d94ad28a3653993b9ba183542d47d3ee74babbcab5634a769b7395b93dd53b12fd0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b0bc0301d6faebed7dbe49a6658c053c79dc95ad631029811ffdbbc98b69cbbe95fd520b08312dfafe7b371f50e4cf9048a9fd480e1ef4cb23032907bcb599da5f4ec7a26a636d87dc109e98346a5032a47499b53cffab8cb7b7657f2d57c59c6d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45dccb9bf43f9d083c44559e3a186f0f472ef7819da2b72b4f0b452edbdeb2c97a6f873577059825b3e8cfb3c3e640fd0778bff46ed4612ef44c15dcb6d39dafe460e0462cdc940444b9ee07efad320250d101f1876a31e9599fc27a90ed652add0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5ffaab906842b46dc11b998c98c6bc7007019d1f8d0bc3f87783b4677903f38eb227ad04e452976ceff8d43484e9710c9b06bd37cf78518760a2b5f11319f04de6c2dd511cb31e213322f7f8c7a684236879246bd57f93f4406736d55abcf425833;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68748e5e23d0738482d4060aa06f3beb46c3d2ae2a5e290a83be37f46ad6ed64ed65c368243c9419b7436a68416e07a813820f04e5625077171e6ba0a7641b979ef1ace395d19ceb0b661908e72e69621b848db073598b22091f35bbf10b81824859;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda410a4f762d28462acf9130cf089aeba7cd7fbcd803405db89e53cad220b60625afdc85ab35ced5dc7e1e0a17c46715b3a190f06efd60e240be04c653d4627d98022493cf31868d203288bd425e4e3fb1d3129069535d22018282f43c3f6b1fd616;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h570ab14dc9007bfa34f987b7d54eec0a700f72fa4ce69a911ef5eedb12500134b05adf4154f8e00ac6c20143d821bda09ff1683d2aa501802684f9c937a2cbb0869ec431f057078e53181cf4173f7e3ae1546d4b1dea19bfaae0fbeafa9e7788efa5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbebe698c7f53f1a3aeedd6c307a954da913516f11efe79df0d34679a66a504fb4fb854e6b9a679bb9583372e0fc0ec5d49586b3df32dba5601d85355ddc72d118697ad4971d148f96930775e91f4d0deed2a75734b8ce8f5ae639474cc1e72136a5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6083bc050c3de98092af28304bd36b2c46036c23305ebc298350248cd0c13b3cc8d16936d9bfc9673183d27a08f2327a03374e0344c3955ff44726479c4aacc0f8691131c76451f5b410b71f4ad12e957a0abb48dbec0515cf3859185400339d805;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77c1651914c3927d25cb160dae1e54a108baff906307948cd6aed39a8037a9a21c93d9d1bec93ef9d1436f598be63d9b532a5289ab875a4a6bbcffd92c6687ecc466786fa2544f9d0768bdb20f41fcb381ea197021499add71a925b8f007f5e68238;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54f1dd3f7fdce349ed3069b122bbecef67a3b82e9624be2be95b38a822317781afd1b94a8ea960698a4a0d883dd1ca5a7425f7547335ab1f691daae809544654773b735f5e67ab383a6387b0b7b059fd06482a026bd2c3f8cb5210e984b6463b78b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81149d0a071ef246638893ecee0b6c0de0ef815a108c67345f23ac910a812ff8cc1e25d0e89e15116a6b2e06803ceb4a5cd3a9e1bcc39934accff8c94f0e6793a42610ae7c3ec3762d1502924b4ce83cfc2f0d375d4e546c73a1d7defd6092689c41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d3d47bca93e065a0b2b507f5b1cef7b6445b5b86b0ab52afd0402e260e23d4c3c23d11fbfb7f69c1073407910d35a0dc7e992c1ffdb1b739a118ead29cf4144573f6247be1f1b5d42ec2e17a4b81f4975eb37536e4ec2b443fdf3e2dc34f943152e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7b1a1bb90c5999dea55d7596093bc6299bd4c64e0f1c09d657b5fc2cf6df85009110e71bab9424e94b73dfe936f8240b32073606e678c9a61a6aa99dbfe320474500160956416f69a3d15c0bb46a85df68f1fc182068182b96670d64ad761beb774;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2d284a33e6920a46a63a249c2a20f6bd587e4a66cae15b537bcdb58fa0c373c7a022286bb775bd3378f7bc12c896121f88cb787987dfb2acebee82f40b67a2ddeba15780a3b63e35a25f2876253043ab7ff3a6fdb379966f417be19665e4c8452d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb0e3f19f36ae3a5dfd136ba68d6846c3617d6a88a46ed55a4f3de0f4480caf3eeac78699ad783f2be18898037a7769078fcb500abe97f5a06937ae6e781cdae245c72c62606116653623108a1d139a1eb3138ec2ed1bf05090a8378247436220bf2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1c6d3266e06ed6dd1f6b7431c27fe5e52aedad4afd0ba917e6d2bc5a58dae4eea3fdce426b4e28a0c45233f29f05e3b8f30bf78ccc8c4a6bc4c4acb23fb1c4dd03395bf0ad1763f44939b1764151493a1babdbd8b6bdd3b20aa0afdb358613e434;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb771adb1db56690182945e8e6b7f74f1d20e5ba8cbff53c120e7c60012c1bc5a0dcc8c304bd787e9910adff2311f90478e7b1eb8dd11079fc28396b513bacd1b55009ad85a842b0314be3b080d9d73a1a798d82f03a39bd87b4b96a0d51c0c89accd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19a5d1d00ae33d0e1ca31697258bddc3d3aa3f4b910f9cd86f787b7afbf9141de852b3937cfcf01ca64f1524e7c78d9423c748ac6b174efdae6af109d67b8a8b966ec357837c96cee41e16876ec0b1c102c276ea135004ebedfdf71cf26f44e84254;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ec7e3bf77db6dc2e5749272919c8fb7908b2873e572147c5b5b5027a40507353ca0474c33f64b131e2df7be69a0a798c63fa875171dd7e1f0c225f882018449962d5b0abba7cd06f9a1286dca2649a533b370059296955e3c9f0b54180f735a9a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23dc8e319456f428965da6ad5d132d9b80effbdbdc304be94e163e9f5e524d446fa1be5a10176a17b8fe2a5f8cd3bc81b9a19cb779ee0ee9e1885070f8334bab86ba565f4d6d9552a57cfd0bd448cd4505828f448d3b273da76fbe537a4b531898bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedb3fc34aba7a391fe156ce0d9ae4734e150b19727023401b9422a30344db2b211d0c543bb12507fc3c3ff8114a75e5198372c7070f74056d95f993ce1f4c3eddc4375585e2357dbc1f0334268417036b4ebbdb889b44f5e90603bfd709e3df792ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h825b7092e933488bddd8473b6d5c5a3f5ba747bfec020e210baf9947d452e4345f9d50487c85cce61ffd191a874f28c8ccb81ad3bf35fd8d8ab5c31a912f61337017ed9cf5f075789de349ea5aa0ab3d08b8cca1af2f55c0ffae705275636842b1e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9339d9ca2669d2c6fd638741d7bf7ab3e43e17d734f22b25ff66f84f683a8ff1fd413b43e0f9422b27dac8d6cba9e20489216c966356264446b17aa6587ba9a1f90a6f8058d2c7f16838a3a03a2a611b1acc4718e7868225829f8661c67e9dd79514;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1f1fc6c82e73d245a6403673d4ac903a3a3b57e2d9b0d51391a6093942a26004018a0e75c48f51c11c3df5b265b090c065fbc07afd4dc5b710a5c79271d6b8104b60428314d0944201aeff0dc95ae8dd5732852b0efeb744f9b2aeefa285fd5fbe4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32e94b7cb0f1cc9c0ea4537320e01c52c3c2d52c714a267015c1ece9ca34d57a346b2518417fc127febae09cf6dd977aed09abdc622ae71c86f31b14dc377056a7cf23c97a196e404b87408734b458b8003882bce0a06a6a3ca90b9bed1a5ff17a55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91e8c75e7a8ed9032cbf5d0516f2a8323b7d48276fb8f34fe2648180af5704c35e03a87466f3f5b93730c0cf16f8236fce1fba2707d5592149916a9249e164684c8b5eb8bde20280b296cf0c453339398f4fa7b794ed6924fb1d21e6f71cf8e7f194;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10828941bd93bbe864f76ab38251e9df9ddc7bcad9a4556951467374b4572f61dd66f4bcd331b2c7ed926e42641183dbb6c7ed77daa7e8c6bc65d9fe9164a2b1698fa74c3807e5ce97d55f2a526814c075c294a5c0d3221e24a9e6a5b3a29e70085a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c2f9c0d0bfca25acc7790fd2265808bb996f31a02f99914c6d6dc543ebbdfd9c3d9672d81b785b728b24e2ea5e4a0273f651805b36090cd4883c5c7477435dcc04a6d19c63f3861bb45f28a5cff0aae592f07d5ebd8b6ac1628c4bdb1059cb78c9e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21be8e06984962e2353b53786d2f902e41a6926bc975d6d0dc9a19312fc7d190b02cc88d975901ae1ed75409e10741370a9e628faebabf654e3db82c9f086eb6be1a28fa36791073f43af53b87aa896b15be503ab7333d3b62a90e48b81a8f5ed2ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49dbcd9b35db57c8a9107190c86555a14079e24ce55bee81628c3cb04f4e488fd2f36e86747419ca2eb0989b19e1b8a93f9f306aef1ce90b7b3c43c194305d82733f2f29f67144b1ae0ea9f7bb00eca15ae5332e7bc355060d3223fcabd4f58e90b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4160dec98d286ddf42a24104dafefc81a132dc23dfe106b42c55281f701b59548e042ffddc21899645ad239f8b03d892539eceec4359ad6cf9c83d7a25c8ac33241fc54945f9c1e98106e68cf20eed6556e7af3f86aa3bd98d62d8eb69648b878653;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb133fb5caf13e8990a392b1f7a0d0ab5b189d741d99104e6aa89c6ac23c62aaf0129d6e79051029a0060123c30d47e740727836d63a3aed3e586c50e45a22c179186b5e047c7d4af4acc0404b801b7953f019b2f4f81f4b87f1bdec7968c0d34ea8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fdb41a7896cc63f115fbb95d0d0058e01ec3f1f290fe9b04f7a147ff957ede09c9a2d1cded3020e480bb8dab4e7dcb1b5a90ec952ad5071fd29f63c0011b1cd253ff9c1300824b00277c62bd33b559111bd5245a744949d8cf43d1d76aa63cef06c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d0cb066d6d8ede7cfcd215c90e12dcf612287658d7de6c04792d1a78edb6aa36db19d2f1c783ada346a2a97d33321167514e172fa93a2a4ecf1ec0b663bb04c32b8f019ae6e9852421d9d4f866f72a20e2787eb8a5e4b519d9c3345c8131d1ba3a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37cc1ba7e00c065ffe2442542a91fc2582a562863045d9358ddc37e0b2b9c12d7da2101ab0373e83bb49415d1cddb941391cf72b385870134383b5b5a6867432a18e2bab444459b491a97e12b549aa8cd4a1712cbc83ee90609f87e762f3d1903490;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he047332dfba5327db56c117f29f35c51b53a10328d2316af0b5ead36521052833d1d18cee5cff5c29058c082040aba783c2324be5e6fd45cb11725368194025abae4b6e046214ed51a806834598b928e59f33c37f98ae77ce1bbef0649ed2168f5e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72aeb3ec294a12a04b8cf167a384655b6b8bb71952d1bc72c00ce1188454d72d5c42e90eb91793898514e049e3206e1a2fd20273690071061dd7a5a4555a03cadce8dfdaf3b1505f704679afe2c4d452c08a3c363345003cf34cd42fb0818cb62ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h395bb04c5bd8f41824eb1deea623c7ba8d7f4720b5addfb0265aa5f896be2594f665cef3e97a2b219ccd345247acd7acfb1dcb47ee67d76bc70311940e62e35768f24bd2ff0aa3d6efccbafc4f558d9bc7d82710d6e2f15c19e6c500b73d2bd21703;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h387d6ae99204dc46c273eef5baf06bff38816a539129d57128e76caae36c853c92ae11ae741e400605b96b3753f15555253661c5f21e2d10cecd4b420483af41bb0a4f756d05c11dc23c9d54120ee1d9d1f7db2c4969a31e7818e76b41fd3281b64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6c0c2a2f5433a4db0511e5cb6049842264dc8c827d629e1866946b1e29e98502e5322f317c949b2b1c4ee3d1ab9171af944fa23e489d440336e76edc6bffe0db21000a5ec9aa4e81ac4ca1bd528d8cb7d4ae691a312f985de2c58f30e8ab84c30bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce2b01611835530e7ff427d4208e075abb4575e07d40e262181534444be01713c608979d4155745651694000221861215e2c2529275aa5babed8e4d818d657ac5becf7629ee199a1eedcffa96e14a5a52b30e3159bb6304885005c72d18341530a17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he015f92cedb3f5c962603023792bfa4efe6234454ece34d1ba091dfd1da9b97e39929ffe06e3e701fb409f149f14ff6a5fbb8fb4e636f7f0a9cf2c2f96a9611bba9db4cda0d6105ed3975f29601fb05ff8ef5bf83e75f76e5672f2290e8fd75b6744;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd73af344cd713ac6a6ace4d6c3a6e09a96e98f5ddef3144e5bc9ffa9d7f32cf7e9b1439ce241732101e90b61da1910c0f28f8eed9e025fc5956058778c5a8b09aaea5396ef4d4ec52998edba76b4d859bc49d35f628d8a2e73be16a613cd5dae4e9c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8db5dac4702bf369a93ef2137eeb6f35b135c947c81be1a6a0e51b86b7d3482b7627ef230ed24b2f254640eab9541f30cb52c59a5b4889632061e3a18427553717c5fc21cc9ccc0c3afc124128440b9b8b067744670283efddf96884d79cc99fb00;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32da2578c54793048cee2c423713c1d307a540e671bf1e6fe7e609295c5132736276d2071d2ff39cd90d16852e62b8fb75e36428d8b292accbe3e9ecf6f6168f24fa0af0bc1dbfe8264148b7de4654481a993421a7982ea056a9755650087f823e66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h401ec15fc17b9564352002b224853b1acdd23c0a191b9fe62194c6811c649f63ae4dbaa8c9a251a68b34f30781e97498f69948b5ec62e5fc07e6d0a41f30102827e12de4e9d8cd2c7ed194138921bbc433b4a8ddb2a4005e81a7b9fadc173dcdc39e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbc948e6992521b504874edf116ded63a0d2081b170023818c26047b36e9df228c46108720ce68c76ac0c2fff545bed12402b07991978a0c92cbd889519a6fa66015c89fdb64bb952675b55e484b582e47e249ab38c7eae6d5a3104b7e4e43cce2f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h782d44e11ea512a32e4b4aac991fe5966a0176005f997572c46075ff19a3599fbf4c84d0f05ecbc842d29a06442858653b65b0af932a8bb10c5a3f0682609a85145097b0a1fb358b7c2825172d0285fc9bd5204bd420c821b9466b576f6822dd8fba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90313b58ae740b189493c20f13ee61c0bffb57db58ec6d97925d4d9b1ba238509b7b51d4c215925c9ea2801f6fa9249ca572b370e021852e9d61ca7132b1ad99d6928af724370c3fb08a807ca4b05cb7e812a045ff73b57a56f188a7e64b58f5af16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d6034608db7c80b864a354b29048d0e851c0f1f0375a0f230c4b1da61a408799d3c7d359ef9780cdba2f64e700ce3f0ffff89ba631ba3bd83b437ec84a1c58121a3987df04e2175e8f57e573146899a3b7b1031db6ae3c088fa446a84d63a838a6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ea8639b90957734074636089857d95b5a1060fc4fb8f94ab25d140ba5de857ea56620fb8dd47e4e443389dbd27aafba4d1a9f01a05087443d70651c247c53df020829c700ef54af63a80f1d7de299352bae3c1d3184ec48d5fa5f9ed3df52010de4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9d2ff3e0a3716ac4f1c0e1cd9d387254fde912c40085aa732aa70c439a29d72270d02e0e9b25be5a61eab3394ed38cb6d12ec71adb3593468e81a92e3563c5ed638d994fa7b7c9ab38d8be1c4363fcf9f3c7b144ba0d2aa6b87ff6f87d7cd73334b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cbddbfd5c3e9aaabf401f5c8be4d5c3dd36657db7f3deaa3fb0ec904ea6aa959d7a7d1150e87716eda08bfe7b9325b9bef830eca70ebee3a3c737c7ee2656c1f64008e2479fc0b9ac140fa3611cee6c9b0bac79fefc6dd0fc6dfc3b0945dd73045;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46b825e5aafabce752ffa7cac4a1cd7133414855ef6bd56dfb6f50dee9a9cbc6d7e7ca3170d1cd2e5fc1264de060cd550ed534dc940436393d0968771ea6917b9df425b8d8750f35b23a3d3017dd4171c37af7a3f7f223038ea7c207f52c3799b0c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60123d2cbb15fc26c3d2e7eeeab7518d631c38722b778d2f17da695f3a51a84efec1006fada5b417ca6485f6d3f91c404143fd6ebb6e2b39dcb85297f17dacee523fcedfe8bfd5969a177c0d0427a1add2e70a2bffd9078d647cd546c2e93071712c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0108dddbb32e0997a1a9f1d09d2c0fb321157ab5a25b4697aef2f56d1edfc134d9e522432d946942f7d349b2a997bd03ca99f4d8472227563ba29a34c0d910be3fe2518385ee31bca393ab6d992b9d83e8dd4cd8fdae842125da44fa03998b8162a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c3452b686f7c5e308f0c3ff3c6a838c62ab083b929d9d252a622b72ef3515811d628ccbffa43b1013088ea2334e4fffd72735a021f7a554bcad9ce919323224173864f0c090f156ae5df7e4e982ae2884bdf610610d5d8c2b07e50e73f384da8bc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d82b2b7006e1370194b99a1a3c7e4435c076fdfdbd6e8f11966410ab012e4dc08681f3b5b5fe80434f62b9935ac9dbfb2fbcd9bf98ac30aea02e0179220bcdf1d1c4b11a30332b25c70322865555c9509c038ef5548a22507f8adadbe900e39de6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac1c18f62db3f3b27f75876f3888c0458a9ce8c064d05ede0943993e4070757fcb6e55a506e878021bff05a9f3d29937a9a44dbe801f003b82a5d154d0398028ce5a7674a30bdbf9ccc0653c78f2faec9347064ad2e8977a6a4ab52d95c7458968e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8abb5d7ac4e9dad4481e8c1c5aad02616b1b38995bab1a010d08b1733f12938ed02757a93283cfb44ff3130dea306a4b4619044fb010fbab033bba430b2215088b61e965d47293c1d6bd5c745f89c25f3906eea1eaba751ebe1c09bd1f052be909e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a9a218ab909ea89ef3b2d98bc50a60ea6bace57f607176dd0e2adbcb275525d98c1d19423fd6bd356f5e2e0216c916fdfe5da605cb27ae40236a61b6a1fa093dccbe5669c3b62454b9c3d4ec03c8fe5b03539c2110890df1f4b08fa407961953606;
        #1
        $finish();
    end
endmodule
