module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    compressor_CLA64_64 compressor_CLA64_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
        src16 <= 64'h0;
        src17 <= 64'h0;
        src18 <= 64'h0;
        src19 <= 64'h0;
        src20 <= 64'h0;
        src21 <= 64'h0;
        src22 <= 64'h0;
        src23 <= 64'h0;
        src24 <= 64'h0;
        src25 <= 64'h0;
        src26 <= 64'h0;
        src27 <= 64'h0;
        src28 <= 64'h0;
        src29 <= 64'h0;
        src30 <= 64'h0;
        src31 <= 64'h0;
        src32 <= 64'h0;
        src33 <= 64'h0;
        src34 <= 64'h0;
        src35 <= 64'h0;
        src36 <= 64'h0;
        src37 <= 64'h0;
        src38 <= 64'h0;
        src39 <= 64'h0;
        src40 <= 64'h0;
        src41 <= 64'h0;
        src42 <= 64'h0;
        src43 <= 64'h0;
        src44 <= 64'h0;
        src45 <= 64'h0;
        src46 <= 64'h0;
        src47 <= 64'h0;
        src48 <= 64'h0;
        src49 <= 64'h0;
        src50 <= 64'h0;
        src51 <= 64'h0;
        src52 <= 64'h0;
        src53 <= 64'h0;
        src54 <= 64'h0;
        src55 <= 64'h0;
        src56 <= 64'h0;
        src57 <= 64'h0;
        src58 <= 64'h0;
        src59 <= 64'h0;
        src60 <= 64'h0;
        src61 <= 64'h0;
        src62 <= 64'h0;
        src63 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA64_64(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    input [63:0]src16,
    input [63:0]src17,
    input [63:0]src18,
    input [63:0]src19,
    input [63:0]src20,
    input [63:0]src21,
    input [63:0]src22,
    input [63:0]src23,
    input [63:0]src24,
    input [63:0]src25,
    input [63:0]src26,
    input [63:0]src27,
    input [63:0]src28,
    input [63:0]src29,
    input [63:0]src30,
    input [63:0]src31,
    input [63:0]src32,
    input [63:0]src33,
    input [63:0]src34,
    input [63:0]src35,
    input [63:0]src36,
    input [63:0]src37,
    input [63:0]src38,
    input [63:0]src39,
    input [63:0]src40,
    input [63:0]src41,
    input [63:0]src42,
    input [63:0]src43,
    input [63:0]src44,
    input [63:0]src45,
    input [63:0]src46,
    input [63:0]src47,
    input [63:0]src48,
    input [63:0]src49,
    input [63:0]src50,
    input [63:0]src51,
    input [63:0]src52,
    input [63:0]src53,
    input [63:0]src54,
    input [63:0]src55,
    input [63:0]src56,
    input [63:0]src57,
    input [63:0]src58,
    input [63:0]src59,
    input [63:0]src60,
    input [63:0]src61,
    input [63:0]src62,
    input [63:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [0:0] comp_out67;
    wire [1:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out68[1], 1'h0, comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      input wire [63:0] src32,
      input wire [63:0] src33,
      input wire [63:0] src34,
      input wire [63:0] src35,
      input wire [63:0] src36,
      input wire [63:0] src37,
      input wire [63:0] src38,
      input wire [63:0] src39,
      input wire [63:0] src40,
      input wire [63:0] src41,
      input wire [63:0] src42,
      input wire [63:0] src43,
      input wire [63:0] src44,
      input wire [63:0] src45,
      input wire [63:0] src46,
      input wire [63:0] src47,
      input wire [63:0] src48,
      input wire [63:0] src49,
      input wire [63:0] src50,
      input wire [63:0] src51,
      input wire [63:0] src52,
      input wire [63:0] src53,
      input wire [63:0] src54,
      input wire [63:0] src55,
      input wire [63:0] src56,
      input wire [63:0] src57,
      input wire [63:0] src58,
      input wire [63:0] src59,
      input wire [63:0] src60,
      input wire [63:0] src61,
      input wire [63:0] src62,
      input wire [63:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [0:0] dst67,
      output wire [1:0] dst68,
      output wire [0:0] dst69);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [63:0] stage0_16;
   wire [63:0] stage0_17;
   wire [63:0] stage0_18;
   wire [63:0] stage0_19;
   wire [63:0] stage0_20;
   wire [63:0] stage0_21;
   wire [63:0] stage0_22;
   wire [63:0] stage0_23;
   wire [63:0] stage0_24;
   wire [63:0] stage0_25;
   wire [63:0] stage0_26;
   wire [63:0] stage0_27;
   wire [63:0] stage0_28;
   wire [63:0] stage0_29;
   wire [63:0] stage0_30;
   wire [63:0] stage0_31;
   wire [63:0] stage0_32;
   wire [63:0] stage0_33;
   wire [63:0] stage0_34;
   wire [63:0] stage0_35;
   wire [63:0] stage0_36;
   wire [63:0] stage0_37;
   wire [63:0] stage0_38;
   wire [63:0] stage0_39;
   wire [63:0] stage0_40;
   wire [63:0] stage0_41;
   wire [63:0] stage0_42;
   wire [63:0] stage0_43;
   wire [63:0] stage0_44;
   wire [63:0] stage0_45;
   wire [63:0] stage0_46;
   wire [63:0] stage0_47;
   wire [63:0] stage0_48;
   wire [63:0] stage0_49;
   wire [63:0] stage0_50;
   wire [63:0] stage0_51;
   wire [63:0] stage0_52;
   wire [63:0] stage0_53;
   wire [63:0] stage0_54;
   wire [63:0] stage0_55;
   wire [63:0] stage0_56;
   wire [63:0] stage0_57;
   wire [63:0] stage0_58;
   wire [63:0] stage0_59;
   wire [63:0] stage0_60;
   wire [63:0] stage0_61;
   wire [63:0] stage0_62;
   wire [63:0] stage0_63;
   wire [18:0] stage1_0;
   wire [47:0] stage1_1;
   wire [23:0] stage1_2;
   wire [27:0] stage1_3;
   wire [37:0] stage1_4;
   wire [26:0] stage1_5;
   wire [21:0] stage1_6;
   wire [35:0] stage1_7;
   wire [26:0] stage1_8;
   wire [28:0] stage1_9;
   wire [33:0] stage1_10;
   wire [32:0] stage1_11;
   wire [26:0] stage1_12;
   wire [30:0] stage1_13;
   wire [24:0] stage1_14;
   wire [44:0] stage1_15;
   wire [30:0] stage1_16;
   wire [44:0] stage1_17;
   wire [22:0] stage1_18;
   wire [28:0] stage1_19;
   wire [40:0] stage1_20;
   wire [32:0] stage1_21;
   wire [30:0] stage1_22;
   wire [34:0] stage1_23;
   wire [26:0] stage1_24;
   wire [44:0] stage1_25;
   wire [28:0] stage1_26;
   wire [40:0] stage1_27;
   wire [26:0] stage1_28;
   wire [28:0] stage1_29;
   wire [25:0] stage1_30;
   wire [22:0] stage1_31;
   wire [30:0] stage1_32;
   wire [37:0] stage1_33;
   wire [23:0] stage1_34;
   wire [29:0] stage1_35;
   wire [43:0] stage1_36;
   wire [23:0] stage1_37;
   wire [41:0] stage1_38;
   wire [22:0] stage1_39;
   wire [26:0] stage1_40;
   wire [35:0] stage1_41;
   wire [28:0] stage1_42;
   wire [35:0] stage1_43;
   wire [32:0] stage1_44;
   wire [47:0] stage1_45;
   wire [16:0] stage1_46;
   wire [40:0] stage1_47;
   wire [31:0] stage1_48;
   wire [24:0] stage1_49;
   wire [24:0] stage1_50;
   wire [31:0] stage1_51;
   wire [42:0] stage1_52;
   wire [26:0] stage1_53;
   wire [32:0] stage1_54;
   wire [24:0] stage1_55;
   wire [25:0] stage1_56;
   wire [25:0] stage1_57;
   wire [40:0] stage1_58;
   wire [41:0] stage1_59;
   wire [32:0] stage1_60;
   wire [30:0] stage1_61;
   wire [32:0] stage1_62;
   wire [27:0] stage1_63;
   wire [15:0] stage1_64;
   wire [8:0] stage1_65;
   wire [5:0] stage2_0;
   wire [8:0] stage2_1;
   wire [11:0] stage2_2;
   wire [11:0] stage2_3;
   wire [25:0] stage2_4;
   wire [21:0] stage2_5;
   wire [13:0] stage2_6;
   wire [19:0] stage2_7;
   wire [19:0] stage2_8;
   wire [10:0] stage2_9;
   wire [30:0] stage2_10;
   wire [15:0] stage2_11;
   wire [18:0] stage2_12;
   wire [8:0] stage2_13;
   wire [15:0] stage2_14;
   wire [20:0] stage2_15;
   wire [15:0] stage2_16;
   wire [21:0] stage2_17;
   wire [18:0] stage2_18;
   wire [14:0] stage2_19;
   wire [23:0] stage2_20;
   wire [12:0] stage2_21;
   wire [10:0] stage2_22;
   wire [16:0] stage2_23;
   wire [13:0] stage2_24;
   wire [13:0] stage2_25;
   wire [19:0] stage2_26;
   wire [25:0] stage2_27;
   wire [15:0] stage2_28;
   wire [9:0] stage2_29;
   wire [19:0] stage2_30;
   wire [12:0] stage2_31;
   wire [18:0] stage2_32;
   wire [22:0] stage2_33;
   wire [12:0] stage2_34;
   wire [12:0] stage2_35;
   wire [17:0] stage2_36;
   wire [17:0] stage2_37;
   wire [23:0] stage2_38;
   wire [12:0] stage2_39;
   wire [11:0] stage2_40;
   wire [19:0] stage2_41;
   wire [14:0] stage2_42;
   wire [12:0] stage2_43;
   wire [17:0] stage2_44;
   wire [13:0] stage2_45;
   wire [11:0] stage2_46;
   wire [18:0] stage2_47;
   wire [16:0] stage2_48;
   wire [10:0] stage2_49;
   wire [11:0] stage2_50;
   wire [15:0] stage2_51;
   wire [11:0] stage2_52;
   wire [17:0] stage2_53;
   wire [14:0] stage2_54;
   wire [16:0] stage2_55;
   wire [9:0] stage2_56;
   wire [13:0] stage2_57;
   wire [17:0] stage2_58;
   wire [19:0] stage2_59;
   wire [13:0] stage2_60;
   wire [14:0] stage2_61;
   wire [12:0] stage2_62;
   wire [12:0] stage2_63;
   wire [10:0] stage2_64;
   wire [7:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage2_67;
   wire [5:0] stage3_0;
   wire [3:0] stage3_1;
   wire [2:0] stage3_2;
   wire [4:0] stage3_3;
   wire [6:0] stage3_4;
   wire [8:0] stage3_5;
   wire [7:0] stage3_6;
   wire [10:0] stage3_7;
   wire [8:0] stage3_8;
   wire [11:0] stage3_9;
   wire [6:0] stage3_10;
   wire [8:0] stage3_11;
   wire [7:0] stage3_12;
   wire [8:0] stage3_13;
   wire [6:0] stage3_14;
   wire [8:0] stage3_15;
   wire [7:0] stage3_16;
   wire [6:0] stage3_17;
   wire [12:0] stage3_18;
   wire [6:0] stage3_19;
   wire [5:0] stage3_20;
   wire [8:0] stage3_21;
   wire [6:0] stage3_22;
   wire [7:0] stage3_23;
   wire [6:0] stage3_24;
   wire [7:0] stage3_25;
   wire [6:0] stage3_26;
   wire [6:0] stage3_27;
   wire [8:0] stage3_28;
   wire [8:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [6:0] stage3_32;
   wire [16:0] stage3_33;
   wire [6:0] stage3_34;
   wire [5:0] stage3_35;
   wire [9:0] stage3_36;
   wire [5:0] stage3_37;
   wire [10:0] stage3_38;
   wire [6:0] stage3_39;
   wire [5:0] stage3_40;
   wire [13:0] stage3_41;
   wire [3:0] stage3_42;
   wire [5:0] stage3_43;
   wire [16:0] stage3_44;
   wire [4:0] stage3_45;
   wire [6:0] stage3_46;
   wire [8:0] stage3_47;
   wire [5:0] stage3_48;
   wire [5:0] stage3_49;
   wire [6:0] stage3_50;
   wire [8:0] stage3_51;
   wire [6:0] stage3_52;
   wire [5:0] stage3_53;
   wire [5:0] stage3_54;
   wire [9:0] stage3_55;
   wire [5:0] stage3_56;
   wire [7:0] stage3_57;
   wire [7:0] stage3_58;
   wire [7:0] stage3_59;
   wire [13:0] stage3_60;
   wire [6:0] stage3_61;
   wire [4:0] stage3_62;
   wire [5:0] stage3_63;
   wire [4:0] stage3_64;
   wire [5:0] stage3_65;
   wire [2:0] stage3_66;
   wire [2:0] stage3_67;
   wire [0:0] stage3_68;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [2:0] stage4_2;
   wire [1:0] stage4_3;
   wire [3:0] stage4_4;
   wire [1:0] stage4_5;
   wire [2:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [4:0] stage4_11;
   wire [2:0] stage4_12;
   wire [3:0] stage4_13;
   wire [3:0] stage4_14;
   wire [3:0] stage4_15;
   wire [4:0] stage4_16;
   wire [2:0] stage4_17;
   wire [3:0] stage4_18;
   wire [2:0] stage4_19;
   wire [3:0] stage4_20;
   wire [7:0] stage4_21;
   wire [1:0] stage4_22;
   wire [3:0] stage4_23;
   wire [3:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [3:0] stage4_27;
   wire [3:0] stage4_28;
   wire [3:0] stage4_29;
   wire [2:0] stage4_30;
   wire [2:0] stage4_31;
   wire [3:0] stage4_32;
   wire [5:0] stage4_33;
   wire [4:0] stage4_34;
   wire [2:0] stage4_35;
   wire [3:0] stage4_36;
   wire [4:0] stage4_37;
   wire [2:0] stage4_38;
   wire [2:0] stage4_39;
   wire [2:0] stage4_40;
   wire [3:0] stage4_41;
   wire [3:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [2:0] stage4_45;
   wire [3:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [3:0] stage4_49;
   wire [3:0] stage4_50;
   wire [5:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [2:0] stage4_54;
   wire [6:0] stage4_55;
   wire [1:0] stage4_56;
   wire [3:0] stage4_57;
   wire [5:0] stage4_58;
   wire [2:0] stage4_59;
   wire [5:0] stage4_60;
   wire [4:0] stage4_61;
   wire [2:0] stage4_62;
   wire [1:0] stage4_63;
   wire [6:0] stage4_64;
   wire [2:0] stage4_65;
   wire [1:0] stage4_66;
   wire [0:0] stage4_67;
   wire [0:0] stage4_68;
   wire [0:0] stage4_69;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [0:0] stage5_67;
   wire [1:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc615_5 gpc14 (
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[5],stage1_4[14],stage1_3[14]}
   );
   gpc615_5 gpc15 (
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[6],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[7],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[8],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc18 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[5],stage1_5[10],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[6],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[7],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[8],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[9],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[10],stage1_5[15],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[11],stage1_5[16],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[12],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[13],stage1_6[13],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[14],stage1_6[14],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[15],stage1_6[15],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[16],stage1_6[16],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[17],stage1_6[17],stage1_5[22]}
   );
   gpc615_5 gpc32 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[30]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[5],stage1_8[13],stage1_7[18],stage1_6[18]}
   );
   gpc615_5 gpc33 (
      {stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_7[31]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[6],stage1_8[14],stage1_7[19],stage1_6[19]}
   );
   gpc615_5 gpc34 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62]},
      {stage0_7[32]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[7],stage1_8[15],stage1_7[20],stage1_6[20]}
   );
   gpc615_5 gpc35 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[8],stage1_8[16],stage1_7[21]}
   );
   gpc615_5 gpc36 (
      {stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42]},
      {stage0_8[19]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[9],stage1_8[17],stage1_7[22]}
   );
   gpc615_5 gpc37 (
      {stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage0_8[20]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[10],stage1_8[18],stage1_7[23]}
   );
   gpc615_5 gpc38 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52]},
      {stage0_8[21]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[11],stage1_8[19],stage1_7[24]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[4],stage1_10[7],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[5],stage1_10[8],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[6],stage1_10[9],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc42 (
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[7],stage1_10[10],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc43 (
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[8],stage1_10[11],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc44 (
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[9],stage1_10[12],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc45 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[10],stage1_10[13],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc46 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[11],stage1_10[14],stage1_9[19]}
   );
   gpc606_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[12],stage1_10[15],stage1_9[20]}
   );
   gpc606_5 gpc48 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[13],stage1_10[16],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[14],stage1_10[17],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[15],stage1_10[18],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[16],stage1_10[19],stage1_9[24]}
   );
   gpc615_5 gpc52 (
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46]},
      {stage0_11[36]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[6],stage1_12[13],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc53 (
      {stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51]},
      {stage0_11[37]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[7],stage1_12[14],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc54 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[8],stage1_12[15],stage1_11[19]}
   );
   gpc615_5 gpc55 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[9],stage1_12[16],stage1_11[20]}
   );
   gpc615_5 gpc56 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52]},
      {stage0_12[14]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[4],stage1_13[10],stage1_12[17],stage1_11[21]}
   );
   gpc606_5 gpc57 (
      {stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[3],stage1_14[5],stage1_13[11],stage1_12[18]}
   );
   gpc606_5 gpc58 (
      {stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[4],stage1_14[6],stage1_13[12],stage1_12[19]}
   );
   gpc606_5 gpc59 (
      {stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[5],stage1_14[7],stage1_13[13],stage1_12[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[6],stage1_14[8],stage1_13[14],stage1_12[21]}
   );
   gpc606_5 gpc61 (
      {stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[7],stage1_14[9],stage1_13[15],stage1_12[22]}
   );
   gpc606_5 gpc62 (
      {stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[8],stage1_14[10],stage1_13[16],stage1_12[23]}
   );
   gpc606_5 gpc63 (
      {stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[9],stage1_14[11],stage1_13[17],stage1_12[24]}
   );
   gpc606_5 gpc64 (
      {stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[10],stage1_14[12],stage1_13[18],stage1_12[25]}
   );
   gpc2135_5 gpc65 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22]},
      {stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[0]},
      {stage0_16[0], stage0_16[1]},
      {stage1_17[0],stage1_16[8],stage1_15[11],stage1_14[13],stage1_13[19]}
   );
   gpc606_5 gpc66 (
      {stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[1],stage1_16[9],stage1_15[12],stage1_14[14],stage1_13[20]}
   );
   gpc606_5 gpc67 (
      {stage0_13[29], stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[2],stage1_16[10],stage1_15[13],stage1_14[15],stage1_13[21]}
   );
   gpc606_5 gpc68 (
      {stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[3],stage1_16[11],stage1_15[14],stage1_14[16],stage1_13[22]}
   );
   gpc606_5 gpc69 (
      {stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage1_17[4],stage1_16[12],stage1_15[15],stage1_14[17],stage1_13[23]}
   );
   gpc606_5 gpc70 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52]},
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30]},
      {stage1_17[5],stage1_16[13],stage1_15[16],stage1_14[18],stage1_13[24]}
   );
   gpc606_5 gpc71 (
      {stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58]},
      {stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36]},
      {stage1_17[6],stage1_16[14],stage1_15[17],stage1_14[19],stage1_13[25]}
   );
   gpc615_5 gpc72 (
      {stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage0_15[37]},
      {stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7]},
      {stage1_18[0],stage1_17[7],stage1_16[15],stage1_15[18],stage1_14[20]}
   );
   gpc615_5 gpc73 (
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage0_15[38]},
      {stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13]},
      {stage1_18[1],stage1_17[8],stage1_16[16],stage1_15[19],stage1_14[21]}
   );
   gpc606_5 gpc74 (
      {stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[9],stage1_16[17]}
   );
   gpc606_5 gpc75 (
      {stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[10],stage1_16[18]}
   );
   gpc606_5 gpc76 (
      {stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[2],stage1_18[4],stage1_17[11],stage1_16[19]}
   );
   gpc606_5 gpc77 (
      {stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[3],stage1_18[5],stage1_17[12],stage1_16[20]}
   );
   gpc615_5 gpc78 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_17[0]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[4],stage1_18[6],stage1_17[13],stage1_16[21]}
   );
   gpc615_5 gpc79 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage0_17[1]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[5],stage1_18[7],stage1_17[14],stage1_16[22]}
   );
   gpc615_5 gpc80 (
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52]},
      {stage0_17[2]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[6],stage1_18[8],stage1_17[15],stage1_16[23]}
   );
   gpc615_5 gpc81 (
      {stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage0_17[3]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[7],stage1_18[9],stage1_17[16],stage1_16[24]}
   );
   gpc606_5 gpc82 (
      {stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[8],stage1_19[8],stage1_18[10],stage1_17[17]}
   );
   gpc606_5 gpc83 (
      {stage0_17[10], stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[9],stage1_19[9],stage1_18[11],stage1_17[18]}
   );
   gpc606_5 gpc84 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[10],stage1_19[10],stage1_18[12],stage1_17[19]}
   );
   gpc606_5 gpc85 (
      {stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[11],stage1_19[11],stage1_18[13],stage1_17[20]}
   );
   gpc606_5 gpc86 (
      {stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[12],stage1_19[12],stage1_18[14],stage1_17[21]}
   );
   gpc606_5 gpc87 (
      {stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[13],stage1_19[13],stage1_18[15],stage1_17[22]}
   );
   gpc623_5 gpc88 (
      {stage0_17[40], stage0_17[41], stage0_17[42]},
      {stage0_18[48], stage0_18[49]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[14],stage1_19[14],stage1_18[16],stage1_17[23]}
   );
   gpc615_5 gpc89 (
      {stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53], stage0_18[54]},
      {stage0_19[42]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[7],stage1_20[15],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc90 (
      {stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage0_19[43]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[8],stage1_20[16],stage1_19[16],stage1_18[18]}
   );
   gpc615_5 gpc91 (
      {stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[9],stage1_20[17],stage1_19[17]}
   );
   gpc615_5 gpc92 (
      {stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage0_20[13]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[3],stage1_21[10],stage1_20[18],stage1_19[18]}
   );
   gpc615_5 gpc93 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[4],stage1_21[11],stage1_20[19]}
   );
   gpc615_5 gpc94 (
      {stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[5],stage1_21[12],stage1_20[20]}
   );
   gpc615_5 gpc95 (
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[6],stage1_21[13],stage1_20[21]}
   );
   gpc615_5 gpc96 (
      {stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[7],stage1_21[14],stage1_20[22]}
   );
   gpc615_5 gpc97 (
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[8],stage1_21[15],stage1_20[23]}
   );
   gpc615_5 gpc98 (
      {stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[9],stage1_21[16],stage1_20[24]}
   );
   gpc615_5 gpc99 (
      {stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47], stage0_20[48]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[10],stage1_21[17],stage1_20[25]}
   );
   gpc606_5 gpc100 (
      {stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[7],stage1_23[9],stage1_22[11],stage1_21[18]}
   );
   gpc606_5 gpc101 (
      {stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[8],stage1_23[10],stage1_22[12],stage1_21[19]}
   );
   gpc606_5 gpc102 (
      {stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[9],stage1_23[11],stage1_22[13],stage1_21[20]}
   );
   gpc606_5 gpc103 (
      {stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[10],stage1_23[12],stage1_22[14],stage1_21[21]}
   );
   gpc606_5 gpc104 (
      {stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[11],stage1_23[13],stage1_22[15],stage1_21[22]}
   );
   gpc606_5 gpc105 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[12],stage1_23[14],stage1_22[16],stage1_21[23]}
   );
   gpc615_5 gpc106 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46]},
      {stage0_23[36]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[6],stage1_24[13],stage1_23[15],stage1_22[17]}
   );
   gpc615_5 gpc107 (
      {stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51]},
      {stage0_23[37]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[7],stage1_24[14],stage1_23[16],stage1_22[18]}
   );
   gpc615_5 gpc108 (
      {stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage0_24[12]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[2],stage1_25[8],stage1_24[15],stage1_23[17]}
   );
   gpc615_5 gpc109 (
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage0_24[13]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[3],stage1_25[9],stage1_24[16],stage1_23[18]}
   );
   gpc606_5 gpc110 (
      {stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18], stage0_24[19]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[4],stage1_25[10],stage1_24[17]}
   );
   gpc606_5 gpc111 (
      {stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24], stage0_24[25]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[5],stage1_25[11],stage1_24[18]}
   );
   gpc606_5 gpc112 (
      {stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[6],stage1_25[12],stage1_24[19]}
   );
   gpc606_5 gpc113 (
      {stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36], stage0_24[37]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[7],stage1_25[13],stage1_24[20]}
   );
   gpc606_5 gpc114 (
      {stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42], stage0_24[43]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[8],stage1_25[14],stage1_24[21]}
   );
   gpc606_5 gpc115 (
      {stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47], stage0_24[48], stage0_24[49]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[9],stage1_25[15],stage1_24[22]}
   );
   gpc606_5 gpc116 (
      {stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53], stage0_24[54], stage0_24[55]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[10],stage1_25[16],stage1_24[23]}
   );
   gpc606_5 gpc117 (
      {stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59], stage0_24[60], stage0_24[61]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[11],stage1_25[17],stage1_24[24]}
   );
   gpc606_5 gpc118 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[10],stage1_26[12],stage1_25[18]}
   );
   gpc606_5 gpc119 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[11],stage1_26[13],stage1_25[19]}
   );
   gpc606_5 gpc120 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[12],stage1_26[14],stage1_25[20]}
   );
   gpc606_5 gpc121 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[13],stage1_26[15],stage1_25[21]}
   );
   gpc606_5 gpc122 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[14],stage1_26[16],stage1_25[22]}
   );
   gpc615_5 gpc123 (
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52]},
      {stage0_27[30]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[5],stage1_28[13],stage1_27[15],stage1_26[17]}
   );
   gpc615_5 gpc124 (
      {stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage0_28[6]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[6],stage1_28[14],stage1_27[16]}
   );
   gpc615_5 gpc125 (
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40]},
      {stage0_28[7]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[2],stage1_29[7],stage1_28[15],stage1_27[17]}
   );
   gpc606_5 gpc126 (
      {stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[3],stage1_29[8],stage1_28[16]}
   );
   gpc606_5 gpc127 (
      {stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[3],stage1_30[4],stage1_29[9],stage1_28[17]}
   );
   gpc606_5 gpc128 (
      {stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[4],stage1_30[5],stage1_29[10],stage1_28[18]}
   );
   gpc606_5 gpc129 (
      {stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[5],stage1_30[6],stage1_29[11],stage1_28[19]}
   );
   gpc606_5 gpc130 (
      {stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36], stage0_28[37]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[6],stage1_30[7],stage1_29[12],stage1_28[20]}
   );
   gpc606_5 gpc131 (
      {stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42], stage0_28[43]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[7],stage1_30[8],stage1_29[13],stage1_28[21]}
   );
   gpc606_5 gpc132 (
      {stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48], stage0_28[49]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[8],stage1_30[9],stage1_29[14],stage1_28[22]}
   );
   gpc606_5 gpc133 (
      {stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], stage0_28[54], stage0_28[55]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[9],stage1_30[10],stage1_29[15],stage1_28[23]}
   );
   gpc606_5 gpc134 (
      {stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59], stage0_28[60], stage0_28[61]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[10],stage1_30[11],stage1_29[16],stage1_28[24]}
   );
   gpc606_5 gpc135 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[11],stage1_30[12],stage1_29[17]}
   );
   gpc606_5 gpc136 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[12],stage1_30[13],stage1_29[18]}
   );
   gpc606_5 gpc137 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[13],stage1_30[14],stage1_29[19]}
   );
   gpc606_5 gpc138 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[14],stage1_30[15],stage1_29[20]}
   );
   gpc606_5 gpc139 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[15],stage1_30[16],stage1_29[21]}
   );
   gpc606_5 gpc140 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[16],stage1_30[17],stage1_29[22]}
   );
   gpc606_5 gpc141 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[17],stage1_30[18],stage1_29[23]}
   );
   gpc606_5 gpc142 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[18],stage1_30[19],stage1_29[24]}
   );
   gpc615_5 gpc143 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58]},
      {stage0_31[48]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[8],stage1_32[17],stage1_31[19],stage1_30[20]}
   );
   gpc615_5 gpc144 (
      {stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage0_32[6]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[1],stage1_33[9],stage1_32[18],stage1_31[20]}
   );
   gpc615_5 gpc145 (
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58]},
      {stage0_32[7]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[2],stage1_33[10],stage1_32[19],stage1_31[21]}
   );
   gpc615_5 gpc146 (
      {stage0_31[59], stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63]},
      {stage0_32[8]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[3],stage1_33[11],stage1_32[20],stage1_31[22]}
   );
   gpc606_5 gpc147 (
      {stage0_32[9], stage0_32[10], stage0_32[11], stage0_32[12], stage0_32[13], stage0_32[14]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[3],stage1_34[4],stage1_33[12],stage1_32[21]}
   );
   gpc606_5 gpc148 (
      {stage0_32[15], stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[4],stage1_34[5],stage1_33[13],stage1_32[22]}
   );
   gpc606_5 gpc149 (
      {stage0_32[21], stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[5],stage1_34[6],stage1_33[14],stage1_32[23]}
   );
   gpc606_5 gpc150 (
      {stage0_32[27], stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[6],stage1_34[7],stage1_33[15],stage1_32[24]}
   );
   gpc606_5 gpc151 (
      {stage0_32[33], stage0_32[34], stage0_32[35], stage0_32[36], stage0_32[37], stage0_32[38]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[7],stage1_34[8],stage1_33[16],stage1_32[25]}
   );
   gpc606_5 gpc152 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[8],stage1_34[9],stage1_33[17],stage1_32[26]}
   );
   gpc606_5 gpc153 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[9],stage1_34[10],stage1_33[18],stage1_32[27]}
   );
   gpc606_5 gpc154 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[10],stage1_34[11],stage1_33[19],stage1_32[28]}
   );
   gpc606_5 gpc155 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[11],stage1_34[12],stage1_33[20],stage1_32[29]}
   );
   gpc606_5 gpc156 (
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[9],stage1_35[12],stage1_34[13],stage1_33[21]}
   );
   gpc606_5 gpc157 (
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[10],stage1_35[13],stage1_34[14],stage1_33[22]}
   );
   gpc606_5 gpc158 (
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[11],stage1_35[14],stage1_34[15],stage1_33[23]}
   );
   gpc606_5 gpc159 (
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[12],stage1_35[15],stage1_34[16],stage1_33[24]}
   );
   gpc606_5 gpc160 (
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[13],stage1_35[16],stage1_34[17],stage1_33[25]}
   );
   gpc615_5 gpc161 (
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52]},
      {stage0_34[54]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[14],stage1_35[17],stage1_34[18],stage1_33[26]}
   );
   gpc615_5 gpc162 (
      {stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage0_35[36]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[6],stage1_36[15],stage1_35[18],stage1_34[19]}
   );
   gpc615_5 gpc163 (
      {stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage0_36[6]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[1],stage1_37[7],stage1_36[16],stage1_35[19]}
   );
   gpc615_5 gpc164 (
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46]},
      {stage0_36[7]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[2],stage1_37[8],stage1_36[17],stage1_35[20]}
   );
   gpc615_5 gpc165 (
      {stage0_35[47], stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51]},
      {stage0_36[8]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[3],stage1_37[9],stage1_36[18],stage1_35[21]}
   );
   gpc615_5 gpc166 (
      {stage0_35[52], stage0_35[53], stage0_35[54], stage0_35[55], stage0_35[56]},
      {stage0_36[9]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[4],stage1_37[10],stage1_36[19],stage1_35[22]}
   );
   gpc606_5 gpc167 (
      {stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[4],stage1_38[5],stage1_37[11],stage1_36[20]}
   );
   gpc606_5 gpc168 (
      {stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[5],stage1_38[6],stage1_37[12],stage1_36[21]}
   );
   gpc606_5 gpc169 (
      {stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[6],stage1_38[7],stage1_37[13],stage1_36[22]}
   );
   gpc606_5 gpc170 (
      {stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[7],stage1_38[8],stage1_37[14],stage1_36[23]}
   );
   gpc606_5 gpc171 (
      {stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[8],stage1_38[9],stage1_37[15],stage1_36[24]}
   );
   gpc606_5 gpc172 (
      {stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[9],stage1_38[10],stage1_37[16],stage1_36[25]}
   );
   gpc606_5 gpc173 (
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[10],stage1_38[11],stage1_37[17]}
   );
   gpc606_5 gpc174 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[11],stage1_38[12],stage1_37[18]}
   );
   gpc606_5 gpc175 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[12],stage1_38[13],stage1_37[19]}
   );
   gpc606_5 gpc176 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[9],stage1_39[13],stage1_38[14],stage1_37[20]}
   );
   gpc606_5 gpc177 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[10],stage1_39[14],stage1_38[15],stage1_37[21]}
   );
   gpc606_5 gpc178 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[11],stage1_39[15],stage1_38[16],stage1_37[22]}
   );
   gpc606_5 gpc179 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], 1'b0, 1'b0},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[12],stage1_39[16],stage1_38[17],stage1_37[23]}
   );
   gpc615_5 gpc180 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[13],stage1_39[17],stage1_38[18]}
   );
   gpc615_5 gpc181 (
      {stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage0_40[6]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[8],stage1_40[14],stage1_39[18]}
   );
   gpc615_5 gpc182 (
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52]},
      {stage0_40[7]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[2],stage1_41[9],stage1_40[15],stage1_39[19]}
   );
   gpc615_5 gpc183 (
      {stage0_39[53], stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57]},
      {stage0_40[8]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[3],stage1_41[10],stage1_40[16],stage1_39[20]}
   );
   gpc615_5 gpc184 (
      {stage0_39[58], stage0_39[59], stage0_39[60], stage0_39[61], stage0_39[62]},
      {stage0_40[9]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[4],stage1_41[11],stage1_40[17],stage1_39[21]}
   );
   gpc606_5 gpc185 (
      {stage0_40[10], stage0_40[11], stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[4],stage1_42[5],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc186 (
      {stage0_40[16], stage0_40[17], stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[5],stage1_42[6],stage1_41[13],stage1_40[19]}
   );
   gpc606_5 gpc187 (
      {stage0_40[22], stage0_40[23], stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[6],stage1_42[7],stage1_41[14],stage1_40[20]}
   );
   gpc606_5 gpc188 (
      {stage0_40[28], stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[7],stage1_42[8],stage1_41[15],stage1_40[21]}
   );
   gpc606_5 gpc189 (
      {stage0_40[34], stage0_40[35], stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[8],stage1_42[9],stage1_41[16],stage1_40[22]}
   );
   gpc606_5 gpc190 (
      {stage0_40[40], stage0_40[41], stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[9],stage1_42[10],stage1_41[17],stage1_40[23]}
   );
   gpc606_5 gpc191 (
      {stage0_40[46], stage0_40[47], stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[10],stage1_42[11],stage1_41[18],stage1_40[24]}
   );
   gpc606_5 gpc192 (
      {stage0_40[52], stage0_40[53], stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[11],stage1_42[12],stage1_41[19],stage1_40[25]}
   );
   gpc606_5 gpc193 (
      {stage0_40[58], stage0_40[59], stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[12],stage1_42[13],stage1_41[20],stage1_40[26]}
   );
   gpc606_5 gpc194 (
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[9],stage1_43[13],stage1_42[14],stage1_41[21]}
   );
   gpc606_5 gpc195 (
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[10],stage1_43[14],stage1_42[15],stage1_41[22]}
   );
   gpc606_5 gpc196 (
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[11],stage1_43[15],stage1_42[16],stage1_41[23]}
   );
   gpc606_5 gpc197 (
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[12],stage1_43[16],stage1_42[17],stage1_41[24]}
   );
   gpc606_5 gpc198 (
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[13],stage1_43[17],stage1_42[18],stage1_41[25]}
   );
   gpc615_5 gpc199 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[0]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[0],stage1_45[5],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc200 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[1]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[1],stage1_45[6],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc201 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[2]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[2],stage1_45[7],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc202 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[3]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[3],stage1_45[8],stage1_44[17],stage1_43[21]}
   );
   gpc606_5 gpc203 (
      {stage0_44[4], stage0_44[5], stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[4],stage1_46[4],stage1_45[9],stage1_44[18]}
   );
   gpc606_5 gpc204 (
      {stage0_44[10], stage0_44[11], stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[5],stage1_46[5],stage1_45[10],stage1_44[19]}
   );
   gpc606_5 gpc205 (
      {stage0_44[16], stage0_44[17], stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[6],stage1_46[6],stage1_45[11],stage1_44[20]}
   );
   gpc606_5 gpc206 (
      {stage0_44[22], stage0_44[23], stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[7],stage1_46[7],stage1_45[12],stage1_44[21]}
   );
   gpc606_5 gpc207 (
      {stage0_44[28], stage0_44[29], stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[8],stage1_46[8],stage1_45[13],stage1_44[22]}
   );
   gpc606_5 gpc208 (
      {stage0_44[34], stage0_44[35], stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[9],stage1_46[9],stage1_45[14],stage1_44[23]}
   );
   gpc606_5 gpc209 (
      {stage0_44[40], stage0_44[41], stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[10],stage1_46[10],stage1_45[15],stage1_44[24]}
   );
   gpc606_5 gpc210 (
      {stage0_44[46], stage0_44[47], stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[11],stage1_46[11],stage1_45[16],stage1_44[25]}
   );
   gpc606_5 gpc211 (
      {stage0_44[52], stage0_44[53], stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[12],stage1_46[12],stage1_45[17],stage1_44[26]}
   );
   gpc606_5 gpc212 (
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[9],stage1_47[13],stage1_46[13],stage1_45[18]}
   );
   gpc606_5 gpc213 (
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[10],stage1_47[14],stage1_46[14],stage1_45[19]}
   );
   gpc615_5 gpc214 (
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58]},
      {stage0_47[12]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[2],stage1_48[11],stage1_47[15],stage1_46[15]}
   );
   gpc615_5 gpc215 (
      {stage0_46[59], stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63]},
      {stage0_47[13]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[3],stage1_48[12],stage1_47[16],stage1_46[16]}
   );
   gpc606_5 gpc216 (
      {stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[2],stage1_49[4],stage1_48[13],stage1_47[17]}
   );
   gpc606_5 gpc217 (
      {stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[3],stage1_49[5],stage1_48[14],stage1_47[18]}
   );
   gpc615_5 gpc218 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[12]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[4],stage1_49[6],stage1_48[15],stage1_47[19]}
   );
   gpc615_5 gpc219 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[13]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[5],stage1_49[7],stage1_48[16],stage1_47[20]}
   );
   gpc615_5 gpc220 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[14]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[6],stage1_49[8],stage1_48[17],stage1_47[21]}
   );
   gpc615_5 gpc221 (
      {stage0_47[41], stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45]},
      {stage0_48[15]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[7],stage1_49[9],stage1_48[18],stage1_47[22]}
   );
   gpc606_5 gpc222 (
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[8],stage1_49[10],stage1_48[19]}
   );
   gpc606_5 gpc223 (
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[9],stage1_49[11],stage1_48[20]}
   );
   gpc606_5 gpc224 (
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[10],stage1_49[12],stage1_48[21]}
   );
   gpc606_5 gpc225 (
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[9],stage1_50[11],stage1_49[13],stage1_48[22]}
   );
   gpc606_5 gpc226 (
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[10],stage1_50[12],stage1_49[14],stage1_48[23]}
   );
   gpc606_5 gpc227 (
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[11],stage1_50[13],stage1_49[15],stage1_48[24]}
   );
   gpc606_5 gpc228 (
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[12],stage1_50[14],stage1_49[16],stage1_48[25]}
   );
   gpc606_5 gpc229 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[7],stage1_51[13],stage1_50[15],stage1_49[17]}
   );
   gpc606_5 gpc230 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[8],stage1_51[14],stage1_50[16],stage1_49[18]}
   );
   gpc606_5 gpc231 (
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[9],stage1_51[15],stage1_50[17],stage1_49[19]}
   );
   gpc606_5 gpc232 (
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[10],stage1_51[16],stage1_50[18],stage1_49[20]}
   );
   gpc615_5 gpc233 (
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46]},
      {stage0_51[24]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[4],stage1_52[11],stage1_51[17],stage1_50[19]}
   );
   gpc615_5 gpc234 (
      {stage0_50[47], stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51]},
      {stage0_51[25]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[5],stage1_52[12],stage1_51[18],stage1_50[20]}
   );
   gpc615_5 gpc235 (
      {stage0_50[52], stage0_50[53], stage0_50[54], stage0_50[55], stage0_50[56]},
      {stage0_51[26]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[6],stage1_52[13],stage1_51[19],stage1_50[21]}
   );
   gpc615_5 gpc236 (
      {stage0_50[57], stage0_50[58], stage0_50[59], stage0_50[60], stage0_50[61]},
      {stage0_51[27]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[7],stage1_52[14],stage1_51[20],stage1_50[22]}
   );
   gpc606_5 gpc237 (
      {stage0_51[28], stage0_51[29], stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[8],stage1_52[15],stage1_51[21]}
   );
   gpc615_5 gpc238 (
      {stage0_51[34], stage0_51[35], stage0_51[36], stage0_51[37], stage0_51[38]},
      {stage0_52[24]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[9],stage1_52[16],stage1_51[22]}
   );
   gpc615_5 gpc239 (
      {stage0_51[39], stage0_51[40], stage0_51[41], stage0_51[42], stage0_51[43]},
      {stage0_52[25]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[10],stage1_52[17],stage1_51[23]}
   );
   gpc615_5 gpc240 (
      {stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47], stage0_51[48]},
      {stage0_52[26]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[11],stage1_52[18],stage1_51[24]}
   );
   gpc615_5 gpc241 (
      {stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage0_52[27]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[12],stage1_52[19],stage1_51[25]}
   );
   gpc615_5 gpc242 (
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58]},
      {stage0_52[28]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[13],stage1_52[20],stage1_51[26]}
   );
   gpc606_5 gpc243 (
      {stage0_52[29], stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[6],stage1_54[10],stage1_53[14],stage1_52[21]}
   );
   gpc615_5 gpc244 (
      {stage0_52[35], stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39]},
      {stage0_53[36]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[7],stage1_54[11],stage1_53[15],stage1_52[22]}
   );
   gpc615_5 gpc245 (
      {stage0_52[40], stage0_52[41], stage0_52[42], stage0_52[43], stage0_52[44]},
      {stage0_53[37]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[8],stage1_54[12],stage1_53[16],stage1_52[23]}
   );
   gpc615_5 gpc246 (
      {stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41], stage0_53[42]},
      {stage0_54[18]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[3],stage1_55[9],stage1_54[13],stage1_53[17]}
   );
   gpc615_5 gpc247 (
      {stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage0_54[19]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[4],stage1_55[10],stage1_54[14],stage1_53[18]}
   );
   gpc615_5 gpc248 (
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52]},
      {stage0_54[20]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[5],stage1_55[11],stage1_54[15],stage1_53[19]}
   );
   gpc615_5 gpc249 (
      {stage0_53[53], stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57]},
      {stage0_54[21]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[6],stage1_55[12],stage1_54[16],stage1_53[20]}
   );
   gpc606_5 gpc250 (
      {stage0_54[22], stage0_54[23], stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[4],stage1_56[7],stage1_55[13],stage1_54[17]}
   );
   gpc606_5 gpc251 (
      {stage0_54[28], stage0_54[29], stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[5],stage1_56[8],stage1_55[14],stage1_54[18]}
   );
   gpc615_5 gpc252 (
      {stage0_54[34], stage0_54[35], stage0_54[36], stage0_54[37], stage0_54[38]},
      {stage0_55[24]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[6],stage1_56[9],stage1_55[15],stage1_54[19]}
   );
   gpc615_5 gpc253 (
      {stage0_54[39], stage0_54[40], stage0_54[41], stage0_54[42], stage0_54[43]},
      {stage0_55[25]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[7],stage1_56[10],stage1_55[16],stage1_54[20]}
   );
   gpc615_5 gpc254 (
      {stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48]},
      {stage0_55[26]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[8],stage1_56[11],stage1_55[17],stage1_54[21]}
   );
   gpc615_5 gpc255 (
      {stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage0_55[27]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[9],stage1_56[12],stage1_55[18],stage1_54[22]}
   );
   gpc606_5 gpc256 (
      {stage0_55[28], stage0_55[29], stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[10],stage1_56[13],stage1_55[19]}
   );
   gpc606_5 gpc257 (
      {stage0_55[34], stage0_55[35], stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[11],stage1_56[14],stage1_55[20]}
   );
   gpc606_5 gpc258 (
      {stage0_55[40], stage0_55[41], stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[12],stage1_56[15],stage1_55[21]}
   );
   gpc606_5 gpc259 (
      {stage0_55[46], stage0_55[47], stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[13],stage1_56[16],stage1_55[22]}
   );
   gpc606_5 gpc260 (
      {stage0_55[52], stage0_55[53], stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[10],stage1_57[14],stage1_56[17],stage1_55[23]}
   );
   gpc606_5 gpc261 (
      {stage0_55[58], stage0_55[59], stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[11],stage1_57[15],stage1_56[18],stage1_55[24]}
   );
   gpc606_5 gpc262 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[6],stage1_58[12],stage1_57[16],stage1_56[19]}
   );
   gpc615_5 gpc263 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46]},
      {stage0_57[36]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[7],stage1_58[13],stage1_57[17],stage1_56[20]}
   );
   gpc615_5 gpc264 (
      {stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_57[37]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[8],stage1_58[14],stage1_57[18],stage1_56[21]}
   );
   gpc615_5 gpc265 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56]},
      {stage0_57[38]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[9],stage1_58[15],stage1_57[19],stage1_56[22]}
   );
   gpc615_5 gpc266 (
      {stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_57[39]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[10],stage1_58[16],stage1_57[20],stage1_56[23]}
   );
   gpc615_5 gpc267 (
      {stage0_57[40], stage0_57[41], stage0_57[42], stage0_57[43], stage0_57[44]},
      {stage0_58[30]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[5],stage1_59[11],stage1_58[17],stage1_57[21]}
   );
   gpc615_5 gpc268 (
      {stage0_57[45], stage0_57[46], stage0_57[47], stage0_57[48], stage0_57[49]},
      {stage0_58[31]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[6],stage1_59[12],stage1_58[18],stage1_57[22]}
   );
   gpc615_5 gpc269 (
      {stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53], stage0_57[54]},
      {stage0_58[32]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[7],stage1_59[13],stage1_58[19],stage1_57[23]}
   );
   gpc615_5 gpc270 (
      {stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_58[33]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[8],stage1_59[14],stage1_58[20],stage1_57[24]}
   );
   gpc615_5 gpc271 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], 1'b0},
      {stage0_58[34]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[9],stage1_59[15],stage1_58[21],stage1_57[25]}
   );
   gpc1406_5 gpc272 (
      {stage0_58[35], stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3]},
      {stage0_61[0]},
      {stage1_62[0],stage1_61[5],stage1_60[10],stage1_59[16],stage1_58[22]}
   );
   gpc606_5 gpc273 (
      {stage0_58[41], stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46]},
      {stage0_60[4], stage0_60[5], stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9]},
      {stage1_62[1],stage1_61[6],stage1_60[11],stage1_59[17],stage1_58[23]}
   );
   gpc606_5 gpc274 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5], stage0_61[6]},
      {stage1_63[0],stage1_62[2],stage1_61[7],stage1_60[12],stage1_59[18]}
   );
   gpc606_5 gpc275 (
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11], stage0_61[12]},
      {stage1_63[1],stage1_62[3],stage1_61[8],stage1_60[13],stage1_59[19]}
   );
   gpc606_5 gpc276 (
      {stage0_60[10], stage0_60[11], stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[2],stage1_62[4],stage1_61[9],stage1_60[14]}
   );
   gpc606_5 gpc277 (
      {stage0_60[16], stage0_60[17], stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[3],stage1_62[5],stage1_61[10],stage1_60[15]}
   );
   gpc606_5 gpc278 (
      {stage0_60[22], stage0_60[23], stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[4],stage1_62[6],stage1_61[11],stage1_60[16]}
   );
   gpc606_5 gpc279 (
      {stage0_60[28], stage0_60[29], stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[5],stage1_62[7],stage1_61[12],stage1_60[17]}
   );
   gpc606_5 gpc280 (
      {stage0_60[34], stage0_60[35], stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[6],stage1_62[8],stage1_61[13],stage1_60[18]}
   );
   gpc606_5 gpc281 (
      {stage0_60[40], stage0_60[41], stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[7],stage1_62[9],stage1_61[14],stage1_60[19]}
   );
   gpc606_5 gpc282 (
      {stage0_60[46], stage0_60[47], stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[8],stage1_62[10],stage1_61[15],stage1_60[20]}
   );
   gpc615_5 gpc283 (
      {stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_62[42]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[7],stage1_63[9],stage1_62[11],stage1_61[16]}
   );
   gpc615_5 gpc284 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22]},
      {stage0_62[43]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[8],stage1_63[10],stage1_62[12],stage1_61[17]}
   );
   gpc615_5 gpc285 (
      {stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27]},
      {stage0_62[44]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[9],stage1_63[11],stage1_62[13],stage1_61[18]}
   );
   gpc615_5 gpc286 (
      {stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage0_62[45]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[10],stage1_63[12],stage1_62[14],stage1_61[19]}
   );
   gpc615_5 gpc287 (
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37]},
      {stage0_62[46]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[11],stage1_63[13],stage1_62[15],stage1_61[20]}
   );
   gpc615_5 gpc288 (
      {stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42]},
      {stage0_62[47]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[12],stage1_63[14],stage1_62[16],stage1_61[21]}
   );
   gpc615_5 gpc289 (
      {stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_62[48]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[13],stage1_63[15],stage1_62[17],stage1_61[22]}
   );
   gpc615_5 gpc290 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52]},
      {stage0_62[49]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[14],stage1_63[16],stage1_62[18],stage1_61[23]}
   );
   gpc615_5 gpc291 (
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57]},
      {stage0_62[50]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[15],stage1_63[17],stage1_62[19],stage1_61[24]}
   );
   gpc1_1 gpc292 (
      {stage0_0[54]},
      {stage1_0[9]}
   );
   gpc1_1 gpc293 (
      {stage0_0[55]},
      {stage1_0[10]}
   );
   gpc1_1 gpc294 (
      {stage0_0[56]},
      {stage1_0[11]}
   );
   gpc1_1 gpc295 (
      {stage0_0[57]},
      {stage1_0[12]}
   );
   gpc1_1 gpc296 (
      {stage0_0[58]},
      {stage1_0[13]}
   );
   gpc1_1 gpc297 (
      {stage0_0[59]},
      {stage1_0[14]}
   );
   gpc1_1 gpc298 (
      {stage0_0[60]},
      {stage1_0[15]}
   );
   gpc1_1 gpc299 (
      {stage0_0[61]},
      {stage1_0[16]}
   );
   gpc1_1 gpc300 (
      {stage0_0[62]},
      {stage1_0[17]}
   );
   gpc1_1 gpc301 (
      {stage0_0[63]},
      {stage1_0[18]}
   );
   gpc1_1 gpc302 (
      {stage0_1[30]},
      {stage1_1[14]}
   );
   gpc1_1 gpc303 (
      {stage0_1[31]},
      {stage1_1[15]}
   );
   gpc1_1 gpc304 (
      {stage0_1[32]},
      {stage1_1[16]}
   );
   gpc1_1 gpc305 (
      {stage0_1[33]},
      {stage1_1[17]}
   );
   gpc1_1 gpc306 (
      {stage0_1[34]},
      {stage1_1[18]}
   );
   gpc1_1 gpc307 (
      {stage0_1[35]},
      {stage1_1[19]}
   );
   gpc1_1 gpc308 (
      {stage0_1[36]},
      {stage1_1[20]}
   );
   gpc1_1 gpc309 (
      {stage0_1[37]},
      {stage1_1[21]}
   );
   gpc1_1 gpc310 (
      {stage0_1[38]},
      {stage1_1[22]}
   );
   gpc1_1 gpc311 (
      {stage0_1[39]},
      {stage1_1[23]}
   );
   gpc1_1 gpc312 (
      {stage0_1[40]},
      {stage1_1[24]}
   );
   gpc1_1 gpc313 (
      {stage0_1[41]},
      {stage1_1[25]}
   );
   gpc1_1 gpc314 (
      {stage0_1[42]},
      {stage1_1[26]}
   );
   gpc1_1 gpc315 (
      {stage0_1[43]},
      {stage1_1[27]}
   );
   gpc1_1 gpc316 (
      {stage0_1[44]},
      {stage1_1[28]}
   );
   gpc1_1 gpc317 (
      {stage0_1[45]},
      {stage1_1[29]}
   );
   gpc1_1 gpc318 (
      {stage0_1[46]},
      {stage1_1[30]}
   );
   gpc1_1 gpc319 (
      {stage0_1[47]},
      {stage1_1[31]}
   );
   gpc1_1 gpc320 (
      {stage0_1[48]},
      {stage1_1[32]}
   );
   gpc1_1 gpc321 (
      {stage0_1[49]},
      {stage1_1[33]}
   );
   gpc1_1 gpc322 (
      {stage0_1[50]},
      {stage1_1[34]}
   );
   gpc1_1 gpc323 (
      {stage0_1[51]},
      {stage1_1[35]}
   );
   gpc1_1 gpc324 (
      {stage0_1[52]},
      {stage1_1[36]}
   );
   gpc1_1 gpc325 (
      {stage0_1[53]},
      {stage1_1[37]}
   );
   gpc1_1 gpc326 (
      {stage0_1[54]},
      {stage1_1[38]}
   );
   gpc1_1 gpc327 (
      {stage0_1[55]},
      {stage1_1[39]}
   );
   gpc1_1 gpc328 (
      {stage0_1[56]},
      {stage1_1[40]}
   );
   gpc1_1 gpc329 (
      {stage0_1[57]},
      {stage1_1[41]}
   );
   gpc1_1 gpc330 (
      {stage0_1[58]},
      {stage1_1[42]}
   );
   gpc1_1 gpc331 (
      {stage0_1[59]},
      {stage1_1[43]}
   );
   gpc1_1 gpc332 (
      {stage0_1[60]},
      {stage1_1[44]}
   );
   gpc1_1 gpc333 (
      {stage0_1[61]},
      {stage1_1[45]}
   );
   gpc1_1 gpc334 (
      {stage0_1[62]},
      {stage1_1[46]}
   );
   gpc1_1 gpc335 (
      {stage0_1[63]},
      {stage1_1[47]}
   );
   gpc1_1 gpc336 (
      {stage0_2[54]},
      {stage1_2[14]}
   );
   gpc1_1 gpc337 (
      {stage0_2[55]},
      {stage1_2[15]}
   );
   gpc1_1 gpc338 (
      {stage0_2[56]},
      {stage1_2[16]}
   );
   gpc1_1 gpc339 (
      {stage0_2[57]},
      {stage1_2[17]}
   );
   gpc1_1 gpc340 (
      {stage0_2[58]},
      {stage1_2[18]}
   );
   gpc1_1 gpc341 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc342 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc343 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc344 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc345 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc346 (
      {stage0_3[55]},
      {stage1_3[19]}
   );
   gpc1_1 gpc347 (
      {stage0_3[56]},
      {stage1_3[20]}
   );
   gpc1_1 gpc348 (
      {stage0_3[57]},
      {stage1_3[21]}
   );
   gpc1_1 gpc349 (
      {stage0_3[58]},
      {stage1_3[22]}
   );
   gpc1_1 gpc350 (
      {stage0_3[59]},
      {stage1_3[23]}
   );
   gpc1_1 gpc351 (
      {stage0_3[60]},
      {stage1_3[24]}
   );
   gpc1_1 gpc352 (
      {stage0_3[61]},
      {stage1_3[25]}
   );
   gpc1_1 gpc353 (
      {stage0_3[62]},
      {stage1_3[26]}
   );
   gpc1_1 gpc354 (
      {stage0_3[63]},
      {stage1_3[27]}
   );
   gpc1_1 gpc355 (
      {stage0_4[53]},
      {stage1_4[27]}
   );
   gpc1_1 gpc356 (
      {stage0_4[54]},
      {stage1_4[28]}
   );
   gpc1_1 gpc357 (
      {stage0_4[55]},
      {stage1_4[29]}
   );
   gpc1_1 gpc358 (
      {stage0_4[56]},
      {stage1_4[30]}
   );
   gpc1_1 gpc359 (
      {stage0_4[57]},
      {stage1_4[31]}
   );
   gpc1_1 gpc360 (
      {stage0_4[58]},
      {stage1_4[32]}
   );
   gpc1_1 gpc361 (
      {stage0_4[59]},
      {stage1_4[33]}
   );
   gpc1_1 gpc362 (
      {stage0_4[60]},
      {stage1_4[34]}
   );
   gpc1_1 gpc363 (
      {stage0_4[61]},
      {stage1_4[35]}
   );
   gpc1_1 gpc364 (
      {stage0_4[62]},
      {stage1_4[36]}
   );
   gpc1_1 gpc365 (
      {stage0_4[63]},
      {stage1_4[37]}
   );
   gpc1_1 gpc366 (
      {stage0_5[60]},
      {stage1_5[23]}
   );
   gpc1_1 gpc367 (
      {stage0_5[61]},
      {stage1_5[24]}
   );
   gpc1_1 gpc368 (
      {stage0_5[62]},
      {stage1_5[25]}
   );
   gpc1_1 gpc369 (
      {stage0_5[63]},
      {stage1_5[26]}
   );
   gpc1_1 gpc370 (
      {stage0_6[63]},
      {stage1_6[21]}
   );
   gpc1_1 gpc371 (
      {stage0_7[53]},
      {stage1_7[25]}
   );
   gpc1_1 gpc372 (
      {stage0_7[54]},
      {stage1_7[26]}
   );
   gpc1_1 gpc373 (
      {stage0_7[55]},
      {stage1_7[27]}
   );
   gpc1_1 gpc374 (
      {stage0_7[56]},
      {stage1_7[28]}
   );
   gpc1_1 gpc375 (
      {stage0_7[57]},
      {stage1_7[29]}
   );
   gpc1_1 gpc376 (
      {stage0_7[58]},
      {stage1_7[30]}
   );
   gpc1_1 gpc377 (
      {stage0_7[59]},
      {stage1_7[31]}
   );
   gpc1_1 gpc378 (
      {stage0_7[60]},
      {stage1_7[32]}
   );
   gpc1_1 gpc379 (
      {stage0_7[61]},
      {stage1_7[33]}
   );
   gpc1_1 gpc380 (
      {stage0_7[62]},
      {stage1_7[34]}
   );
   gpc1_1 gpc381 (
      {stage0_7[63]},
      {stage1_7[35]}
   );
   gpc1_1 gpc382 (
      {stage0_9[60]},
      {stage1_9[25]}
   );
   gpc1_1 gpc383 (
      {stage0_9[61]},
      {stage1_9[26]}
   );
   gpc1_1 gpc384 (
      {stage0_9[62]},
      {stage1_9[27]}
   );
   gpc1_1 gpc385 (
      {stage0_9[63]},
      {stage1_9[28]}
   );
   gpc1_1 gpc386 (
      {stage0_10[52]},
      {stage1_10[22]}
   );
   gpc1_1 gpc387 (
      {stage0_10[53]},
      {stage1_10[23]}
   );
   gpc1_1 gpc388 (
      {stage0_10[54]},
      {stage1_10[24]}
   );
   gpc1_1 gpc389 (
      {stage0_10[55]},
      {stage1_10[25]}
   );
   gpc1_1 gpc390 (
      {stage0_10[56]},
      {stage1_10[26]}
   );
   gpc1_1 gpc391 (
      {stage0_10[57]},
      {stage1_10[27]}
   );
   gpc1_1 gpc392 (
      {stage0_10[58]},
      {stage1_10[28]}
   );
   gpc1_1 gpc393 (
      {stage0_10[59]},
      {stage1_10[29]}
   );
   gpc1_1 gpc394 (
      {stage0_10[60]},
      {stage1_10[30]}
   );
   gpc1_1 gpc395 (
      {stage0_10[61]},
      {stage1_10[31]}
   );
   gpc1_1 gpc396 (
      {stage0_10[62]},
      {stage1_10[32]}
   );
   gpc1_1 gpc397 (
      {stage0_10[63]},
      {stage1_10[33]}
   );
   gpc1_1 gpc398 (
      {stage0_11[53]},
      {stage1_11[22]}
   );
   gpc1_1 gpc399 (
      {stage0_11[54]},
      {stage1_11[23]}
   );
   gpc1_1 gpc400 (
      {stage0_11[55]},
      {stage1_11[24]}
   );
   gpc1_1 gpc401 (
      {stage0_11[56]},
      {stage1_11[25]}
   );
   gpc1_1 gpc402 (
      {stage0_11[57]},
      {stage1_11[26]}
   );
   gpc1_1 gpc403 (
      {stage0_11[58]},
      {stage1_11[27]}
   );
   gpc1_1 gpc404 (
      {stage0_11[59]},
      {stage1_11[28]}
   );
   gpc1_1 gpc405 (
      {stage0_11[60]},
      {stage1_11[29]}
   );
   gpc1_1 gpc406 (
      {stage0_11[61]},
      {stage1_11[30]}
   );
   gpc1_1 gpc407 (
      {stage0_11[62]},
      {stage1_11[31]}
   );
   gpc1_1 gpc408 (
      {stage0_11[63]},
      {stage1_11[32]}
   );
   gpc1_1 gpc409 (
      {stage0_12[63]},
      {stage1_12[26]}
   );
   gpc1_1 gpc410 (
      {stage0_13[59]},
      {stage1_13[26]}
   );
   gpc1_1 gpc411 (
      {stage0_13[60]},
      {stage1_13[27]}
   );
   gpc1_1 gpc412 (
      {stage0_13[61]},
      {stage1_13[28]}
   );
   gpc1_1 gpc413 (
      {stage0_13[62]},
      {stage1_13[29]}
   );
   gpc1_1 gpc414 (
      {stage0_13[63]},
      {stage1_13[30]}
   );
   gpc1_1 gpc415 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc416 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc417 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc418 (
      {stage0_15[39]},
      {stage1_15[20]}
   );
   gpc1_1 gpc419 (
      {stage0_15[40]},
      {stage1_15[21]}
   );
   gpc1_1 gpc420 (
      {stage0_15[41]},
      {stage1_15[22]}
   );
   gpc1_1 gpc421 (
      {stage0_15[42]},
      {stage1_15[23]}
   );
   gpc1_1 gpc422 (
      {stage0_15[43]},
      {stage1_15[24]}
   );
   gpc1_1 gpc423 (
      {stage0_15[44]},
      {stage1_15[25]}
   );
   gpc1_1 gpc424 (
      {stage0_15[45]},
      {stage1_15[26]}
   );
   gpc1_1 gpc425 (
      {stage0_15[46]},
      {stage1_15[27]}
   );
   gpc1_1 gpc426 (
      {stage0_15[47]},
      {stage1_15[28]}
   );
   gpc1_1 gpc427 (
      {stage0_15[48]},
      {stage1_15[29]}
   );
   gpc1_1 gpc428 (
      {stage0_15[49]},
      {stage1_15[30]}
   );
   gpc1_1 gpc429 (
      {stage0_15[50]},
      {stage1_15[31]}
   );
   gpc1_1 gpc430 (
      {stage0_15[51]},
      {stage1_15[32]}
   );
   gpc1_1 gpc431 (
      {stage0_15[52]},
      {stage1_15[33]}
   );
   gpc1_1 gpc432 (
      {stage0_15[53]},
      {stage1_15[34]}
   );
   gpc1_1 gpc433 (
      {stage0_15[54]},
      {stage1_15[35]}
   );
   gpc1_1 gpc434 (
      {stage0_15[55]},
      {stage1_15[36]}
   );
   gpc1_1 gpc435 (
      {stage0_15[56]},
      {stage1_15[37]}
   );
   gpc1_1 gpc436 (
      {stage0_15[57]},
      {stage1_15[38]}
   );
   gpc1_1 gpc437 (
      {stage0_15[58]},
      {stage1_15[39]}
   );
   gpc1_1 gpc438 (
      {stage0_15[59]},
      {stage1_15[40]}
   );
   gpc1_1 gpc439 (
      {stage0_15[60]},
      {stage1_15[41]}
   );
   gpc1_1 gpc440 (
      {stage0_15[61]},
      {stage1_15[42]}
   );
   gpc1_1 gpc441 (
      {stage0_15[62]},
      {stage1_15[43]}
   );
   gpc1_1 gpc442 (
      {stage0_15[63]},
      {stage1_15[44]}
   );
   gpc1_1 gpc443 (
      {stage0_16[58]},
      {stage1_16[25]}
   );
   gpc1_1 gpc444 (
      {stage0_16[59]},
      {stage1_16[26]}
   );
   gpc1_1 gpc445 (
      {stage0_16[60]},
      {stage1_16[27]}
   );
   gpc1_1 gpc446 (
      {stage0_16[61]},
      {stage1_16[28]}
   );
   gpc1_1 gpc447 (
      {stage0_16[62]},
      {stage1_16[29]}
   );
   gpc1_1 gpc448 (
      {stage0_16[63]},
      {stage1_16[30]}
   );
   gpc1_1 gpc449 (
      {stage0_17[43]},
      {stage1_17[24]}
   );
   gpc1_1 gpc450 (
      {stage0_17[44]},
      {stage1_17[25]}
   );
   gpc1_1 gpc451 (
      {stage0_17[45]},
      {stage1_17[26]}
   );
   gpc1_1 gpc452 (
      {stage0_17[46]},
      {stage1_17[27]}
   );
   gpc1_1 gpc453 (
      {stage0_17[47]},
      {stage1_17[28]}
   );
   gpc1_1 gpc454 (
      {stage0_17[48]},
      {stage1_17[29]}
   );
   gpc1_1 gpc455 (
      {stage0_17[49]},
      {stage1_17[30]}
   );
   gpc1_1 gpc456 (
      {stage0_17[50]},
      {stage1_17[31]}
   );
   gpc1_1 gpc457 (
      {stage0_17[51]},
      {stage1_17[32]}
   );
   gpc1_1 gpc458 (
      {stage0_17[52]},
      {stage1_17[33]}
   );
   gpc1_1 gpc459 (
      {stage0_17[53]},
      {stage1_17[34]}
   );
   gpc1_1 gpc460 (
      {stage0_17[54]},
      {stage1_17[35]}
   );
   gpc1_1 gpc461 (
      {stage0_17[55]},
      {stage1_17[36]}
   );
   gpc1_1 gpc462 (
      {stage0_17[56]},
      {stage1_17[37]}
   );
   gpc1_1 gpc463 (
      {stage0_17[57]},
      {stage1_17[38]}
   );
   gpc1_1 gpc464 (
      {stage0_17[58]},
      {stage1_17[39]}
   );
   gpc1_1 gpc465 (
      {stage0_17[59]},
      {stage1_17[40]}
   );
   gpc1_1 gpc466 (
      {stage0_17[60]},
      {stage1_17[41]}
   );
   gpc1_1 gpc467 (
      {stage0_17[61]},
      {stage1_17[42]}
   );
   gpc1_1 gpc468 (
      {stage0_17[62]},
      {stage1_17[43]}
   );
   gpc1_1 gpc469 (
      {stage0_17[63]},
      {stage1_17[44]}
   );
   gpc1_1 gpc470 (
      {stage0_18[60]},
      {stage1_18[19]}
   );
   gpc1_1 gpc471 (
      {stage0_18[61]},
      {stage1_18[20]}
   );
   gpc1_1 gpc472 (
      {stage0_18[62]},
      {stage1_18[21]}
   );
   gpc1_1 gpc473 (
      {stage0_18[63]},
      {stage1_18[22]}
   );
   gpc1_1 gpc474 (
      {stage0_19[54]},
      {stage1_19[19]}
   );
   gpc1_1 gpc475 (
      {stage0_19[55]},
      {stage1_19[20]}
   );
   gpc1_1 gpc476 (
      {stage0_19[56]},
      {stage1_19[21]}
   );
   gpc1_1 gpc477 (
      {stage0_19[57]},
      {stage1_19[22]}
   );
   gpc1_1 gpc478 (
      {stage0_19[58]},
      {stage1_19[23]}
   );
   gpc1_1 gpc479 (
      {stage0_19[59]},
      {stage1_19[24]}
   );
   gpc1_1 gpc480 (
      {stage0_19[60]},
      {stage1_19[25]}
   );
   gpc1_1 gpc481 (
      {stage0_19[61]},
      {stage1_19[26]}
   );
   gpc1_1 gpc482 (
      {stage0_19[62]},
      {stage1_19[27]}
   );
   gpc1_1 gpc483 (
      {stage0_19[63]},
      {stage1_19[28]}
   );
   gpc1_1 gpc484 (
      {stage0_20[49]},
      {stage1_20[26]}
   );
   gpc1_1 gpc485 (
      {stage0_20[50]},
      {stage1_20[27]}
   );
   gpc1_1 gpc486 (
      {stage0_20[51]},
      {stage1_20[28]}
   );
   gpc1_1 gpc487 (
      {stage0_20[52]},
      {stage1_20[29]}
   );
   gpc1_1 gpc488 (
      {stage0_20[53]},
      {stage1_20[30]}
   );
   gpc1_1 gpc489 (
      {stage0_20[54]},
      {stage1_20[31]}
   );
   gpc1_1 gpc490 (
      {stage0_20[55]},
      {stage1_20[32]}
   );
   gpc1_1 gpc491 (
      {stage0_20[56]},
      {stage1_20[33]}
   );
   gpc1_1 gpc492 (
      {stage0_20[57]},
      {stage1_20[34]}
   );
   gpc1_1 gpc493 (
      {stage0_20[58]},
      {stage1_20[35]}
   );
   gpc1_1 gpc494 (
      {stage0_20[59]},
      {stage1_20[36]}
   );
   gpc1_1 gpc495 (
      {stage0_20[60]},
      {stage1_20[37]}
   );
   gpc1_1 gpc496 (
      {stage0_20[61]},
      {stage1_20[38]}
   );
   gpc1_1 gpc497 (
      {stage0_20[62]},
      {stage1_20[39]}
   );
   gpc1_1 gpc498 (
      {stage0_20[63]},
      {stage1_20[40]}
   );
   gpc1_1 gpc499 (
      {stage0_21[55]},
      {stage1_21[24]}
   );
   gpc1_1 gpc500 (
      {stage0_21[56]},
      {stage1_21[25]}
   );
   gpc1_1 gpc501 (
      {stage0_21[57]},
      {stage1_21[26]}
   );
   gpc1_1 gpc502 (
      {stage0_21[58]},
      {stage1_21[27]}
   );
   gpc1_1 gpc503 (
      {stage0_21[59]},
      {stage1_21[28]}
   );
   gpc1_1 gpc504 (
      {stage0_21[60]},
      {stage1_21[29]}
   );
   gpc1_1 gpc505 (
      {stage0_21[61]},
      {stage1_21[30]}
   );
   gpc1_1 gpc506 (
      {stage0_21[62]},
      {stage1_21[31]}
   );
   gpc1_1 gpc507 (
      {stage0_21[63]},
      {stage1_21[32]}
   );
   gpc1_1 gpc508 (
      {stage0_22[52]},
      {stage1_22[19]}
   );
   gpc1_1 gpc509 (
      {stage0_22[53]},
      {stage1_22[20]}
   );
   gpc1_1 gpc510 (
      {stage0_22[54]},
      {stage1_22[21]}
   );
   gpc1_1 gpc511 (
      {stage0_22[55]},
      {stage1_22[22]}
   );
   gpc1_1 gpc512 (
      {stage0_22[56]},
      {stage1_22[23]}
   );
   gpc1_1 gpc513 (
      {stage0_22[57]},
      {stage1_22[24]}
   );
   gpc1_1 gpc514 (
      {stage0_22[58]},
      {stage1_22[25]}
   );
   gpc1_1 gpc515 (
      {stage0_22[59]},
      {stage1_22[26]}
   );
   gpc1_1 gpc516 (
      {stage0_22[60]},
      {stage1_22[27]}
   );
   gpc1_1 gpc517 (
      {stage0_22[61]},
      {stage1_22[28]}
   );
   gpc1_1 gpc518 (
      {stage0_22[62]},
      {stage1_22[29]}
   );
   gpc1_1 gpc519 (
      {stage0_22[63]},
      {stage1_22[30]}
   );
   gpc1_1 gpc520 (
      {stage0_23[48]},
      {stage1_23[19]}
   );
   gpc1_1 gpc521 (
      {stage0_23[49]},
      {stage1_23[20]}
   );
   gpc1_1 gpc522 (
      {stage0_23[50]},
      {stage1_23[21]}
   );
   gpc1_1 gpc523 (
      {stage0_23[51]},
      {stage1_23[22]}
   );
   gpc1_1 gpc524 (
      {stage0_23[52]},
      {stage1_23[23]}
   );
   gpc1_1 gpc525 (
      {stage0_23[53]},
      {stage1_23[24]}
   );
   gpc1_1 gpc526 (
      {stage0_23[54]},
      {stage1_23[25]}
   );
   gpc1_1 gpc527 (
      {stage0_23[55]},
      {stage1_23[26]}
   );
   gpc1_1 gpc528 (
      {stage0_23[56]},
      {stage1_23[27]}
   );
   gpc1_1 gpc529 (
      {stage0_23[57]},
      {stage1_23[28]}
   );
   gpc1_1 gpc530 (
      {stage0_23[58]},
      {stage1_23[29]}
   );
   gpc1_1 gpc531 (
      {stage0_23[59]},
      {stage1_23[30]}
   );
   gpc1_1 gpc532 (
      {stage0_23[60]},
      {stage1_23[31]}
   );
   gpc1_1 gpc533 (
      {stage0_23[61]},
      {stage1_23[32]}
   );
   gpc1_1 gpc534 (
      {stage0_23[62]},
      {stage1_23[33]}
   );
   gpc1_1 gpc535 (
      {stage0_23[63]},
      {stage1_23[34]}
   );
   gpc1_1 gpc536 (
      {stage0_24[62]},
      {stage1_24[25]}
   );
   gpc1_1 gpc537 (
      {stage0_24[63]},
      {stage1_24[26]}
   );
   gpc1_1 gpc538 (
      {stage0_25[42]},
      {stage1_25[23]}
   );
   gpc1_1 gpc539 (
      {stage0_25[43]},
      {stage1_25[24]}
   );
   gpc1_1 gpc540 (
      {stage0_25[44]},
      {stage1_25[25]}
   );
   gpc1_1 gpc541 (
      {stage0_25[45]},
      {stage1_25[26]}
   );
   gpc1_1 gpc542 (
      {stage0_25[46]},
      {stage1_25[27]}
   );
   gpc1_1 gpc543 (
      {stage0_25[47]},
      {stage1_25[28]}
   );
   gpc1_1 gpc544 (
      {stage0_25[48]},
      {stage1_25[29]}
   );
   gpc1_1 gpc545 (
      {stage0_25[49]},
      {stage1_25[30]}
   );
   gpc1_1 gpc546 (
      {stage0_25[50]},
      {stage1_25[31]}
   );
   gpc1_1 gpc547 (
      {stage0_25[51]},
      {stage1_25[32]}
   );
   gpc1_1 gpc548 (
      {stage0_25[52]},
      {stage1_25[33]}
   );
   gpc1_1 gpc549 (
      {stage0_25[53]},
      {stage1_25[34]}
   );
   gpc1_1 gpc550 (
      {stage0_25[54]},
      {stage1_25[35]}
   );
   gpc1_1 gpc551 (
      {stage0_25[55]},
      {stage1_25[36]}
   );
   gpc1_1 gpc552 (
      {stage0_25[56]},
      {stage1_25[37]}
   );
   gpc1_1 gpc553 (
      {stage0_25[57]},
      {stage1_25[38]}
   );
   gpc1_1 gpc554 (
      {stage0_25[58]},
      {stage1_25[39]}
   );
   gpc1_1 gpc555 (
      {stage0_25[59]},
      {stage1_25[40]}
   );
   gpc1_1 gpc556 (
      {stage0_25[60]},
      {stage1_25[41]}
   );
   gpc1_1 gpc557 (
      {stage0_25[61]},
      {stage1_25[42]}
   );
   gpc1_1 gpc558 (
      {stage0_25[62]},
      {stage1_25[43]}
   );
   gpc1_1 gpc559 (
      {stage0_25[63]},
      {stage1_25[44]}
   );
   gpc1_1 gpc560 (
      {stage0_26[53]},
      {stage1_26[18]}
   );
   gpc1_1 gpc561 (
      {stage0_26[54]},
      {stage1_26[19]}
   );
   gpc1_1 gpc562 (
      {stage0_26[55]},
      {stage1_26[20]}
   );
   gpc1_1 gpc563 (
      {stage0_26[56]},
      {stage1_26[21]}
   );
   gpc1_1 gpc564 (
      {stage0_26[57]},
      {stage1_26[22]}
   );
   gpc1_1 gpc565 (
      {stage0_26[58]},
      {stage1_26[23]}
   );
   gpc1_1 gpc566 (
      {stage0_26[59]},
      {stage1_26[24]}
   );
   gpc1_1 gpc567 (
      {stage0_26[60]},
      {stage1_26[25]}
   );
   gpc1_1 gpc568 (
      {stage0_26[61]},
      {stage1_26[26]}
   );
   gpc1_1 gpc569 (
      {stage0_26[62]},
      {stage1_26[27]}
   );
   gpc1_1 gpc570 (
      {stage0_26[63]},
      {stage1_26[28]}
   );
   gpc1_1 gpc571 (
      {stage0_27[41]},
      {stage1_27[18]}
   );
   gpc1_1 gpc572 (
      {stage0_27[42]},
      {stage1_27[19]}
   );
   gpc1_1 gpc573 (
      {stage0_27[43]},
      {stage1_27[20]}
   );
   gpc1_1 gpc574 (
      {stage0_27[44]},
      {stage1_27[21]}
   );
   gpc1_1 gpc575 (
      {stage0_27[45]},
      {stage1_27[22]}
   );
   gpc1_1 gpc576 (
      {stage0_27[46]},
      {stage1_27[23]}
   );
   gpc1_1 gpc577 (
      {stage0_27[47]},
      {stage1_27[24]}
   );
   gpc1_1 gpc578 (
      {stage0_27[48]},
      {stage1_27[25]}
   );
   gpc1_1 gpc579 (
      {stage0_27[49]},
      {stage1_27[26]}
   );
   gpc1_1 gpc580 (
      {stage0_27[50]},
      {stage1_27[27]}
   );
   gpc1_1 gpc581 (
      {stage0_27[51]},
      {stage1_27[28]}
   );
   gpc1_1 gpc582 (
      {stage0_27[52]},
      {stage1_27[29]}
   );
   gpc1_1 gpc583 (
      {stage0_27[53]},
      {stage1_27[30]}
   );
   gpc1_1 gpc584 (
      {stage0_27[54]},
      {stage1_27[31]}
   );
   gpc1_1 gpc585 (
      {stage0_27[55]},
      {stage1_27[32]}
   );
   gpc1_1 gpc586 (
      {stage0_27[56]},
      {stage1_27[33]}
   );
   gpc1_1 gpc587 (
      {stage0_27[57]},
      {stage1_27[34]}
   );
   gpc1_1 gpc588 (
      {stage0_27[58]},
      {stage1_27[35]}
   );
   gpc1_1 gpc589 (
      {stage0_27[59]},
      {stage1_27[36]}
   );
   gpc1_1 gpc590 (
      {stage0_27[60]},
      {stage1_27[37]}
   );
   gpc1_1 gpc591 (
      {stage0_27[61]},
      {stage1_27[38]}
   );
   gpc1_1 gpc592 (
      {stage0_27[62]},
      {stage1_27[39]}
   );
   gpc1_1 gpc593 (
      {stage0_27[63]},
      {stage1_27[40]}
   );
   gpc1_1 gpc594 (
      {stage0_28[62]},
      {stage1_28[25]}
   );
   gpc1_1 gpc595 (
      {stage0_28[63]},
      {stage1_28[26]}
   );
   gpc1_1 gpc596 (
      {stage0_29[60]},
      {stage1_29[25]}
   );
   gpc1_1 gpc597 (
      {stage0_29[61]},
      {stage1_29[26]}
   );
   gpc1_1 gpc598 (
      {stage0_29[62]},
      {stage1_29[27]}
   );
   gpc1_1 gpc599 (
      {stage0_29[63]},
      {stage1_29[28]}
   );
   gpc1_1 gpc600 (
      {stage0_30[59]},
      {stage1_30[21]}
   );
   gpc1_1 gpc601 (
      {stage0_30[60]},
      {stage1_30[22]}
   );
   gpc1_1 gpc602 (
      {stage0_30[61]},
      {stage1_30[23]}
   );
   gpc1_1 gpc603 (
      {stage0_30[62]},
      {stage1_30[24]}
   );
   gpc1_1 gpc604 (
      {stage0_30[63]},
      {stage1_30[25]}
   );
   gpc1_1 gpc605 (
      {stage0_32[63]},
      {stage1_32[30]}
   );
   gpc1_1 gpc606 (
      {stage0_33[53]},
      {stage1_33[27]}
   );
   gpc1_1 gpc607 (
      {stage0_33[54]},
      {stage1_33[28]}
   );
   gpc1_1 gpc608 (
      {stage0_33[55]},
      {stage1_33[29]}
   );
   gpc1_1 gpc609 (
      {stage0_33[56]},
      {stage1_33[30]}
   );
   gpc1_1 gpc610 (
      {stage0_33[57]},
      {stage1_33[31]}
   );
   gpc1_1 gpc611 (
      {stage0_33[58]},
      {stage1_33[32]}
   );
   gpc1_1 gpc612 (
      {stage0_33[59]},
      {stage1_33[33]}
   );
   gpc1_1 gpc613 (
      {stage0_33[60]},
      {stage1_33[34]}
   );
   gpc1_1 gpc614 (
      {stage0_33[61]},
      {stage1_33[35]}
   );
   gpc1_1 gpc615 (
      {stage0_33[62]},
      {stage1_33[36]}
   );
   gpc1_1 gpc616 (
      {stage0_33[63]},
      {stage1_33[37]}
   );
   gpc1_1 gpc617 (
      {stage0_34[60]},
      {stage1_34[20]}
   );
   gpc1_1 gpc618 (
      {stage0_34[61]},
      {stage1_34[21]}
   );
   gpc1_1 gpc619 (
      {stage0_34[62]},
      {stage1_34[22]}
   );
   gpc1_1 gpc620 (
      {stage0_34[63]},
      {stage1_34[23]}
   );
   gpc1_1 gpc621 (
      {stage0_35[57]},
      {stage1_35[23]}
   );
   gpc1_1 gpc622 (
      {stage0_35[58]},
      {stage1_35[24]}
   );
   gpc1_1 gpc623 (
      {stage0_35[59]},
      {stage1_35[25]}
   );
   gpc1_1 gpc624 (
      {stage0_35[60]},
      {stage1_35[26]}
   );
   gpc1_1 gpc625 (
      {stage0_35[61]},
      {stage1_35[27]}
   );
   gpc1_1 gpc626 (
      {stage0_35[62]},
      {stage1_35[28]}
   );
   gpc1_1 gpc627 (
      {stage0_35[63]},
      {stage1_35[29]}
   );
   gpc1_1 gpc628 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc629 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc630 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc631 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc632 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc633 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc634 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc635 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc636 (
      {stage0_36[54]},
      {stage1_36[34]}
   );
   gpc1_1 gpc637 (
      {stage0_36[55]},
      {stage1_36[35]}
   );
   gpc1_1 gpc638 (
      {stage0_36[56]},
      {stage1_36[36]}
   );
   gpc1_1 gpc639 (
      {stage0_36[57]},
      {stage1_36[37]}
   );
   gpc1_1 gpc640 (
      {stage0_36[58]},
      {stage1_36[38]}
   );
   gpc1_1 gpc641 (
      {stage0_36[59]},
      {stage1_36[39]}
   );
   gpc1_1 gpc642 (
      {stage0_36[60]},
      {stage1_36[40]}
   );
   gpc1_1 gpc643 (
      {stage0_36[61]},
      {stage1_36[41]}
   );
   gpc1_1 gpc644 (
      {stage0_36[62]},
      {stage1_36[42]}
   );
   gpc1_1 gpc645 (
      {stage0_36[63]},
      {stage1_36[43]}
   );
   gpc1_1 gpc646 (
      {stage0_38[41]},
      {stage1_38[19]}
   );
   gpc1_1 gpc647 (
      {stage0_38[42]},
      {stage1_38[20]}
   );
   gpc1_1 gpc648 (
      {stage0_38[43]},
      {stage1_38[21]}
   );
   gpc1_1 gpc649 (
      {stage0_38[44]},
      {stage1_38[22]}
   );
   gpc1_1 gpc650 (
      {stage0_38[45]},
      {stage1_38[23]}
   );
   gpc1_1 gpc651 (
      {stage0_38[46]},
      {stage1_38[24]}
   );
   gpc1_1 gpc652 (
      {stage0_38[47]},
      {stage1_38[25]}
   );
   gpc1_1 gpc653 (
      {stage0_38[48]},
      {stage1_38[26]}
   );
   gpc1_1 gpc654 (
      {stage0_38[49]},
      {stage1_38[27]}
   );
   gpc1_1 gpc655 (
      {stage0_38[50]},
      {stage1_38[28]}
   );
   gpc1_1 gpc656 (
      {stage0_38[51]},
      {stage1_38[29]}
   );
   gpc1_1 gpc657 (
      {stage0_38[52]},
      {stage1_38[30]}
   );
   gpc1_1 gpc658 (
      {stage0_38[53]},
      {stage1_38[31]}
   );
   gpc1_1 gpc659 (
      {stage0_38[54]},
      {stage1_38[32]}
   );
   gpc1_1 gpc660 (
      {stage0_38[55]},
      {stage1_38[33]}
   );
   gpc1_1 gpc661 (
      {stage0_38[56]},
      {stage1_38[34]}
   );
   gpc1_1 gpc662 (
      {stage0_38[57]},
      {stage1_38[35]}
   );
   gpc1_1 gpc663 (
      {stage0_38[58]},
      {stage1_38[36]}
   );
   gpc1_1 gpc664 (
      {stage0_38[59]},
      {stage1_38[37]}
   );
   gpc1_1 gpc665 (
      {stage0_38[60]},
      {stage1_38[38]}
   );
   gpc1_1 gpc666 (
      {stage0_38[61]},
      {stage1_38[39]}
   );
   gpc1_1 gpc667 (
      {stage0_38[62]},
      {stage1_38[40]}
   );
   gpc1_1 gpc668 (
      {stage0_38[63]},
      {stage1_38[41]}
   );
   gpc1_1 gpc669 (
      {stage0_39[63]},
      {stage1_39[22]}
   );
   gpc1_1 gpc670 (
      {stage0_41[54]},
      {stage1_41[26]}
   );
   gpc1_1 gpc671 (
      {stage0_41[55]},
      {stage1_41[27]}
   );
   gpc1_1 gpc672 (
      {stage0_41[56]},
      {stage1_41[28]}
   );
   gpc1_1 gpc673 (
      {stage0_41[57]},
      {stage1_41[29]}
   );
   gpc1_1 gpc674 (
      {stage0_41[58]},
      {stage1_41[30]}
   );
   gpc1_1 gpc675 (
      {stage0_41[59]},
      {stage1_41[31]}
   );
   gpc1_1 gpc676 (
      {stage0_41[60]},
      {stage1_41[32]}
   );
   gpc1_1 gpc677 (
      {stage0_41[61]},
      {stage1_41[33]}
   );
   gpc1_1 gpc678 (
      {stage0_41[62]},
      {stage1_41[34]}
   );
   gpc1_1 gpc679 (
      {stage0_41[63]},
      {stage1_41[35]}
   );
   gpc1_1 gpc680 (
      {stage0_42[54]},
      {stage1_42[19]}
   );
   gpc1_1 gpc681 (
      {stage0_42[55]},
      {stage1_42[20]}
   );
   gpc1_1 gpc682 (
      {stage0_42[56]},
      {stage1_42[21]}
   );
   gpc1_1 gpc683 (
      {stage0_42[57]},
      {stage1_42[22]}
   );
   gpc1_1 gpc684 (
      {stage0_42[58]},
      {stage1_42[23]}
   );
   gpc1_1 gpc685 (
      {stage0_42[59]},
      {stage1_42[24]}
   );
   gpc1_1 gpc686 (
      {stage0_42[60]},
      {stage1_42[25]}
   );
   gpc1_1 gpc687 (
      {stage0_42[61]},
      {stage1_42[26]}
   );
   gpc1_1 gpc688 (
      {stage0_42[62]},
      {stage1_42[27]}
   );
   gpc1_1 gpc689 (
      {stage0_42[63]},
      {stage1_42[28]}
   );
   gpc1_1 gpc690 (
      {stage0_43[50]},
      {stage1_43[22]}
   );
   gpc1_1 gpc691 (
      {stage0_43[51]},
      {stage1_43[23]}
   );
   gpc1_1 gpc692 (
      {stage0_43[52]},
      {stage1_43[24]}
   );
   gpc1_1 gpc693 (
      {stage0_43[53]},
      {stage1_43[25]}
   );
   gpc1_1 gpc694 (
      {stage0_43[54]},
      {stage1_43[26]}
   );
   gpc1_1 gpc695 (
      {stage0_43[55]},
      {stage1_43[27]}
   );
   gpc1_1 gpc696 (
      {stage0_43[56]},
      {stage1_43[28]}
   );
   gpc1_1 gpc697 (
      {stage0_43[57]},
      {stage1_43[29]}
   );
   gpc1_1 gpc698 (
      {stage0_43[58]},
      {stage1_43[30]}
   );
   gpc1_1 gpc699 (
      {stage0_43[59]},
      {stage1_43[31]}
   );
   gpc1_1 gpc700 (
      {stage0_43[60]},
      {stage1_43[32]}
   );
   gpc1_1 gpc701 (
      {stage0_43[61]},
      {stage1_43[33]}
   );
   gpc1_1 gpc702 (
      {stage0_43[62]},
      {stage1_43[34]}
   );
   gpc1_1 gpc703 (
      {stage0_43[63]},
      {stage1_43[35]}
   );
   gpc1_1 gpc704 (
      {stage0_44[58]},
      {stage1_44[27]}
   );
   gpc1_1 gpc705 (
      {stage0_44[59]},
      {stage1_44[28]}
   );
   gpc1_1 gpc706 (
      {stage0_44[60]},
      {stage1_44[29]}
   );
   gpc1_1 gpc707 (
      {stage0_44[61]},
      {stage1_44[30]}
   );
   gpc1_1 gpc708 (
      {stage0_44[62]},
      {stage1_44[31]}
   );
   gpc1_1 gpc709 (
      {stage0_44[63]},
      {stage1_44[32]}
   );
   gpc1_1 gpc710 (
      {stage0_45[36]},
      {stage1_45[20]}
   );
   gpc1_1 gpc711 (
      {stage0_45[37]},
      {stage1_45[21]}
   );
   gpc1_1 gpc712 (
      {stage0_45[38]},
      {stage1_45[22]}
   );
   gpc1_1 gpc713 (
      {stage0_45[39]},
      {stage1_45[23]}
   );
   gpc1_1 gpc714 (
      {stage0_45[40]},
      {stage1_45[24]}
   );
   gpc1_1 gpc715 (
      {stage0_45[41]},
      {stage1_45[25]}
   );
   gpc1_1 gpc716 (
      {stage0_45[42]},
      {stage1_45[26]}
   );
   gpc1_1 gpc717 (
      {stage0_45[43]},
      {stage1_45[27]}
   );
   gpc1_1 gpc718 (
      {stage0_45[44]},
      {stage1_45[28]}
   );
   gpc1_1 gpc719 (
      {stage0_45[45]},
      {stage1_45[29]}
   );
   gpc1_1 gpc720 (
      {stage0_45[46]},
      {stage1_45[30]}
   );
   gpc1_1 gpc721 (
      {stage0_45[47]},
      {stage1_45[31]}
   );
   gpc1_1 gpc722 (
      {stage0_45[48]},
      {stage1_45[32]}
   );
   gpc1_1 gpc723 (
      {stage0_45[49]},
      {stage1_45[33]}
   );
   gpc1_1 gpc724 (
      {stage0_45[50]},
      {stage1_45[34]}
   );
   gpc1_1 gpc725 (
      {stage0_45[51]},
      {stage1_45[35]}
   );
   gpc1_1 gpc726 (
      {stage0_45[52]},
      {stage1_45[36]}
   );
   gpc1_1 gpc727 (
      {stage0_45[53]},
      {stage1_45[37]}
   );
   gpc1_1 gpc728 (
      {stage0_45[54]},
      {stage1_45[38]}
   );
   gpc1_1 gpc729 (
      {stage0_45[55]},
      {stage1_45[39]}
   );
   gpc1_1 gpc730 (
      {stage0_45[56]},
      {stage1_45[40]}
   );
   gpc1_1 gpc731 (
      {stage0_45[57]},
      {stage1_45[41]}
   );
   gpc1_1 gpc732 (
      {stage0_45[58]},
      {stage1_45[42]}
   );
   gpc1_1 gpc733 (
      {stage0_45[59]},
      {stage1_45[43]}
   );
   gpc1_1 gpc734 (
      {stage0_45[60]},
      {stage1_45[44]}
   );
   gpc1_1 gpc735 (
      {stage0_45[61]},
      {stage1_45[45]}
   );
   gpc1_1 gpc736 (
      {stage0_45[62]},
      {stage1_45[46]}
   );
   gpc1_1 gpc737 (
      {stage0_45[63]},
      {stage1_45[47]}
   );
   gpc1_1 gpc738 (
      {stage0_47[46]},
      {stage1_47[23]}
   );
   gpc1_1 gpc739 (
      {stage0_47[47]},
      {stage1_47[24]}
   );
   gpc1_1 gpc740 (
      {stage0_47[48]},
      {stage1_47[25]}
   );
   gpc1_1 gpc741 (
      {stage0_47[49]},
      {stage1_47[26]}
   );
   gpc1_1 gpc742 (
      {stage0_47[50]},
      {stage1_47[27]}
   );
   gpc1_1 gpc743 (
      {stage0_47[51]},
      {stage1_47[28]}
   );
   gpc1_1 gpc744 (
      {stage0_47[52]},
      {stage1_47[29]}
   );
   gpc1_1 gpc745 (
      {stage0_47[53]},
      {stage1_47[30]}
   );
   gpc1_1 gpc746 (
      {stage0_47[54]},
      {stage1_47[31]}
   );
   gpc1_1 gpc747 (
      {stage0_47[55]},
      {stage1_47[32]}
   );
   gpc1_1 gpc748 (
      {stage0_47[56]},
      {stage1_47[33]}
   );
   gpc1_1 gpc749 (
      {stage0_47[57]},
      {stage1_47[34]}
   );
   gpc1_1 gpc750 (
      {stage0_47[58]},
      {stage1_47[35]}
   );
   gpc1_1 gpc751 (
      {stage0_47[59]},
      {stage1_47[36]}
   );
   gpc1_1 gpc752 (
      {stage0_47[60]},
      {stage1_47[37]}
   );
   gpc1_1 gpc753 (
      {stage0_47[61]},
      {stage1_47[38]}
   );
   gpc1_1 gpc754 (
      {stage0_47[62]},
      {stage1_47[39]}
   );
   gpc1_1 gpc755 (
      {stage0_47[63]},
      {stage1_47[40]}
   );
   gpc1_1 gpc756 (
      {stage0_48[58]},
      {stage1_48[26]}
   );
   gpc1_1 gpc757 (
      {stage0_48[59]},
      {stage1_48[27]}
   );
   gpc1_1 gpc758 (
      {stage0_48[60]},
      {stage1_48[28]}
   );
   gpc1_1 gpc759 (
      {stage0_48[61]},
      {stage1_48[29]}
   );
   gpc1_1 gpc760 (
      {stage0_48[62]},
      {stage1_48[30]}
   );
   gpc1_1 gpc761 (
      {stage0_48[63]},
      {stage1_48[31]}
   );
   gpc1_1 gpc762 (
      {stage0_49[60]},
      {stage1_49[21]}
   );
   gpc1_1 gpc763 (
      {stage0_49[61]},
      {stage1_49[22]}
   );
   gpc1_1 gpc764 (
      {stage0_49[62]},
      {stage1_49[23]}
   );
   gpc1_1 gpc765 (
      {stage0_49[63]},
      {stage1_49[24]}
   );
   gpc1_1 gpc766 (
      {stage0_50[62]},
      {stage1_50[23]}
   );
   gpc1_1 gpc767 (
      {stage0_50[63]},
      {stage1_50[24]}
   );
   gpc1_1 gpc768 (
      {stage0_51[59]},
      {stage1_51[27]}
   );
   gpc1_1 gpc769 (
      {stage0_51[60]},
      {stage1_51[28]}
   );
   gpc1_1 gpc770 (
      {stage0_51[61]},
      {stage1_51[29]}
   );
   gpc1_1 gpc771 (
      {stage0_51[62]},
      {stage1_51[30]}
   );
   gpc1_1 gpc772 (
      {stage0_51[63]},
      {stage1_51[31]}
   );
   gpc1_1 gpc773 (
      {stage0_52[45]},
      {stage1_52[24]}
   );
   gpc1_1 gpc774 (
      {stage0_52[46]},
      {stage1_52[25]}
   );
   gpc1_1 gpc775 (
      {stage0_52[47]},
      {stage1_52[26]}
   );
   gpc1_1 gpc776 (
      {stage0_52[48]},
      {stage1_52[27]}
   );
   gpc1_1 gpc777 (
      {stage0_52[49]},
      {stage1_52[28]}
   );
   gpc1_1 gpc778 (
      {stage0_52[50]},
      {stage1_52[29]}
   );
   gpc1_1 gpc779 (
      {stage0_52[51]},
      {stage1_52[30]}
   );
   gpc1_1 gpc780 (
      {stage0_52[52]},
      {stage1_52[31]}
   );
   gpc1_1 gpc781 (
      {stage0_52[53]},
      {stage1_52[32]}
   );
   gpc1_1 gpc782 (
      {stage0_52[54]},
      {stage1_52[33]}
   );
   gpc1_1 gpc783 (
      {stage0_52[55]},
      {stage1_52[34]}
   );
   gpc1_1 gpc784 (
      {stage0_52[56]},
      {stage1_52[35]}
   );
   gpc1_1 gpc785 (
      {stage0_52[57]},
      {stage1_52[36]}
   );
   gpc1_1 gpc786 (
      {stage0_52[58]},
      {stage1_52[37]}
   );
   gpc1_1 gpc787 (
      {stage0_52[59]},
      {stage1_52[38]}
   );
   gpc1_1 gpc788 (
      {stage0_52[60]},
      {stage1_52[39]}
   );
   gpc1_1 gpc789 (
      {stage0_52[61]},
      {stage1_52[40]}
   );
   gpc1_1 gpc790 (
      {stage0_52[62]},
      {stage1_52[41]}
   );
   gpc1_1 gpc791 (
      {stage0_52[63]},
      {stage1_52[42]}
   );
   gpc1_1 gpc792 (
      {stage0_53[58]},
      {stage1_53[21]}
   );
   gpc1_1 gpc793 (
      {stage0_53[59]},
      {stage1_53[22]}
   );
   gpc1_1 gpc794 (
      {stage0_53[60]},
      {stage1_53[23]}
   );
   gpc1_1 gpc795 (
      {stage0_53[61]},
      {stage1_53[24]}
   );
   gpc1_1 gpc796 (
      {stage0_53[62]},
      {stage1_53[25]}
   );
   gpc1_1 gpc797 (
      {stage0_53[63]},
      {stage1_53[26]}
   );
   gpc1_1 gpc798 (
      {stage0_54[54]},
      {stage1_54[23]}
   );
   gpc1_1 gpc799 (
      {stage0_54[55]},
      {stage1_54[24]}
   );
   gpc1_1 gpc800 (
      {stage0_54[56]},
      {stage1_54[25]}
   );
   gpc1_1 gpc801 (
      {stage0_54[57]},
      {stage1_54[26]}
   );
   gpc1_1 gpc802 (
      {stage0_54[58]},
      {stage1_54[27]}
   );
   gpc1_1 gpc803 (
      {stage0_54[59]},
      {stage1_54[28]}
   );
   gpc1_1 gpc804 (
      {stage0_54[60]},
      {stage1_54[29]}
   );
   gpc1_1 gpc805 (
      {stage0_54[61]},
      {stage1_54[30]}
   );
   gpc1_1 gpc806 (
      {stage0_54[62]},
      {stage1_54[31]}
   );
   gpc1_1 gpc807 (
      {stage0_54[63]},
      {stage1_54[32]}
   );
   gpc1_1 gpc808 (
      {stage0_56[62]},
      {stage1_56[24]}
   );
   gpc1_1 gpc809 (
      {stage0_56[63]},
      {stage1_56[25]}
   );
   gpc1_1 gpc810 (
      {stage0_58[47]},
      {stage1_58[24]}
   );
   gpc1_1 gpc811 (
      {stage0_58[48]},
      {stage1_58[25]}
   );
   gpc1_1 gpc812 (
      {stage0_58[49]},
      {stage1_58[26]}
   );
   gpc1_1 gpc813 (
      {stage0_58[50]},
      {stage1_58[27]}
   );
   gpc1_1 gpc814 (
      {stage0_58[51]},
      {stage1_58[28]}
   );
   gpc1_1 gpc815 (
      {stage0_58[52]},
      {stage1_58[29]}
   );
   gpc1_1 gpc816 (
      {stage0_58[53]},
      {stage1_58[30]}
   );
   gpc1_1 gpc817 (
      {stage0_58[54]},
      {stage1_58[31]}
   );
   gpc1_1 gpc818 (
      {stage0_58[55]},
      {stage1_58[32]}
   );
   gpc1_1 gpc819 (
      {stage0_58[56]},
      {stage1_58[33]}
   );
   gpc1_1 gpc820 (
      {stage0_58[57]},
      {stage1_58[34]}
   );
   gpc1_1 gpc821 (
      {stage0_58[58]},
      {stage1_58[35]}
   );
   gpc1_1 gpc822 (
      {stage0_58[59]},
      {stage1_58[36]}
   );
   gpc1_1 gpc823 (
      {stage0_58[60]},
      {stage1_58[37]}
   );
   gpc1_1 gpc824 (
      {stage0_58[61]},
      {stage1_58[38]}
   );
   gpc1_1 gpc825 (
      {stage0_58[62]},
      {stage1_58[39]}
   );
   gpc1_1 gpc826 (
      {stage0_58[63]},
      {stage1_58[40]}
   );
   gpc1_1 gpc827 (
      {stage0_59[42]},
      {stage1_59[20]}
   );
   gpc1_1 gpc828 (
      {stage0_59[43]},
      {stage1_59[21]}
   );
   gpc1_1 gpc829 (
      {stage0_59[44]},
      {stage1_59[22]}
   );
   gpc1_1 gpc830 (
      {stage0_59[45]},
      {stage1_59[23]}
   );
   gpc1_1 gpc831 (
      {stage0_59[46]},
      {stage1_59[24]}
   );
   gpc1_1 gpc832 (
      {stage0_59[47]},
      {stage1_59[25]}
   );
   gpc1_1 gpc833 (
      {stage0_59[48]},
      {stage1_59[26]}
   );
   gpc1_1 gpc834 (
      {stage0_59[49]},
      {stage1_59[27]}
   );
   gpc1_1 gpc835 (
      {stage0_59[50]},
      {stage1_59[28]}
   );
   gpc1_1 gpc836 (
      {stage0_59[51]},
      {stage1_59[29]}
   );
   gpc1_1 gpc837 (
      {stage0_59[52]},
      {stage1_59[30]}
   );
   gpc1_1 gpc838 (
      {stage0_59[53]},
      {stage1_59[31]}
   );
   gpc1_1 gpc839 (
      {stage0_59[54]},
      {stage1_59[32]}
   );
   gpc1_1 gpc840 (
      {stage0_59[55]},
      {stage1_59[33]}
   );
   gpc1_1 gpc841 (
      {stage0_59[56]},
      {stage1_59[34]}
   );
   gpc1_1 gpc842 (
      {stage0_59[57]},
      {stage1_59[35]}
   );
   gpc1_1 gpc843 (
      {stage0_59[58]},
      {stage1_59[36]}
   );
   gpc1_1 gpc844 (
      {stage0_59[59]},
      {stage1_59[37]}
   );
   gpc1_1 gpc845 (
      {stage0_59[60]},
      {stage1_59[38]}
   );
   gpc1_1 gpc846 (
      {stage0_59[61]},
      {stage1_59[39]}
   );
   gpc1_1 gpc847 (
      {stage0_59[62]},
      {stage1_59[40]}
   );
   gpc1_1 gpc848 (
      {stage0_59[63]},
      {stage1_59[41]}
   );
   gpc1_1 gpc849 (
      {stage0_60[52]},
      {stage1_60[21]}
   );
   gpc1_1 gpc850 (
      {stage0_60[53]},
      {stage1_60[22]}
   );
   gpc1_1 gpc851 (
      {stage0_60[54]},
      {stage1_60[23]}
   );
   gpc1_1 gpc852 (
      {stage0_60[55]},
      {stage1_60[24]}
   );
   gpc1_1 gpc853 (
      {stage0_60[56]},
      {stage1_60[25]}
   );
   gpc1_1 gpc854 (
      {stage0_60[57]},
      {stage1_60[26]}
   );
   gpc1_1 gpc855 (
      {stage0_60[58]},
      {stage1_60[27]}
   );
   gpc1_1 gpc856 (
      {stage0_60[59]},
      {stage1_60[28]}
   );
   gpc1_1 gpc857 (
      {stage0_60[60]},
      {stage1_60[29]}
   );
   gpc1_1 gpc858 (
      {stage0_60[61]},
      {stage1_60[30]}
   );
   gpc1_1 gpc859 (
      {stage0_60[62]},
      {stage1_60[31]}
   );
   gpc1_1 gpc860 (
      {stage0_60[63]},
      {stage1_60[32]}
   );
   gpc1_1 gpc861 (
      {stage0_61[58]},
      {stage1_61[25]}
   );
   gpc1_1 gpc862 (
      {stage0_61[59]},
      {stage1_61[26]}
   );
   gpc1_1 gpc863 (
      {stage0_61[60]},
      {stage1_61[27]}
   );
   gpc1_1 gpc864 (
      {stage0_61[61]},
      {stage1_61[28]}
   );
   gpc1_1 gpc865 (
      {stage0_61[62]},
      {stage1_61[29]}
   );
   gpc1_1 gpc866 (
      {stage0_61[63]},
      {stage1_61[30]}
   );
   gpc1_1 gpc867 (
      {stage0_62[51]},
      {stage1_62[20]}
   );
   gpc1_1 gpc868 (
      {stage0_62[52]},
      {stage1_62[21]}
   );
   gpc1_1 gpc869 (
      {stage0_62[53]},
      {stage1_62[22]}
   );
   gpc1_1 gpc870 (
      {stage0_62[54]},
      {stage1_62[23]}
   );
   gpc1_1 gpc871 (
      {stage0_62[55]},
      {stage1_62[24]}
   );
   gpc1_1 gpc872 (
      {stage0_62[56]},
      {stage1_62[25]}
   );
   gpc1_1 gpc873 (
      {stage0_62[57]},
      {stage1_62[26]}
   );
   gpc1_1 gpc874 (
      {stage0_62[58]},
      {stage1_62[27]}
   );
   gpc1_1 gpc875 (
      {stage0_62[59]},
      {stage1_62[28]}
   );
   gpc1_1 gpc876 (
      {stage0_62[60]},
      {stage1_62[29]}
   );
   gpc1_1 gpc877 (
      {stage0_62[61]},
      {stage1_62[30]}
   );
   gpc1_1 gpc878 (
      {stage0_62[62]},
      {stage1_62[31]}
   );
   gpc1_1 gpc879 (
      {stage0_62[63]},
      {stage1_62[32]}
   );
   gpc1_1 gpc880 (
      {stage0_63[54]},
      {stage1_63[18]}
   );
   gpc1_1 gpc881 (
      {stage0_63[55]},
      {stage1_63[19]}
   );
   gpc1_1 gpc882 (
      {stage0_63[56]},
      {stage1_63[20]}
   );
   gpc1_1 gpc883 (
      {stage0_63[57]},
      {stage1_63[21]}
   );
   gpc1_1 gpc884 (
      {stage0_63[58]},
      {stage1_63[22]}
   );
   gpc1_1 gpc885 (
      {stage0_63[59]},
      {stage1_63[23]}
   );
   gpc1_1 gpc886 (
      {stage0_63[60]},
      {stage1_63[24]}
   );
   gpc1_1 gpc887 (
      {stage0_63[61]},
      {stage1_63[25]}
   );
   gpc1_1 gpc888 (
      {stage0_63[62]},
      {stage1_63[26]}
   );
   gpc1_1 gpc889 (
      {stage0_63[63]},
      {stage1_63[27]}
   );
   gpc1163_5 gpc890 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc891 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc892 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc893 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc894 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc895 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], 1'b0, 1'b0},
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc896 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc897 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc898 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc899 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc900 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc901 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[12]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[11],stage2_3[11]}
   );
   gpc1163_5 gpc902 (
      {stage1_4[13], stage1_4[14], stage1_4[15]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[12]}
   );
   gpc606_5 gpc903 (
      {stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[13]}
   );
   gpc1325_5 gpc904 (
      {stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_5[12], stage1_5[13]},
      {stage1_6[7], stage1_6[8], stage1_6[9]},
      {stage1_7[1]},
      {stage2_8[2],stage2_7[3],stage2_6[5],stage2_5[8],stage2_4[14]}
   );
   gpc615_5 gpc905 (
      {stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13], stage1_6[14]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[3],stage2_7[4],stage2_6[6]}
   );
   gpc117_4 gpc906 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage1_8[6]},
      {stage1_9[0]},
      {stage2_10[1],stage2_9[1],stage2_8[4],stage2_7[5]}
   );
   gpc615_5 gpc907 (
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14]},
      {stage1_8[7]},
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[5],stage2_7[6]}
   );
   gpc615_5 gpc908 (
      {stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage1_8[8]},
      {stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11], stage1_9[12]},
      {stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[6],stage2_7[7]}
   );
   gpc615_5 gpc909 (
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage1_8[9]},
      {stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18]},
      {stage2_11[2],stage2_10[4],stage2_9[4],stage2_8[7],stage2_7[8]}
   );
   gpc606_5 gpc910 (
      {stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[3],stage2_10[5],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc911 (
      {stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc912 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[5],stage2_10[7]}
   );
   gpc615_5 gpc913 (
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[6]}
   );
   gpc615_5 gpc914 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4],stage2_11[7]}
   );
   gpc615_5 gpc915 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[4],stage2_12[5],stage2_11[8]}
   );
   gpc615_5 gpc916 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[5],stage2_12[6],stage2_11[9]}
   );
   gpc606_5 gpc917 (
      {stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[4],stage2_14[5],stage2_13[6],stage2_12[7]}
   );
   gpc615_5 gpc918 (
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28]},
      {stage1_14[6]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[5],stage2_14[6],stage2_13[7]}
   );
   gpc615_5 gpc919 (
      {stage1_13[29], stage1_13[30], 1'b0, 1'b0, 1'b0},
      {stage1_14[7]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[2],stage2_15[6],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc920 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[3],stage2_15[7],stage2_14[8]}
   );
   gpc615_5 gpc921 (
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[12]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[4],stage2_15[8],stage2_14[9]}
   );
   gpc615_5 gpc922 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[12]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[5],stage2_15[9]}
   );
   gpc615_5 gpc923 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22]},
      {stage1_16[13]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[6],stage2_15[10]}
   );
   gpc615_5 gpc924 (
      {stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage1_16[14]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[7],stage2_15[11]}
   );
   gpc615_5 gpc925 (
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32]},
      {stage1_16[15]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[8],stage2_15[12]}
   );
   gpc615_5 gpc926 (
      {stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[16]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[9],stage2_15[13]}
   );
   gpc615_5 gpc927 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21]},
      {stage1_17[30]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[10]}
   );
   gpc615_5 gpc928 (
      {stage1_16[22], stage1_16[23], stage1_16[24], stage1_16[25], stage1_16[26]},
      {stage1_17[31]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[11]}
   );
   gpc623_5 gpc929 (
      {stage1_17[32], stage1_17[33], stage1_17[34]},
      {stage1_18[12], stage1_18[13]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[7],stage2_18[9],stage2_17[11]}
   );
   gpc615_5 gpc930 (
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[8]}
   );
   gpc615_5 gpc931 (
      {stage1_19[11], stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[2],stage2_20[4],stage2_19[9]}
   );
   gpc615_5 gpc932 (
      {stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19], stage1_19[20]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[3],stage2_20[5],stage2_19[10]}
   );
   gpc615_5 gpc933 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[4],stage2_20[6],stage2_19[11]}
   );
   gpc606_5 gpc934 (
      {stage1_20[4], stage1_20[5], stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[4],stage2_22[4],stage2_21[5],stage2_20[7]}
   );
   gpc606_5 gpc935 (
      {stage1_20[10], stage1_20[11], stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[5],stage2_22[5],stage2_21[6],stage2_20[8]}
   );
   gpc606_5 gpc936 (
      {stage1_20[16], stage1_20[17], stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[6],stage2_22[6],stage2_21[7],stage2_20[9]}
   );
   gpc606_5 gpc937 (
      {stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[7],stage2_22[7],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc938 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[4],stage2_23[8],stage2_22[8],stage2_21[9]}
   );
   gpc1415_5 gpc939 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[6]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[1],stage2_24[5],stage2_23[9],stage2_22[9]}
   );
   gpc623_5 gpc940 (
      {stage1_22[29], stage1_22[30], 1'b0},
      {stage1_23[7], stage1_23[8]},
      {stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9]},
      {stage2_26[1],stage2_25[2],stage2_24[6],stage2_23[10],stage2_22[10]}
   );
   gpc615_5 gpc941 (
      {stage1_23[9], stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13]},
      {stage1_24[10]},
      {stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[7],stage2_23[11]}
   );
   gpc615_5 gpc942 (
      {stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17], stage1_23[18]},
      {stage1_24[11]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[8],stage2_23[12]}
   );
   gpc615_5 gpc943 (
      {stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage1_24[12]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[9],stage2_23[13]}
   );
   gpc615_5 gpc944 (
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28]},
      {stage1_24[13]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[3],stage2_26[5],stage2_25[6],stage2_24[10],stage2_23[14]}
   );
   gpc615_5 gpc945 (
      {stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33]},
      {stage1_24[14]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[4],stage2_26[6],stage2_25[7],stage2_24[11],stage2_23[15]}
   );
   gpc606_5 gpc946 (
      {stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19], stage1_24[20]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[7],stage2_25[8],stage2_24[12]}
   );
   gpc606_5 gpc947 (
      {stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25], stage1_24[26]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[8],stage2_25[9],stage2_24[13]}
   );
   gpc606_5 gpc948 (
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[9],stage2_25[10]}
   );
   gpc606_5 gpc949 (
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[10],stage2_25[11]}
   );
   gpc615_5 gpc950 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16]},
      {stage1_27[12]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[11]}
   );
   gpc615_5 gpc951 (
      {stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21]},
      {stage1_27[13]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[12]}
   );
   gpc615_5 gpc952 (
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18]},
      {stage1_28[12]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[2],stage2_29[4],stage2_28[6],stage2_27[11]}
   );
   gpc615_5 gpc953 (
      {stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage1_28[13]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[3],stage2_29[5],stage2_28[7],stage2_27[12]}
   );
   gpc615_5 gpc954 (
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28]},
      {stage1_28[14]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[4],stage2_29[6],stage2_28[8],stage2_27[13]}
   );
   gpc606_5 gpc955 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[3],stage2_30[5],stage2_29[7],stage2_28[9]}
   );
   gpc606_5 gpc956 (
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[4],stage2_30[6],stage2_29[8]}
   );
   gpc606_5 gpc957 (
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], 1'b0},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[5],stage2_30[7],stage2_29[9]}
   );
   gpc615_5 gpc958 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10]},
      {stage1_31[12]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[2],stage2_32[3],stage2_31[6],stage2_30[8]}
   );
   gpc615_5 gpc959 (
      {stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15]},
      {stage1_31[13]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[3],stage2_32[4],stage2_31[7],stage2_30[9]}
   );
   gpc615_5 gpc960 (
      {stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17], stage1_31[18]},
      {stage1_32[12]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[4],stage2_32[5],stage2_31[8]}
   );
   gpc606_5 gpc961 (
      {stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17], stage1_32[18]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[1],stage2_34[3],stage2_33[5],stage2_32[6]}
   );
   gpc606_5 gpc962 (
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[1],stage2_35[2],stage2_34[4],stage2_33[6]}
   );
   gpc606_5 gpc963 (
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[2],stage2_35[3],stage2_34[5],stage2_33[7]}
   );
   gpc606_5 gpc964 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[3],stage2_35[4],stage2_34[6],stage2_33[8]}
   );
   gpc615_5 gpc965 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[18]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[3],stage2_36[4],stage2_35[5],stage2_34[7]}
   );
   gpc615_5 gpc966 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[19]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[4],stage2_36[5],stage2_35[6],stage2_34[8]}
   );
   gpc615_5 gpc967 (
      {stage1_34[16], stage1_34[17], stage1_34[18], stage1_34[19], stage1_34[20]},
      {stage1_35[20]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[5],stage2_36[6],stage2_35[7],stage2_34[9]}
   );
   gpc615_5 gpc968 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[6],stage2_36[7],stage2_35[8]}
   );
   gpc606_5 gpc969 (
      {stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[1],stage2_38[4],stage2_37[7],stage2_36[8]}
   );
   gpc606_5 gpc970 (
      {stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30]},
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11]},
      {stage2_40[1],stage2_39[2],stage2_38[5],stage2_37[8],stage2_36[9]}
   );
   gpc606_5 gpc971 (
      {stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36]},
      {stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17]},
      {stage2_40[2],stage2_39[3],stage2_38[6],stage2_37[9],stage2_36[10]}
   );
   gpc606_5 gpc972 (
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[3],stage2_39[4],stage2_38[7],stage2_37[10]}
   );
   gpc606_5 gpc973 (
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[4],stage2_39[5],stage2_38[8],stage2_37[11]}
   );
   gpc1406_5 gpc974 (
      {stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3]},
      {stage1_41[0]},
      {stage2_42[0],stage2_41[2],stage2_40[5],stage2_39[6],stage2_38[9]}
   );
   gpc1325_5 gpc975 (
      {stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28]},
      {stage1_39[12], stage1_39[13]},
      {stage1_40[4], stage1_40[5], stage1_40[6]},
      {stage1_41[1]},
      {stage2_42[1],stage2_41[3],stage2_40[6],stage2_39[7],stage2_38[10]}
   );
   gpc615_5 gpc976 (
      {stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage1_40[7]},
      {stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5], stage1_41[6], stage1_41[7]},
      {stage2_43[0],stage2_42[2],stage2_41[4],stage2_40[7],stage2_39[8]}
   );
   gpc606_5 gpc977 (
      {stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11], stage1_40[12], stage1_40[13]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[1],stage2_42[3],stage2_41[5],stage2_40[8]}
   );
   gpc606_5 gpc978 (
      {stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17], stage1_40[18], stage1_40[19]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[2],stage2_42[4],stage2_41[6],stage2_40[9]}
   );
   gpc606_5 gpc979 (
      {stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23], stage1_40[24], stage1_40[25]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[3],stage2_42[5],stage2_41[7],stage2_40[10]}
   );
   gpc7_3 gpc980 (
      {stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11], stage1_41[12], stage1_41[13], stage1_41[14]},
      {stage2_43[4],stage2_42[6],stage2_41[8]}
   );
   gpc606_5 gpc981 (
      {stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19], stage1_41[20]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[3],stage2_43[5],stage2_42[7],stage2_41[9]}
   );
   gpc606_5 gpc982 (
      {stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24], stage1_41[25], stage1_41[26]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[4],stage2_43[6],stage2_42[8],stage2_41[10]}
   );
   gpc606_5 gpc983 (
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[2],stage2_44[5],stage2_43[7],stage2_42[9]}
   );
   gpc615_5 gpc984 (
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[3],stage2_44[6],stage2_43[8]}
   );
   gpc615_5 gpc985 (
      {stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[4],stage2_44[7],stage2_43[9]}
   );
   gpc615_5 gpc986 (
      {stage1_43[22], stage1_43[23], stage1_43[24], stage1_43[25], stage1_43[26]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[5],stage2_44[8],stage2_43[10]}
   );
   gpc615_5 gpc987 (
      {stage1_43[27], stage1_43[28], stage1_43[29], stage1_43[30], stage1_43[31]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[6],stage2_44[9],stage2_43[11]}
   );
   gpc615_5 gpc988 (
      {stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35], 1'b0},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[7],stage2_44[10],stage2_43[12]}
   );
   gpc606_5 gpc989 (
      {stage1_44[11], stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[5],stage2_46[6],stage2_45[8],stage2_44[11]}
   );
   gpc606_5 gpc990 (
      {stage1_44[17], stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[6],stage2_46[7],stage2_45[9],stage2_44[12]}
   );
   gpc606_5 gpc991 (
      {stage1_44[23], stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], 1'b0},
      {stage2_48[2],stage2_47[7],stage2_46[8],stage2_45[10],stage2_44[13]}
   );
   gpc606_5 gpc992 (
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[8],stage2_46[9],stage2_45[11]}
   );
   gpc606_5 gpc993 (
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[9],stage2_46[10],stage2_45[12]}
   );
   gpc606_5 gpc994 (
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[5],stage2_47[10],stage2_46[11],stage2_45[13]}
   );
   gpc606_5 gpc995 (
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[3],stage2_48[6],stage2_47[11]}
   );
   gpc606_5 gpc996 (
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[4],stage2_48[7],stage2_47[12]}
   );
   gpc606_5 gpc997 (
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[2],stage2_49[5],stage2_48[8],stage2_47[13]}
   );
   gpc117_4 gpc998 (
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6]},
      {stage1_49[18]},
      {stage1_50[0]},
      {stage2_51[3],stage2_50[3],stage2_49[6],stage2_48[9]}
   );
   gpc117_4 gpc999 (
      {stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_49[19]},
      {stage1_50[1]},
      {stage2_51[4],stage2_50[4],stage2_49[7],stage2_48[10]}
   );
   gpc117_4 gpc1000 (
      {stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17], stage1_48[18], stage1_48[19], stage1_48[20]},
      {stage1_49[20]},
      {stage1_50[2]},
      {stage2_51[5],stage2_50[5],stage2_49[8],stage2_48[11]}
   );
   gpc207_4 gpc1001 (
      {stage1_48[21], stage1_48[22], stage1_48[23], stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27]},
      {stage1_50[3], stage1_50[4]},
      {stage2_51[6],stage2_50[6],stage2_49[9],stage2_48[12]}
   );
   gpc606_5 gpc1002 (
      {stage1_49[21], stage1_49[22], stage1_49[23], stage1_49[24], 1'b0, 1'b0},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[0],stage2_51[7],stage2_50[7],stage2_49[10]}
   );
   gpc615_5 gpc1003 (
      {stage1_50[5], stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9]},
      {stage1_51[6]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[1],stage2_52[1],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc1004 (
      {stage1_50[10], stage1_50[11], stage1_50[12], stage1_50[13], stage1_50[14]},
      {stage1_51[7]},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage2_54[1],stage2_53[2],stage2_52[2],stage2_51[9],stage2_50[9]}
   );
   gpc615_5 gpc1005 (
      {stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18], stage1_50[19]},
      {stage1_51[8]},
      {stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17]},
      {stage2_54[2],stage2_53[3],stage2_52[3],stage2_51[10],stage2_50[10]}
   );
   gpc615_5 gpc1006 (
      {stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_51[9]},
      {stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23]},
      {stage2_54[3],stage2_53[4],stage2_52[4],stage2_51[11],stage2_50[11]}
   );
   gpc2116_5 gpc1007 (
      {stage1_51[10], stage1_51[11], stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15]},
      {stage1_52[24]},
      {stage1_53[0]},
      {stage1_54[0], stage1_54[1]},
      {stage2_55[0],stage2_54[4],stage2_53[5],stage2_52[5],stage2_51[12]}
   );
   gpc2116_5 gpc1008 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_52[25]},
      {stage1_53[1]},
      {stage1_54[2], stage1_54[3]},
      {stage2_55[1],stage2_54[5],stage2_53[6],stage2_52[6],stage2_51[13]}
   );
   gpc615_5 gpc1009 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26]},
      {stage1_52[26]},
      {stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5], stage1_53[6], stage1_53[7]},
      {stage2_55[2],stage2_54[6],stage2_53[7],stage2_52[7],stage2_51[14]}
   );
   gpc615_5 gpc1010 (
      {stage1_51[27], stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31]},
      {stage1_52[27]},
      {stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13]},
      {stage2_55[3],stage2_54[7],stage2_53[8],stage2_52[8],stage2_51[15]}
   );
   gpc615_5 gpc1011 (
      {stage1_52[28], stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32]},
      {stage1_53[14]},
      {stage1_54[4], stage1_54[5], stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9]},
      {stage2_56[0],stage2_55[4],stage2_54[8],stage2_53[9],stage2_52[9]}
   );
   gpc615_5 gpc1012 (
      {stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36], stage1_52[37]},
      {stage1_53[15]},
      {stage1_54[10], stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage2_56[1],stage2_55[5],stage2_54[9],stage2_53[10],stage2_52[10]}
   );
   gpc615_5 gpc1013 (
      {stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_53[16]},
      {stage1_54[16], stage1_54[17], stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21]},
      {stage2_56[2],stage2_55[6],stage2_54[10],stage2_53[11],stage2_52[11]}
   );
   gpc615_5 gpc1014 (
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage1_54[22]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[3],stage2_55[7],stage2_54[11],stage2_53[12]}
   );
   gpc1163_5 gpc1015 (
      {stage1_54[23], stage1_54[24], stage1_54[25]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage1_56[0]},
      {stage1_57[0]},
      {stage2_58[0],stage2_57[1],stage2_56[4],stage2_55[8],stage2_54[12]}
   );
   gpc1163_5 gpc1016 (
      {stage1_54[26], stage1_54[27], stage1_54[28]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[1]},
      {stage1_57[1]},
      {stage2_58[1],stage2_57[2],stage2_56[5],stage2_55[9],stage2_54[13]}
   );
   gpc615_5 gpc1017 (
      {stage1_54[29], stage1_54[30], stage1_54[31], stage1_54[32], 1'b0},
      {stage1_55[18]},
      {stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5], stage1_56[6], stage1_56[7]},
      {stage2_58[2],stage2_57[3],stage2_56[6],stage2_55[10],stage2_54[14]}
   );
   gpc606_5 gpc1018 (
      {stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11], stage1_56[12], stage1_56[13]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[0],stage2_58[3],stage2_57[4],stage2_56[7]}
   );
   gpc606_5 gpc1019 (
      {stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17], stage1_56[18], stage1_56[19]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[1],stage2_58[4],stage2_57[5],stage2_56[8]}
   );
   gpc606_5 gpc1020 (
      {stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[2],stage2_58[5],stage2_57[6],stage2_56[9]}
   );
   gpc606_5 gpc1021 (
      {stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5], stage1_57[6], stage1_57[7]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[3],stage2_59[3],stage2_58[6],stage2_57[7]}
   );
   gpc615_5 gpc1022 (
      {stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11], stage1_57[12]},
      {stage1_58[18]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[4],stage2_59[4],stage2_58[7],stage2_57[8]}
   );
   gpc615_5 gpc1023 (
      {stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage1_58[19]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[5],stage2_59[5],stage2_58[8],stage2_57[9]}
   );
   gpc615_5 gpc1024 (
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22]},
      {stage1_58[20]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[6],stage2_59[6],stage2_58[9],stage2_57[10]}
   );
   gpc615_5 gpc1025 (
      {stage1_58[21], stage1_58[22], stage1_58[23], stage1_58[24], stage1_58[25]},
      {stage1_59[24]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[4],stage2_60[7],stage2_59[7],stage2_58[10]}
   );
   gpc615_5 gpc1026 (
      {stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29], stage1_58[30]},
      {stage1_59[25]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[5],stage2_60[8],stage2_59[8],stage2_58[11]}
   );
   gpc615_5 gpc1027 (
      {stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage1_59[26]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[6],stage2_60[9],stage2_59[9],stage2_58[12]}
   );
   gpc606_5 gpc1028 (
      {stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30], stage1_59[31], stage1_59[32]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[3],stage2_61[7],stage2_60[10],stage2_59[10]}
   );
   gpc615_5 gpc1029 (
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22]},
      {stage1_61[6]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[1],stage2_62[4],stage2_61[8],stage2_60[11]}
   );
   gpc615_5 gpc1030 (
      {stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage1_61[7]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[2],stage2_62[5],stage2_61[9],stage2_60[12]}
   );
   gpc615_5 gpc1031 (
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32]},
      {stage1_61[8]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[3],stage2_62[6],stage2_61[10],stage2_60[13]}
   );
   gpc2135_5 gpc1032 (
      {stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12], stage1_61[13]},
      {stage1_62[18], stage1_62[19], stage1_62[20]},
      {stage1_63[0]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[0],stage2_64[3],stage2_63[4],stage2_62[7],stage2_61[11]}
   );
   gpc2135_5 gpc1033 (
      {stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage1_63[1]},
      {stage1_64[2], stage1_64[3]},
      {stage2_65[1],stage2_64[4],stage2_63[5],stage2_62[8],stage2_61[12]}
   );
   gpc606_5 gpc1034 (
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6], stage1_63[7]},
      {stage2_65[2],stage2_64[5],stage2_63[6],stage2_62[9],stage2_61[13]}
   );
   gpc606_5 gpc1035 (
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12], stage1_63[13]},
      {stage2_65[3],stage2_64[6],stage2_63[7],stage2_62[10],stage2_61[14]}
   );
   gpc606_5 gpc1036 (
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9]},
      {stage2_66[0],stage2_65[4],stage2_64[7],stage2_63[8],stage2_62[11]}
   );
   gpc615_5 gpc1037 (
      {stage1_62[30], stage1_62[31], stage1_62[32], 1'b0, 1'b0},
      {stage1_63[14]},
      {stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15]},
      {stage2_66[1],stage2_65[5],stage2_64[8],stage2_63[9],stage2_62[12]}
   );
   gpc606_5 gpc1038 (
      {stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_65[0], stage1_65[1], stage1_65[2], stage1_65[3], stage1_65[4], stage1_65[5]},
      {stage2_67[0],stage2_66[2],stage2_65[6],stage2_64[9],stage2_63[10]}
   );
   gpc606_5 gpc1039 (
      {stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_65[6], stage1_65[7], stage1_65[8], 1'b0, 1'b0, 1'b0},
      {stage2_67[1],stage2_66[3],stage2_65[7],stage2_64[10],stage2_63[11]}
   );
   gpc1_1 gpc1040 (
      {stage1_2[23]},
      {stage2_2[11]}
   );
   gpc1_1 gpc1041 (
      {stage1_4[27]},
      {stage2_4[15]}
   );
   gpc1_1 gpc1042 (
      {stage1_4[28]},
      {stage2_4[16]}
   );
   gpc1_1 gpc1043 (
      {stage1_4[29]},
      {stage2_4[17]}
   );
   gpc1_1 gpc1044 (
      {stage1_4[30]},
      {stage2_4[18]}
   );
   gpc1_1 gpc1045 (
      {stage1_4[31]},
      {stage2_4[19]}
   );
   gpc1_1 gpc1046 (
      {stage1_4[32]},
      {stage2_4[20]}
   );
   gpc1_1 gpc1047 (
      {stage1_4[33]},
      {stage2_4[21]}
   );
   gpc1_1 gpc1048 (
      {stage1_4[34]},
      {stage2_4[22]}
   );
   gpc1_1 gpc1049 (
      {stage1_4[35]},
      {stage2_4[23]}
   );
   gpc1_1 gpc1050 (
      {stage1_4[36]},
      {stage2_4[24]}
   );
   gpc1_1 gpc1051 (
      {stage1_4[37]},
      {stage2_4[25]}
   );
   gpc1_1 gpc1052 (
      {stage1_5[14]},
      {stage2_5[9]}
   );
   gpc1_1 gpc1053 (
      {stage1_5[15]},
      {stage2_5[10]}
   );
   gpc1_1 gpc1054 (
      {stage1_5[16]},
      {stage2_5[11]}
   );
   gpc1_1 gpc1055 (
      {stage1_5[17]},
      {stage2_5[12]}
   );
   gpc1_1 gpc1056 (
      {stage1_5[18]},
      {stage2_5[13]}
   );
   gpc1_1 gpc1057 (
      {stage1_5[19]},
      {stage2_5[14]}
   );
   gpc1_1 gpc1058 (
      {stage1_5[20]},
      {stage2_5[15]}
   );
   gpc1_1 gpc1059 (
      {stage1_5[21]},
      {stage2_5[16]}
   );
   gpc1_1 gpc1060 (
      {stage1_5[22]},
      {stage2_5[17]}
   );
   gpc1_1 gpc1061 (
      {stage1_5[23]},
      {stage2_5[18]}
   );
   gpc1_1 gpc1062 (
      {stage1_5[24]},
      {stage2_5[19]}
   );
   gpc1_1 gpc1063 (
      {stage1_5[25]},
      {stage2_5[20]}
   );
   gpc1_1 gpc1064 (
      {stage1_5[26]},
      {stage2_5[21]}
   );
   gpc1_1 gpc1065 (
      {stage1_6[15]},
      {stage2_6[7]}
   );
   gpc1_1 gpc1066 (
      {stage1_6[16]},
      {stage2_6[8]}
   );
   gpc1_1 gpc1067 (
      {stage1_6[17]},
      {stage2_6[9]}
   );
   gpc1_1 gpc1068 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc1069 (
      {stage1_6[19]},
      {stage2_6[11]}
   );
   gpc1_1 gpc1070 (
      {stage1_6[20]},
      {stage2_6[12]}
   );
   gpc1_1 gpc1071 (
      {stage1_6[21]},
      {stage2_6[13]}
   );
   gpc1_1 gpc1072 (
      {stage1_7[25]},
      {stage2_7[9]}
   );
   gpc1_1 gpc1073 (
      {stage1_7[26]},
      {stage2_7[10]}
   );
   gpc1_1 gpc1074 (
      {stage1_7[27]},
      {stage2_7[11]}
   );
   gpc1_1 gpc1075 (
      {stage1_7[28]},
      {stage2_7[12]}
   );
   gpc1_1 gpc1076 (
      {stage1_7[29]},
      {stage2_7[13]}
   );
   gpc1_1 gpc1077 (
      {stage1_7[30]},
      {stage2_7[14]}
   );
   gpc1_1 gpc1078 (
      {stage1_7[31]},
      {stage2_7[15]}
   );
   gpc1_1 gpc1079 (
      {stage1_7[32]},
      {stage2_7[16]}
   );
   gpc1_1 gpc1080 (
      {stage1_7[33]},
      {stage2_7[17]}
   );
   gpc1_1 gpc1081 (
      {stage1_7[34]},
      {stage2_7[18]}
   );
   gpc1_1 gpc1082 (
      {stage1_7[35]},
      {stage2_7[19]}
   );
   gpc1_1 gpc1083 (
      {stage1_8[16]},
      {stage2_8[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_8[17]},
      {stage2_8[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_8[18]},
      {stage2_8[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_8[19]},
      {stage2_8[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_8[20]},
      {stage2_8[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_8[21]},
      {stage2_8[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_8[22]},
      {stage2_8[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_8[23]},
      {stage2_8[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_8[24]},
      {stage2_8[17]}
   );
   gpc1_1 gpc1092 (
      {stage1_8[25]},
      {stage2_8[18]}
   );
   gpc1_1 gpc1093 (
      {stage1_8[26]},
      {stage2_8[19]}
   );
   gpc1_1 gpc1094 (
      {stage1_9[25]},
      {stage2_9[7]}
   );
   gpc1_1 gpc1095 (
      {stage1_9[26]},
      {stage2_9[8]}
   );
   gpc1_1 gpc1096 (
      {stage1_9[27]},
      {stage2_9[9]}
   );
   gpc1_1 gpc1097 (
      {stage1_9[28]},
      {stage2_9[10]}
   );
   gpc1_1 gpc1098 (
      {stage1_10[11]},
      {stage2_10[8]}
   );
   gpc1_1 gpc1099 (
      {stage1_10[12]},
      {stage2_10[9]}
   );
   gpc1_1 gpc1100 (
      {stage1_10[13]},
      {stage2_10[10]}
   );
   gpc1_1 gpc1101 (
      {stage1_10[14]},
      {stage2_10[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_10[15]},
      {stage2_10[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_10[16]},
      {stage2_10[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_10[17]},
      {stage2_10[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_10[18]},
      {stage2_10[15]}
   );
   gpc1_1 gpc1106 (
      {stage1_10[19]},
      {stage2_10[16]}
   );
   gpc1_1 gpc1107 (
      {stage1_10[20]},
      {stage2_10[17]}
   );
   gpc1_1 gpc1108 (
      {stage1_10[21]},
      {stage2_10[18]}
   );
   gpc1_1 gpc1109 (
      {stage1_10[22]},
      {stage2_10[19]}
   );
   gpc1_1 gpc1110 (
      {stage1_10[23]},
      {stage2_10[20]}
   );
   gpc1_1 gpc1111 (
      {stage1_10[24]},
      {stage2_10[21]}
   );
   gpc1_1 gpc1112 (
      {stage1_10[25]},
      {stage2_10[22]}
   );
   gpc1_1 gpc1113 (
      {stage1_10[26]},
      {stage2_10[23]}
   );
   gpc1_1 gpc1114 (
      {stage1_10[27]},
      {stage2_10[24]}
   );
   gpc1_1 gpc1115 (
      {stage1_10[28]},
      {stage2_10[25]}
   );
   gpc1_1 gpc1116 (
      {stage1_10[29]},
      {stage2_10[26]}
   );
   gpc1_1 gpc1117 (
      {stage1_10[30]},
      {stage2_10[27]}
   );
   gpc1_1 gpc1118 (
      {stage1_10[31]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1119 (
      {stage1_10[32]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1120 (
      {stage1_10[33]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1121 (
      {stage1_11[27]},
      {stage2_11[10]}
   );
   gpc1_1 gpc1122 (
      {stage1_11[28]},
      {stage2_11[11]}
   );
   gpc1_1 gpc1123 (
      {stage1_11[29]},
      {stage2_11[12]}
   );
   gpc1_1 gpc1124 (
      {stage1_11[30]},
      {stage2_11[13]}
   );
   gpc1_1 gpc1125 (
      {stage1_11[31]},
      {stage2_11[14]}
   );
   gpc1_1 gpc1126 (
      {stage1_11[32]},
      {stage2_11[15]}
   );
   gpc1_1 gpc1127 (
      {stage1_12[16]},
      {stage2_12[8]}
   );
   gpc1_1 gpc1128 (
      {stage1_12[17]},
      {stage2_12[9]}
   );
   gpc1_1 gpc1129 (
      {stage1_12[18]},
      {stage2_12[10]}
   );
   gpc1_1 gpc1130 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc1131 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc1132 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc1133 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc1134 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc1135 (
      {stage1_12[24]},
      {stage2_12[16]}
   );
   gpc1_1 gpc1136 (
      {stage1_12[25]},
      {stage2_12[17]}
   );
   gpc1_1 gpc1137 (
      {stage1_12[26]},
      {stage2_12[18]}
   );
   gpc1_1 gpc1138 (
      {stage1_14[19]},
      {stage2_14[10]}
   );
   gpc1_1 gpc1139 (
      {stage1_14[20]},
      {stage2_14[11]}
   );
   gpc1_1 gpc1140 (
      {stage1_14[21]},
      {stage2_14[12]}
   );
   gpc1_1 gpc1141 (
      {stage1_14[22]},
      {stage2_14[13]}
   );
   gpc1_1 gpc1142 (
      {stage1_14[23]},
      {stage2_14[14]}
   );
   gpc1_1 gpc1143 (
      {stage1_14[24]},
      {stage2_14[15]}
   );
   gpc1_1 gpc1144 (
      {stage1_15[38]},
      {stage2_15[14]}
   );
   gpc1_1 gpc1145 (
      {stage1_15[39]},
      {stage2_15[15]}
   );
   gpc1_1 gpc1146 (
      {stage1_15[40]},
      {stage2_15[16]}
   );
   gpc1_1 gpc1147 (
      {stage1_15[41]},
      {stage2_15[17]}
   );
   gpc1_1 gpc1148 (
      {stage1_15[42]},
      {stage2_15[18]}
   );
   gpc1_1 gpc1149 (
      {stage1_15[43]},
      {stage2_15[19]}
   );
   gpc1_1 gpc1150 (
      {stage1_15[44]},
      {stage2_15[20]}
   );
   gpc1_1 gpc1151 (
      {stage1_16[27]},
      {stage2_16[12]}
   );
   gpc1_1 gpc1152 (
      {stage1_16[28]},
      {stage2_16[13]}
   );
   gpc1_1 gpc1153 (
      {stage1_16[29]},
      {stage2_16[14]}
   );
   gpc1_1 gpc1154 (
      {stage1_16[30]},
      {stage2_16[15]}
   );
   gpc1_1 gpc1155 (
      {stage1_17[35]},
      {stage2_17[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_17[36]},
      {stage2_17[13]}
   );
   gpc1_1 gpc1157 (
      {stage1_17[37]},
      {stage2_17[14]}
   );
   gpc1_1 gpc1158 (
      {stage1_17[38]},
      {stage2_17[15]}
   );
   gpc1_1 gpc1159 (
      {stage1_17[39]},
      {stage2_17[16]}
   );
   gpc1_1 gpc1160 (
      {stage1_17[40]},
      {stage2_17[17]}
   );
   gpc1_1 gpc1161 (
      {stage1_17[41]},
      {stage2_17[18]}
   );
   gpc1_1 gpc1162 (
      {stage1_17[42]},
      {stage2_17[19]}
   );
   gpc1_1 gpc1163 (
      {stage1_17[43]},
      {stage2_17[20]}
   );
   gpc1_1 gpc1164 (
      {stage1_17[44]},
      {stage2_17[21]}
   );
   gpc1_1 gpc1165 (
      {stage1_18[14]},
      {stage2_18[10]}
   );
   gpc1_1 gpc1166 (
      {stage1_18[15]},
      {stage2_18[11]}
   );
   gpc1_1 gpc1167 (
      {stage1_18[16]},
      {stage2_18[12]}
   );
   gpc1_1 gpc1168 (
      {stage1_18[17]},
      {stage2_18[13]}
   );
   gpc1_1 gpc1169 (
      {stage1_18[18]},
      {stage2_18[14]}
   );
   gpc1_1 gpc1170 (
      {stage1_18[19]},
      {stage2_18[15]}
   );
   gpc1_1 gpc1171 (
      {stage1_18[20]},
      {stage2_18[16]}
   );
   gpc1_1 gpc1172 (
      {stage1_18[21]},
      {stage2_18[17]}
   );
   gpc1_1 gpc1173 (
      {stage1_18[22]},
      {stage2_18[18]}
   );
   gpc1_1 gpc1174 (
      {stage1_19[26]},
      {stage2_19[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_19[27]},
      {stage2_19[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_19[28]},
      {stage2_19[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_20[28]},
      {stage2_20[11]}
   );
   gpc1_1 gpc1178 (
      {stage1_20[29]},
      {stage2_20[12]}
   );
   gpc1_1 gpc1179 (
      {stage1_20[30]},
      {stage2_20[13]}
   );
   gpc1_1 gpc1180 (
      {stage1_20[31]},
      {stage2_20[14]}
   );
   gpc1_1 gpc1181 (
      {stage1_20[32]},
      {stage2_20[15]}
   );
   gpc1_1 gpc1182 (
      {stage1_20[33]},
      {stage2_20[16]}
   );
   gpc1_1 gpc1183 (
      {stage1_20[34]},
      {stage2_20[17]}
   );
   gpc1_1 gpc1184 (
      {stage1_20[35]},
      {stage2_20[18]}
   );
   gpc1_1 gpc1185 (
      {stage1_20[36]},
      {stage2_20[19]}
   );
   gpc1_1 gpc1186 (
      {stage1_20[37]},
      {stage2_20[20]}
   );
   gpc1_1 gpc1187 (
      {stage1_20[38]},
      {stage2_20[21]}
   );
   gpc1_1 gpc1188 (
      {stage1_20[39]},
      {stage2_20[22]}
   );
   gpc1_1 gpc1189 (
      {stage1_20[40]},
      {stage2_20[23]}
   );
   gpc1_1 gpc1190 (
      {stage1_21[30]},
      {stage2_21[10]}
   );
   gpc1_1 gpc1191 (
      {stage1_21[31]},
      {stage2_21[11]}
   );
   gpc1_1 gpc1192 (
      {stage1_21[32]},
      {stage2_21[12]}
   );
   gpc1_1 gpc1193 (
      {stage1_23[34]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1194 (
      {stage1_25[43]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1195 (
      {stage1_25[44]},
      {stage2_25[13]}
   );
   gpc1_1 gpc1196 (
      {stage1_26[22]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1197 (
      {stage1_26[23]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1198 (
      {stage1_26[24]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1199 (
      {stage1_26[25]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1200 (
      {stage1_26[26]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1201 (
      {stage1_26[27]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1202 (
      {stage1_26[28]},
      {stage2_26[19]}
   );
   gpc1_1 gpc1203 (
      {stage1_27[29]},
      {stage2_27[14]}
   );
   gpc1_1 gpc1204 (
      {stage1_27[30]},
      {stage2_27[15]}
   );
   gpc1_1 gpc1205 (
      {stage1_27[31]},
      {stage2_27[16]}
   );
   gpc1_1 gpc1206 (
      {stage1_27[32]},
      {stage2_27[17]}
   );
   gpc1_1 gpc1207 (
      {stage1_27[33]},
      {stage2_27[18]}
   );
   gpc1_1 gpc1208 (
      {stage1_27[34]},
      {stage2_27[19]}
   );
   gpc1_1 gpc1209 (
      {stage1_27[35]},
      {stage2_27[20]}
   );
   gpc1_1 gpc1210 (
      {stage1_27[36]},
      {stage2_27[21]}
   );
   gpc1_1 gpc1211 (
      {stage1_27[37]},
      {stage2_27[22]}
   );
   gpc1_1 gpc1212 (
      {stage1_27[38]},
      {stage2_27[23]}
   );
   gpc1_1 gpc1213 (
      {stage1_27[39]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1214 (
      {stage1_27[40]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1215 (
      {stage1_28[21]},
      {stage2_28[10]}
   );
   gpc1_1 gpc1216 (
      {stage1_28[22]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1217 (
      {stage1_28[23]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1218 (
      {stage1_28[24]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1219 (
      {stage1_28[25]},
      {stage2_28[14]}
   );
   gpc1_1 gpc1220 (
      {stage1_28[26]},
      {stage2_28[15]}
   );
   gpc1_1 gpc1221 (
      {stage1_30[16]},
      {stage2_30[10]}
   );
   gpc1_1 gpc1222 (
      {stage1_30[17]},
      {stage2_30[11]}
   );
   gpc1_1 gpc1223 (
      {stage1_30[18]},
      {stage2_30[12]}
   );
   gpc1_1 gpc1224 (
      {stage1_30[19]},
      {stage2_30[13]}
   );
   gpc1_1 gpc1225 (
      {stage1_30[20]},
      {stage2_30[14]}
   );
   gpc1_1 gpc1226 (
      {stage1_30[21]},
      {stage2_30[15]}
   );
   gpc1_1 gpc1227 (
      {stage1_30[22]},
      {stage2_30[16]}
   );
   gpc1_1 gpc1228 (
      {stage1_30[23]},
      {stage2_30[17]}
   );
   gpc1_1 gpc1229 (
      {stage1_30[24]},
      {stage2_30[18]}
   );
   gpc1_1 gpc1230 (
      {stage1_30[25]},
      {stage2_30[19]}
   );
   gpc1_1 gpc1231 (
      {stage1_31[19]},
      {stage2_31[9]}
   );
   gpc1_1 gpc1232 (
      {stage1_31[20]},
      {stage2_31[10]}
   );
   gpc1_1 gpc1233 (
      {stage1_31[21]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1234 (
      {stage1_31[22]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1235 (
      {stage1_32[19]},
      {stage2_32[7]}
   );
   gpc1_1 gpc1236 (
      {stage1_32[20]},
      {stage2_32[8]}
   );
   gpc1_1 gpc1237 (
      {stage1_32[21]},
      {stage2_32[9]}
   );
   gpc1_1 gpc1238 (
      {stage1_32[22]},
      {stage2_32[10]}
   );
   gpc1_1 gpc1239 (
      {stage1_32[23]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1240 (
      {stage1_32[24]},
      {stage2_32[12]}
   );
   gpc1_1 gpc1241 (
      {stage1_32[25]},
      {stage2_32[13]}
   );
   gpc1_1 gpc1242 (
      {stage1_32[26]},
      {stage2_32[14]}
   );
   gpc1_1 gpc1243 (
      {stage1_32[27]},
      {stage2_32[15]}
   );
   gpc1_1 gpc1244 (
      {stage1_32[28]},
      {stage2_32[16]}
   );
   gpc1_1 gpc1245 (
      {stage1_32[29]},
      {stage2_32[17]}
   );
   gpc1_1 gpc1246 (
      {stage1_32[30]},
      {stage2_32[18]}
   );
   gpc1_1 gpc1247 (
      {stage1_33[24]},
      {stage2_33[9]}
   );
   gpc1_1 gpc1248 (
      {stage1_33[25]},
      {stage2_33[10]}
   );
   gpc1_1 gpc1249 (
      {stage1_33[26]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1250 (
      {stage1_33[27]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1251 (
      {stage1_33[28]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1252 (
      {stage1_33[29]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1253 (
      {stage1_33[30]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1254 (
      {stage1_33[31]},
      {stage2_33[16]}
   );
   gpc1_1 gpc1255 (
      {stage1_33[32]},
      {stage2_33[17]}
   );
   gpc1_1 gpc1256 (
      {stage1_33[33]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1257 (
      {stage1_33[34]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1258 (
      {stage1_33[35]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1259 (
      {stage1_33[36]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1260 (
      {stage1_33[37]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1261 (
      {stage1_34[21]},
      {stage2_34[10]}
   );
   gpc1_1 gpc1262 (
      {stage1_34[22]},
      {stage2_34[11]}
   );
   gpc1_1 gpc1263 (
      {stage1_34[23]},
      {stage2_34[12]}
   );
   gpc1_1 gpc1264 (
      {stage1_35[26]},
      {stage2_35[9]}
   );
   gpc1_1 gpc1265 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1266 (
      {stage1_35[28]},
      {stage2_35[11]}
   );
   gpc1_1 gpc1267 (
      {stage1_35[29]},
      {stage2_35[12]}
   );
   gpc1_1 gpc1268 (
      {stage1_36[37]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1269 (
      {stage1_36[38]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1270 (
      {stage1_36[39]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1271 (
      {stage1_36[40]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1272 (
      {stage1_36[41]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1273 (
      {stage1_36[42]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1274 (
      {stage1_36[43]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1275 (
      {stage1_37[18]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1276 (
      {stage1_37[19]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1277 (
      {stage1_37[20]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1278 (
      {stage1_37[21]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1279 (
      {stage1_37[22]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1280 (
      {stage1_37[23]},
      {stage2_37[17]}
   );
   gpc1_1 gpc1281 (
      {stage1_38[29]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1282 (
      {stage1_38[30]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1283 (
      {stage1_38[31]},
      {stage2_38[13]}
   );
   gpc1_1 gpc1284 (
      {stage1_38[32]},
      {stage2_38[14]}
   );
   gpc1_1 gpc1285 (
      {stage1_38[33]},
      {stage2_38[15]}
   );
   gpc1_1 gpc1286 (
      {stage1_38[34]},
      {stage2_38[16]}
   );
   gpc1_1 gpc1287 (
      {stage1_38[35]},
      {stage2_38[17]}
   );
   gpc1_1 gpc1288 (
      {stage1_38[36]},
      {stage2_38[18]}
   );
   gpc1_1 gpc1289 (
      {stage1_38[37]},
      {stage2_38[19]}
   );
   gpc1_1 gpc1290 (
      {stage1_38[38]},
      {stage2_38[20]}
   );
   gpc1_1 gpc1291 (
      {stage1_38[39]},
      {stage2_38[21]}
   );
   gpc1_1 gpc1292 (
      {stage1_38[40]},
      {stage2_38[22]}
   );
   gpc1_1 gpc1293 (
      {stage1_38[41]},
      {stage2_38[23]}
   );
   gpc1_1 gpc1294 (
      {stage1_39[19]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1295 (
      {stage1_39[20]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1296 (
      {stage1_39[21]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1297 (
      {stage1_39[22]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1298 (
      {stage1_40[26]},
      {stage2_40[11]}
   );
   gpc1_1 gpc1299 (
      {stage1_41[27]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1300 (
      {stage1_41[28]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1301 (
      {stage1_41[29]},
      {stage2_41[13]}
   );
   gpc1_1 gpc1302 (
      {stage1_41[30]},
      {stage2_41[14]}
   );
   gpc1_1 gpc1303 (
      {stage1_41[31]},
      {stage2_41[15]}
   );
   gpc1_1 gpc1304 (
      {stage1_41[32]},
      {stage2_41[16]}
   );
   gpc1_1 gpc1305 (
      {stage1_41[33]},
      {stage2_41[17]}
   );
   gpc1_1 gpc1306 (
      {stage1_41[34]},
      {stage2_41[18]}
   );
   gpc1_1 gpc1307 (
      {stage1_41[35]},
      {stage2_41[19]}
   );
   gpc1_1 gpc1308 (
      {stage1_42[24]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1309 (
      {stage1_42[25]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1310 (
      {stage1_42[26]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1311 (
      {stage1_42[27]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1312 (
      {stage1_42[28]},
      {stage2_42[14]}
   );
   gpc1_1 gpc1313 (
      {stage1_44[29]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1314 (
      {stage1_44[30]},
      {stage2_44[15]}
   );
   gpc1_1 gpc1315 (
      {stage1_44[31]},
      {stage2_44[16]}
   );
   gpc1_1 gpc1316 (
      {stage1_44[32]},
      {stage2_44[17]}
   );
   gpc1_1 gpc1317 (
      {stage1_47[36]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1318 (
      {stage1_47[37]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1319 (
      {stage1_47[38]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1320 (
      {stage1_47[39]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1321 (
      {stage1_47[40]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1322 (
      {stage1_48[28]},
      {stage2_48[13]}
   );
   gpc1_1 gpc1323 (
      {stage1_48[29]},
      {stage2_48[14]}
   );
   gpc1_1 gpc1324 (
      {stage1_48[30]},
      {stage2_48[15]}
   );
   gpc1_1 gpc1325 (
      {stage1_48[31]},
      {stage2_48[16]}
   );
   gpc1_1 gpc1326 (
      {stage1_53[22]},
      {stage2_53[13]}
   );
   gpc1_1 gpc1327 (
      {stage1_53[23]},
      {stage2_53[14]}
   );
   gpc1_1 gpc1328 (
      {stage1_53[24]},
      {stage2_53[15]}
   );
   gpc1_1 gpc1329 (
      {stage1_53[25]},
      {stage2_53[16]}
   );
   gpc1_1 gpc1330 (
      {stage1_53[26]},
      {stage2_53[17]}
   );
   gpc1_1 gpc1331 (
      {stage1_55[19]},
      {stage2_55[11]}
   );
   gpc1_1 gpc1332 (
      {stage1_55[20]},
      {stage2_55[12]}
   );
   gpc1_1 gpc1333 (
      {stage1_55[21]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1334 (
      {stage1_55[22]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1335 (
      {stage1_55[23]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1336 (
      {stage1_55[24]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1337 (
      {stage1_57[23]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1338 (
      {stage1_57[24]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1339 (
      {stage1_57[25]},
      {stage2_57[13]}
   );
   gpc1_1 gpc1340 (
      {stage1_58[36]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1341 (
      {stage1_58[37]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1342 (
      {stage1_58[38]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1343 (
      {stage1_58[39]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1344 (
      {stage1_58[40]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1345 (
      {stage1_59[33]},
      {stage2_59[11]}
   );
   gpc1_1 gpc1346 (
      {stage1_59[34]},
      {stage2_59[12]}
   );
   gpc1_1 gpc1347 (
      {stage1_59[35]},
      {stage2_59[13]}
   );
   gpc1_1 gpc1348 (
      {stage1_59[36]},
      {stage2_59[14]}
   );
   gpc1_1 gpc1349 (
      {stage1_59[37]},
      {stage2_59[15]}
   );
   gpc1_1 gpc1350 (
      {stage1_59[38]},
      {stage2_59[16]}
   );
   gpc1_1 gpc1351 (
      {stage1_59[39]},
      {stage2_59[17]}
   );
   gpc1_1 gpc1352 (
      {stage1_59[40]},
      {stage2_59[18]}
   );
   gpc1_1 gpc1353 (
      {stage1_59[41]},
      {stage2_59[19]}
   );
   gpc1_1 gpc1354 (
      {stage1_63[27]},
      {stage2_63[12]}
   );
   gpc606_5 gpc1355 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc1356 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc1357 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1358 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc606_5 gpc1359 (
      {stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4]}
   );
   gpc606_5 gpc1360 (
      {stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5]}
   );
   gpc606_5 gpc1361 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc606_5 gpc1362 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc1325_5 gpc1363 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], 1'b0},
      {stage2_6[12], stage2_6[13]},
      {stage2_7[12], stage2_7[13], stage2_7[14]},
      {stage2_8[0]},
      {stage3_9[2],stage3_8[4],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc606_5 gpc1364 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc1365 (
      {stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc1366 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[7]}
   );
   gpc606_5 gpc1367 (
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[3],stage3_10[3],stage3_9[6]}
   );
   gpc1163_5 gpc1368 (
      {stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[1],stage3_12[4],stage3_11[4],stage3_10[4]}
   );
   gpc615_5 gpc1369 (
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25]},
      {stage2_11[12]},
      {stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6]},
      {stage3_14[1],stage3_13[2],stage3_12[5],stage3_11[5],stage3_10[5]}
   );
   gpc615_5 gpc1370 (
      {stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_11[13]},
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage3_14[2],stage3_13[3],stage3_12[6],stage3_11[6],stage3_10[6]}
   );
   gpc606_5 gpc1371 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[7]}
   );
   gpc615_5 gpc1372 (
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_14[6]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[1],stage3_14[4],stage3_13[5]}
   );
   gpc615_5 gpc1373 (
      {stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[2],stage3_15[2],stage3_14[5]}
   );
   gpc615_5 gpc1374 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], 1'b0},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[3],stage3_15[3],stage3_14[6]}
   );
   gpc615_5 gpc1375 (
      {stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12]},
      {stage2_16[12]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[3],stage3_16[4],stage3_15[4]}
   );
   gpc615_5 gpc1376 (
      {stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage2_16[13]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[3],stage3_17[4],stage3_16[5],stage3_15[5]}
   );
   gpc606_5 gpc1377 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[2],stage3_18[4],stage3_17[5]}
   );
   gpc606_5 gpc1378 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], 1'b0, 1'b0},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[3],stage3_18[5],stage3_17[6]}
   );
   gpc615_5 gpc1379 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[2],stage3_20[2],stage3_19[4],stage3_18[6]}
   );
   gpc615_5 gpc1380 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[13]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[3],stage3_20[3],stage3_19[5],stage3_18[7]}
   );
   gpc615_5 gpc1381 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[14]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[4],stage3_20[4],stage3_19[6],stage3_18[8]}
   );
   gpc606_5 gpc1382 (
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[3],stage3_21[5],stage3_20[5]}
   );
   gpc606_5 gpc1383 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[1],stage3_22[4],stage3_21[6]}
   );
   gpc606_5 gpc1384 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[2],stage3_22[5],stage3_21[7]}
   );
   gpc615_5 gpc1385 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[3],stage3_23[3],stage3_22[6]}
   );
   gpc606_5 gpc1386 (
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[3],stage3_24[4]}
   );
   gpc606_5 gpc1387 (
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[4]}
   );
   gpc606_5 gpc1388 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[5]}
   );
   gpc135_4 gpc1389 (
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10]},
      {stage2_27[12], stage2_27[13], stage2_27[14]},
      {stage2_28[0]},
      {stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc135_4 gpc1390 (
      {stage2_26[11], stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15]},
      {stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage2_28[1]},
      {stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc135_4 gpc1391 (
      {stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20]},
      {stage2_28[2]},
      {stage3_29[4],stage3_28[5],stage3_27[5],stage3_26[6]}
   );
   gpc615_5 gpc1392 (
      {stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25]},
      {stage2_28[3]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[5],stage3_28[6],stage3_27[6]}
   );
   gpc606_5 gpc1393 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[1],stage3_29[6],stage3_28[7]}
   );
   gpc606_5 gpc1394 (
      {stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[2],stage3_29[7],stage3_28[8]}
   );
   gpc606_5 gpc1395 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], 1'b0, 1'b0},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[2],stage3_31[3],stage3_30[3],stage3_29[8]}
   );
   gpc615_5 gpc1396 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[3],stage3_31[4],stage3_30[4]}
   );
   gpc615_5 gpc1397 (
      {stage2_30[17], stage2_30[18], stage2_30[19], 1'b0, 1'b0},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[4],stage3_31[5],stage3_30[5]}
   );
   gpc615_5 gpc1398 (
      {stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12]},
      {stage2_32[12]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[2],stage3_33[3],stage3_32[5],stage3_31[6]}
   );
   gpc606_5 gpc1399 (
      {stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[1],stage3_34[3],stage3_33[4],stage3_32[6]}
   );
   gpc606_5 gpc1400 (
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[2],stage3_34[4],stage3_33[5]}
   );
   gpc615_5 gpc1401 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10]},
      {stage2_35[6]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[2],stage3_35[3],stage3_34[5]}
   );
   gpc615_5 gpc1402 (
      {stage2_34[11], stage2_34[12], 1'b0, 1'b0, 1'b0},
      {stage2_35[7]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[3],stage3_35[4],stage3_34[6]}
   );
   gpc615_5 gpc1403 (
      {stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[4],stage3_35[5]}
   );
   gpc606_5 gpc1404 (
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4]}
   );
   gpc606_5 gpc1405 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc207_4 gpc1406 (
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6]},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[2],stage3_39[3],stage3_38[5]}
   );
   gpc207_4 gpc1407 (
      {stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage2_40[2], stage2_40[3]},
      {stage3_41[3],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc207_4 gpc1408 (
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_40[4], stage2_40[5]},
      {stage3_41[4],stage3_40[4],stage3_39[5],stage3_38[7]}
   );
   gpc606_5 gpc1409 (
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[0],stage3_42[0],stage3_41[5],stage3_40[5]}
   );
   gpc135_4 gpc1410 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4]},
      {stage2_42[6], stage2_42[7], stage2_42[8]},
      {stage2_43[0]},
      {stage3_44[1],stage3_43[1],stage3_42[1],stage3_41[6]}
   );
   gpc135_4 gpc1411 (
      {stage2_41[5], stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9]},
      {stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage2_43[1]},
      {stage3_44[2],stage3_43[2],stage3_42[2],stage3_41[7]}
   );
   gpc135_4 gpc1412 (
      {stage2_41[10], stage2_41[11], stage2_41[12], stage2_41[13], stage2_41[14]},
      {stage2_42[12], stage2_42[13], stage2_42[14]},
      {stage2_43[2]},
      {stage3_44[3],stage3_43[3],stage3_42[3],stage3_41[8]}
   );
   gpc615_5 gpc1413 (
      {stage2_43[3], stage2_43[4], stage2_43[5], stage2_43[6], stage2_43[7]},
      {stage2_44[0]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[4]}
   );
   gpc615_5 gpc1414 (
      {stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11], stage2_43[12]},
      {stage2_44[1]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[5]}
   );
   gpc606_5 gpc1415 (
      {stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5], stage2_44[6], stage2_44[7]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[2],stage3_46[2],stage3_45[2],stage3_44[6]}
   );
   gpc1163_5 gpc1416 (
      {stage2_46[6], stage2_46[7], stage2_46[8]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[0],stage3_48[1],stage3_47[3],stage3_46[3]}
   );
   gpc1325_5 gpc1417 (
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10]},
      {stage2_48[1], stage2_48[2]},
      {stage2_49[1], stage2_49[2], stage2_49[3]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[1],stage3_49[1],stage3_48[2],stage3_47[4]}
   );
   gpc1325_5 gpc1418 (
      {stage2_47[11], stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15]},
      {stage2_48[3], stage2_48[4]},
      {stage2_49[4], stage2_49[5], stage2_49[6]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[2],stage3_49[2],stage3_48[3],stage3_47[5]}
   );
   gpc1406_5 gpc1419 (
      {stage2_48[5], stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[2],stage3_50[3],stage3_49[3],stage3_48[4]}
   );
   gpc1406_5 gpc1420 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9]},
      {stage2_51[1]},
      {stage3_52[1],stage3_51[3],stage3_50[4],stage3_49[4],stage3_48[5]}
   );
   gpc615_5 gpc1421 (
      {stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], 1'b0},
      {stage2_50[10]},
      {stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7]},
      {stage3_53[0],stage3_52[2],stage3_51[4],stage3_50[5],stage3_49[5]}
   );
   gpc615_5 gpc1422 (
      {stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[1],stage3_52[3],stage3_51[5]}
   );
   gpc615_5 gpc1423 (
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage2_53[6]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[1],stage3_54[1],stage3_53[2],stage3_52[4]}
   );
   gpc615_5 gpc1424 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10]},
      {stage2_53[7]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[2],stage3_54[2],stage3_53[3],stage3_52[5]}
   );
   gpc615_5 gpc1425 (
      {stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11], stage2_53[12]},
      {stage2_54[12]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[2],stage3_55[3],stage3_54[3],stage3_53[4]}
   );
   gpc615_5 gpc1426 (
      {stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage2_54[13]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[3],stage3_55[4],stage3_54[4],stage3_53[5]}
   );
   gpc615_5 gpc1427 (
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[2],stage3_56[4]}
   );
   gpc615_5 gpc1428 (
      {stage2_56[5], stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[3],stage3_56[5]}
   );
   gpc615_5 gpc1429 (
      {stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6]},
      {stage2_58[12]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[4]}
   );
   gpc615_5 gpc1430 (
      {stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage2_58[13]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[5]}
   );
   gpc615_5 gpc1431 (
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16]},
      {stage2_60[0]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[0],stage3_61[2],stage3_60[4],stage3_59[4]}
   );
   gpc615_5 gpc1432 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_61[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[1],stage3_62[1],stage3_61[3],stage3_60[5]}
   );
   gpc606_5 gpc1433 (
      {stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[1],stage3_63[2],stage3_62[2],stage3_61[4]}
   );
   gpc606_5 gpc1434 (
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[2],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1435 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[3],stage3_63[4]}
   );
   gpc1406_5 gpc1436 (
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], 1'b0},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3]},
      {stage2_67[0]},
      {stage3_68[0],stage3_67[1],stage3_66[2],stage3_65[3],stage3_64[4]}
   );
   gpc1_1 gpc1437 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc1438 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1439 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1440 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1441 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1442 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1443 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc1444 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1445 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1446 (
      {stage2_3[11]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1447 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1448 (
      {stage2_7[15]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1449 (
      {stage2_7[16]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1450 (
      {stage2_7[17]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1451 (
      {stage2_7[18]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1452 (
      {stage2_7[19]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1453 (
      {stage2_8[19]},
      {stage3_8[8]}
   );
   gpc1_1 gpc1454 (
      {stage2_9[6]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1455 (
      {stage2_9[7]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1456 (
      {stage2_9[8]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1457 (
      {stage2_9[9]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1458 (
      {stage2_9[10]},
      {stage3_9[11]}
   );
   gpc1_1 gpc1459 (
      {stage2_11[14]},
      {stage3_11[7]}
   );
   gpc1_1 gpc1460 (
      {stage2_11[15]},
      {stage3_11[8]}
   );
   gpc1_1 gpc1461 (
      {stage2_13[6]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1462 (
      {stage2_13[7]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1463 (
      {stage2_13[8]},
      {stage3_13[8]}
   );
   gpc1_1 gpc1464 (
      {stage2_15[18]},
      {stage3_15[6]}
   );
   gpc1_1 gpc1465 (
      {stage2_15[19]},
      {stage3_15[7]}
   );
   gpc1_1 gpc1466 (
      {stage2_15[20]},
      {stage3_15[8]}
   );
   gpc1_1 gpc1467 (
      {stage2_16[14]},
      {stage3_16[6]}
   );
   gpc1_1 gpc1468 (
      {stage2_16[15]},
      {stage3_16[7]}
   );
   gpc1_1 gpc1469 (
      {stage2_18[15]},
      {stage3_18[9]}
   );
   gpc1_1 gpc1470 (
      {stage2_18[16]},
      {stage3_18[10]}
   );
   gpc1_1 gpc1471 (
      {stage2_18[17]},
      {stage3_18[11]}
   );
   gpc1_1 gpc1472 (
      {stage2_18[18]},
      {stage3_18[12]}
   );
   gpc1_1 gpc1473 (
      {stage2_21[12]},
      {stage3_21[8]}
   );
   gpc1_1 gpc1474 (
      {stage2_23[13]},
      {stage3_23[4]}
   );
   gpc1_1 gpc1475 (
      {stage2_23[14]},
      {stage3_23[5]}
   );
   gpc1_1 gpc1476 (
      {stage2_23[15]},
      {stage3_23[6]}
   );
   gpc1_1 gpc1477 (
      {stage2_23[16]},
      {stage3_23[7]}
   );
   gpc1_1 gpc1478 (
      {stage2_24[12]},
      {stage3_24[5]}
   );
   gpc1_1 gpc1479 (
      {stage2_24[13]},
      {stage3_24[6]}
   );
   gpc1_1 gpc1480 (
      {stage2_25[12]},
      {stage3_25[6]}
   );
   gpc1_1 gpc1481 (
      {stage2_25[13]},
      {stage3_25[7]}
   );
   gpc1_1 gpc1482 (
      {stage2_33[12]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1483 (
      {stage2_33[13]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1484 (
      {stage2_33[14]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1485 (
      {stage2_33[15]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1486 (
      {stage2_33[16]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1487 (
      {stage2_33[17]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1488 (
      {stage2_33[18]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1489 (
      {stage2_33[19]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1490 (
      {stage2_33[20]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1491 (
      {stage2_33[21]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1492 (
      {stage2_33[22]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1493 (
      {stage2_36[13]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1494 (
      {stage2_36[14]},
      {stage3_36[6]}
   );
   gpc1_1 gpc1495 (
      {stage2_36[15]},
      {stage3_36[7]}
   );
   gpc1_1 gpc1496 (
      {stage2_36[16]},
      {stage3_36[8]}
   );
   gpc1_1 gpc1497 (
      {stage2_36[17]},
      {stage3_36[9]}
   );
   gpc1_1 gpc1498 (
      {stage2_38[21]},
      {stage3_38[8]}
   );
   gpc1_1 gpc1499 (
      {stage2_38[22]},
      {stage3_38[9]}
   );
   gpc1_1 gpc1500 (
      {stage2_38[23]},
      {stage3_38[10]}
   );
   gpc1_1 gpc1501 (
      {stage2_39[12]},
      {stage3_39[6]}
   );
   gpc1_1 gpc1502 (
      {stage2_41[15]},
      {stage3_41[9]}
   );
   gpc1_1 gpc1503 (
      {stage2_41[16]},
      {stage3_41[10]}
   );
   gpc1_1 gpc1504 (
      {stage2_41[17]},
      {stage3_41[11]}
   );
   gpc1_1 gpc1505 (
      {stage2_41[18]},
      {stage3_41[12]}
   );
   gpc1_1 gpc1506 (
      {stage2_41[19]},
      {stage3_41[13]}
   );
   gpc1_1 gpc1507 (
      {stage2_44[8]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1508 (
      {stage2_44[9]},
      {stage3_44[8]}
   );
   gpc1_1 gpc1509 (
      {stage2_44[10]},
      {stage3_44[9]}
   );
   gpc1_1 gpc1510 (
      {stage2_44[11]},
      {stage3_44[10]}
   );
   gpc1_1 gpc1511 (
      {stage2_44[12]},
      {stage3_44[11]}
   );
   gpc1_1 gpc1512 (
      {stage2_44[13]},
      {stage3_44[12]}
   );
   gpc1_1 gpc1513 (
      {stage2_44[14]},
      {stage3_44[13]}
   );
   gpc1_1 gpc1514 (
      {stage2_44[15]},
      {stage3_44[14]}
   );
   gpc1_1 gpc1515 (
      {stage2_44[16]},
      {stage3_44[15]}
   );
   gpc1_1 gpc1516 (
      {stage2_44[17]},
      {stage3_44[16]}
   );
   gpc1_1 gpc1517 (
      {stage2_45[12]},
      {stage3_45[3]}
   );
   gpc1_1 gpc1518 (
      {stage2_45[13]},
      {stage3_45[4]}
   );
   gpc1_1 gpc1519 (
      {stage2_46[9]},
      {stage3_46[4]}
   );
   gpc1_1 gpc1520 (
      {stage2_46[10]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1521 (
      {stage2_46[11]},
      {stage3_46[6]}
   );
   gpc1_1 gpc1522 (
      {stage2_47[16]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1523 (
      {stage2_47[17]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1524 (
      {stage2_47[18]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1525 (
      {stage2_50[11]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1526 (
      {stage2_51[13]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1527 (
      {stage2_51[14]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1528 (
      {stage2_51[15]},
      {stage3_51[8]}
   );
   gpc1_1 gpc1529 (
      {stage2_52[11]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1530 (
      {stage2_54[14]},
      {stage3_54[5]}
   );
   gpc1_1 gpc1531 (
      {stage2_55[12]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1532 (
      {stage2_55[13]},
      {stage3_55[6]}
   );
   gpc1_1 gpc1533 (
      {stage2_55[14]},
      {stage3_55[7]}
   );
   gpc1_1 gpc1534 (
      {stage2_55[15]},
      {stage3_55[8]}
   );
   gpc1_1 gpc1535 (
      {stage2_55[16]},
      {stage3_55[9]}
   );
   gpc1_1 gpc1536 (
      {stage2_57[12]},
      {stage3_57[6]}
   );
   gpc1_1 gpc1537 (
      {stage2_57[13]},
      {stage3_57[7]}
   );
   gpc1_1 gpc1538 (
      {stage2_58[14]},
      {stage3_58[4]}
   );
   gpc1_1 gpc1539 (
      {stage2_58[15]},
      {stage3_58[5]}
   );
   gpc1_1 gpc1540 (
      {stage2_58[16]},
      {stage3_58[6]}
   );
   gpc1_1 gpc1541 (
      {stage2_58[17]},
      {stage3_58[7]}
   );
   gpc1_1 gpc1542 (
      {stage2_59[17]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1543 (
      {stage2_59[18]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1544 (
      {stage2_59[19]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1545 (
      {stage2_60[6]},
      {stage3_60[6]}
   );
   gpc1_1 gpc1546 (
      {stage2_60[7]},
      {stage3_60[7]}
   );
   gpc1_1 gpc1547 (
      {stage2_60[8]},
      {stage3_60[8]}
   );
   gpc1_1 gpc1548 (
      {stage2_60[9]},
      {stage3_60[9]}
   );
   gpc1_1 gpc1549 (
      {stage2_60[10]},
      {stage3_60[10]}
   );
   gpc1_1 gpc1550 (
      {stage2_60[11]},
      {stage3_60[11]}
   );
   gpc1_1 gpc1551 (
      {stage2_60[12]},
      {stage3_60[12]}
   );
   gpc1_1 gpc1552 (
      {stage2_60[13]},
      {stage3_60[13]}
   );
   gpc1_1 gpc1553 (
      {stage2_61[13]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1554 (
      {stage2_61[14]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1555 (
      {stage2_62[12]},
      {stage3_62[4]}
   );
   gpc1_1 gpc1556 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1557 (
      {stage2_65[6]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1558 (
      {stage2_65[7]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1559 (
      {stage2_67[1]},
      {stage3_67[2]}
   );
   gpc135_4 gpc1560 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[0]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1325_5 gpc1561 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[1]}
   );
   gpc1163_5 gpc1562 (
      {stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[1]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc1563 (
      {stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc1564 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1565 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc207_4 gpc1566 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1567 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4]},
      {stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3]}
   );
   gpc135_4 gpc1568 (
      {stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], 1'b0},
      {stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[1]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4]}
   );
   gpc117_4 gpc1569 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc7_3 gpc1570 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], 1'b0},
      {stage4_16[1],stage4_15[1],stage4_14[3]}
   );
   gpc117_4 gpc1571 (
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7]},
      {stage3_16[0]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[2],stage4_15[2]}
   );
   gpc606_5 gpc1572 (
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1],stage4_16[3]}
   );
   gpc606_5 gpc1573 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[2]}
   );
   gpc117_4 gpc1574 (
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage3_19[6]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[2],stage4_19[2],stage4_18[3]}
   );
   gpc606_5 gpc1575 (
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5], 1'b0},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[3]}
   );
   gpc215_4 gpc1576 (
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4]},
      {stage3_22[6]},
      {stage3_23[0], stage3_23[1]},
      {stage4_24[1],stage4_23[1],stage4_22[1],stage4_21[3]}
   );
   gpc615_5 gpc1577 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[2]}
   );
   gpc606_5 gpc1578 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[1],stage4_26[1],stage4_25[1],stage4_24[3]}
   );
   gpc606_5 gpc1579 (
      {stage3_25[6], stage3_25[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[1],stage4_27[2],stage4_26[2],stage4_25[2]}
   );
   gpc2135_5 gpc1580 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[2]}
   );
   gpc2135_5 gpc1581 (
      {stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8], 1'b0},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[2],stage4_28[3]}
   );
   gpc1343_5 gpc1582 (
      {stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc7_3 gpc1583 (
      {stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5], stage3_32[6], 1'b0},
      {stage4_34[0],stage4_33[1],stage4_32[3]}
   );
   gpc2135_5 gpc1584 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[2]}
   );
   gpc2135_5 gpc1585 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[3]}
   );
   gpc606_5 gpc1586 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15]},
      {stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5], 1'b0, 1'b0},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1587 (
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3],stage4_36[3]}
   );
   gpc606_5 gpc1588 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[1],stage4_39[1],stage4_38[1],stage4_37[4]}
   );
   gpc615_5 gpc1589 (
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10]},
      {stage3_39[6]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[1],stage4_40[2],stage4_39[2],stage4_38[2]}
   );
   gpc207_4 gpc1590 (
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[1],stage4_41[2]}
   );
   gpc207_4 gpc1591 (
      {stage3_41[7], stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[2],stage4_41[3]}
   );
   gpc615_5 gpc1592 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], 1'b0},
      {stage3_43[4]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[3]}
   );
   gpc2135_5 gpc1593 (
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10]},
      {stage3_45[0], stage3_45[1], stage3_45[2]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc2135_5 gpc1594 (
      {stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage3_45[3], stage3_45[4], 1'b0},
      {stage3_46[1]},
      {stage3_47[2], stage3_47[3]},
      {stage4_48[1],stage4_47[1],stage4_46[2],stage4_45[2],stage4_44[4]}
   );
   gpc615_5 gpc1595 (
      {stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_47[4]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[2],stage4_47[2],stage4_46[3]}
   );
   gpc1406_5 gpc1596 (
      {stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8], 1'b0, 1'b0},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3]},
      {stage3_50[0]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[3],stage4_47[3]}
   );
   gpc615_5 gpc1597 (
      {stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[0],stage4_51[1],stage4_50[2]}
   );
   gpc615_5 gpc1598 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage3_52[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[1],stage4_51[2]}
   );
   gpc606_5 gpc1599 (
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[0],stage4_55[1],stage4_54[2]}
   );
   gpc606_5 gpc1600 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[1],stage4_55[2]}
   );
   gpc615_5 gpc1601 (
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4]},
      {stage3_59[0]},
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage4_62[0],stage4_61[0],stage4_60[0],stage4_59[1],stage4_58[2]}
   );
   gpc7_3 gpc1602 (
      {stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7]},
      {stage4_61[1],stage4_60[1],stage4_59[2]}
   );
   gpc615_5 gpc1603 (
      {stage3_60[6], stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10]},
      {stage3_61[0]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], 1'b0},
      {stage4_64[0],stage4_63[0],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc615_5 gpc1604 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {1'b0},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[1],stage4_63[1],stage4_62[2],stage4_61[3]}
   );
   gpc1325_5 gpc1605 (
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4]},
      {stage3_66[0], stage3_66[1]},
      {stage3_67[0], stage3_67[1], stage3_67[2]},
      {stage3_68[0]},
      {stage4_69[0],stage4_68[0],stage4_67[0],stage4_66[0],stage4_65[1]}
   );
   gpc1_1 gpc1606 (
      {stage3_0[5]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1607 (
      {stage3_1[3]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1608 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc1609 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1610 (
      {stage3_4[5]},
      {stage4_4[2]}
   );
   gpc1_1 gpc1611 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1612 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc1613 (
      {stage3_15[8]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1614 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc1615 (
      {stage3_21[5]},
      {stage4_21[4]}
   );
   gpc1_1 gpc1616 (
      {stage3_21[6]},
      {stage4_21[5]}
   );
   gpc1_1 gpc1617 (
      {stage3_21[7]},
      {stage4_21[6]}
   );
   gpc1_1 gpc1618 (
      {stage3_21[8]},
      {stage4_21[7]}
   );
   gpc1_1 gpc1619 (
      {stage3_23[7]},
      {stage4_23[3]}
   );
   gpc1_1 gpc1620 (
      {stage3_26[6]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1621 (
      {stage3_27[6]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1622 (
      {stage3_33[16]},
      {stage4_33[5]}
   );
   gpc1_1 gpc1623 (
      {stage3_34[6]},
      {stage4_34[4]}
   );
   gpc1_1 gpc1624 (
      {stage3_43[5]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1625 (
      {stage3_44[16]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1626 (
      {stage3_49[4]},
      {stage4_49[2]}
   );
   gpc1_1 gpc1627 (
      {stage3_49[5]},
      {stage4_49[3]}
   );
   gpc1_1 gpc1628 (
      {stage3_50[6]},
      {stage4_50[3]}
   );
   gpc1_1 gpc1629 (
      {stage3_51[6]},
      {stage4_51[3]}
   );
   gpc1_1 gpc1630 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1631 (
      {stage3_51[8]},
      {stage4_51[5]}
   );
   gpc1_1 gpc1632 (
      {stage3_55[6]},
      {stage4_55[3]}
   );
   gpc1_1 gpc1633 (
      {stage3_55[7]},
      {stage4_55[4]}
   );
   gpc1_1 gpc1634 (
      {stage3_55[8]},
      {stage4_55[5]}
   );
   gpc1_1 gpc1635 (
      {stage3_55[9]},
      {stage4_55[6]}
   );
   gpc1_1 gpc1636 (
      {stage3_57[6]},
      {stage4_57[2]}
   );
   gpc1_1 gpc1637 (
      {stage3_57[7]},
      {stage4_57[3]}
   );
   gpc1_1 gpc1638 (
      {stage3_58[5]},
      {stage4_58[3]}
   );
   gpc1_1 gpc1639 (
      {stage3_58[6]},
      {stage4_58[4]}
   );
   gpc1_1 gpc1640 (
      {stage3_58[7]},
      {stage4_58[5]}
   );
   gpc1_1 gpc1641 (
      {stage3_60[11]},
      {stage4_60[3]}
   );
   gpc1_1 gpc1642 (
      {stage3_60[12]},
      {stage4_60[4]}
   );
   gpc1_1 gpc1643 (
      {stage3_60[13]},
      {stage4_60[5]}
   );
   gpc1_1 gpc1644 (
      {stage3_61[6]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1645 (
      {stage3_64[0]},
      {stage4_64[2]}
   );
   gpc1_1 gpc1646 (
      {stage3_64[1]},
      {stage4_64[3]}
   );
   gpc1_1 gpc1647 (
      {stage3_64[2]},
      {stage4_64[4]}
   );
   gpc1_1 gpc1648 (
      {stage3_64[3]},
      {stage4_64[5]}
   );
   gpc1_1 gpc1649 (
      {stage3_64[4]},
      {stage4_64[6]}
   );
   gpc1_1 gpc1650 (
      {stage3_65[5]},
      {stage4_65[2]}
   );
   gpc1_1 gpc1651 (
      {stage3_66[2]},
      {stage4_66[1]}
   );
   gpc1343_5 gpc1652 (
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0], stage4_3[1], 1'b0, 1'b0},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc623_5 gpc1653 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], 1'b0},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1]}
   );
   gpc3_2 gpc1654 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage5_8[1],stage5_7[1]}
   );
   gpc1343_5 gpc1655 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1423_5 gpc1656 (
      {stage4_11[3], stage4_11[4], 1'b0},
      {stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1343_5 gpc1657 (
      {stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc1658 (
      {stage4_16[3], stage4_16[4], 1'b0},
      {stage4_17[1], stage4_17[2]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc1659 (
      {stage4_19[1], stage4_19[2], 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc615_5 gpc1660 (
      {stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6], stage4_21[7]},
      {stage4_22[1]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], 1'b0, 1'b0},
      {stage5_25[0],stage5_24[0],stage5_23[1],stage5_22[1],stage5_21[1]}
   );
   gpc135_4 gpc1661 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc1343_5 gpc1662 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1], stage4_28[2]},
      {stage4_29[0]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[1],stage5_26[1]}
   );
   gpc135_4 gpc1663 (
      {stage4_29[1], stage4_29[2], stage4_29[3], 1'b0, 1'b0},
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[1]}
   );
   gpc1343_5 gpc1664 (
      {stage4_31[1], stage4_31[2], 1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0], stage4_33[1], stage4_33[2]},
      {stage4_34[0]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[1],stage5_31[1]}
   );
   gpc1343_5 gpc1665 (
      {stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[1],stage5_33[1]}
   );
   gpc1163_5 gpc1666 (
      {stage4_36[1], stage4_36[2], stage4_36[3]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], 1'b0},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc1423_5 gpc1667 (
      {stage4_38[1], stage4_38[2], 1'b0},
      {stage4_39[1], stage4_39[2]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1668 (
      {stage4_41[1], stage4_41[2], stage4_41[3]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3]},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1669 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1670 (
      {stage4_46[1], stage4_46[2], stage4_46[3]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1163_5 gpc1671 (
      {stage4_49[1], stage4_49[2], stage4_49[3]},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], 1'b0, 1'b0},
      {stage4_51[0]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc215_4 gpc1672 (
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5]},
      {stage4_52[1]},
      {stage4_53[0], stage4_53[1]},
      {stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc3_2 gpc1673 (
      {stage4_54[0], stage4_54[1], stage4_54[2]},
      {stage5_55[0],stage5_54[1]}
   );
   gpc7_3 gpc1674 (
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5], stage4_55[6]},
      {stage5_57[0],stage5_56[0],stage5_55[1]}
   );
   gpc1343_5 gpc1675 (
      {stage4_56[0], stage4_56[1], 1'b0},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3]},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[0],stage5_57[1],stage5_56[1]}
   );
   gpc623_5 gpc1676 (
      {stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage4_59[1], stage4_59[2]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[1]}
   );
   gpc2135_5 gpc1677 (
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc2135_5 gpc1678 (
      {stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2]},
      {stage4_66[0]},
      {stage4_67[0], 1'b0},
      {stage5_68[0],stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1]}
   );
   gpc1_1 gpc1679 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1680 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1681 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1682 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1683 (
      {stage4_4[3]},
      {stage5_4[1]}
   );
   gpc1_1 gpc1684 (
      {stage4_5[1]},
      {stage5_5[1]}
   );
   gpc1_1 gpc1685 (
      {stage4_28[3]},
      {stage5_28[1]}
   );
   gpc1_1 gpc1686 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1687 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
   gpc1_1 gpc1688 (
      {stage4_63[1]},
      {stage5_63[1]}
   );
   gpc1_1 gpc1689 (
      {stage4_66[1]},
      {stage5_66[1]}
   );
   gpc1_1 gpc1690 (
      {stage4_68[0]},
      {stage5_68[1]}
   );
   gpc1_1 gpc1691 (
      {stage4_69[0]},
      {stage5_69[0]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor_CLA64_64 compressor_CLA64_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hae93cab343848eacf9a9ec52f8f3b1069b2203a2a36adb12cfd7e049da1f853e46a027ef51f05349b9deb4b8294017b71880934784a90320feebee51f24d6607638d3b0d01851d3c0f9cf73042b61b749f841f6a050d2ecf5515f82ad16943dca7dfac95a909dd28470cc40c8202286afbebdea8cd50935597d0efcd737bd627610d358ae35ac00989ee824282fd967946a5d0938d8268f8c189f8a9fadee89db028ea986f322a30b49842ac8eeec5c73c397d901e07914121b1feab44b83914c66fdd4776e928ad40ba39b256af9d372d5363f760db08e7803f7da4020d9f8676f6e1b455892780be6467e27e20493cdd390bfe53ca6cf0f7513f3e7e3aa5cdd3d2a2d80ccd1409359ef874a0c501f80ee399b93c2858c00a2183e15b0847c472600c6ead4646083bc2d5e4c698841bcdf5669a5609e76be927a789005c5ed868df3e59cd296f5383daa75ef1b1fe7209f3a8b9aa526a39959e2c84b7145286e1e20027487d62539d2d998cdb39d087643be1be93329f4a783aea5c5ffd34da61950361fd4e227e8e49f6ab54ff08642d083c5fe8ed8a1ec5bf97fb88842b1b3aa9ca3aefc7eff66102fd20c3d703d940e227e173329d53c45c5bb1a165f0ce09ddec9dfaff332dfd9cfb46a57f6f3432c47b2665cbcb7f0b0753722ba7b9e8007a291090814a9682bf2e2a125555c4652c32e173126bcac4a8fbf96b917df6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hef89032916406d32ad6c99b4517808b0ed4818ddc9cc43a847ba6b6da5f5e5835d4b1c606767b1ad9e8eb73a177c948b6554336f9bc482056006323ed72e4c06f376fb7abd8e46934f7bd1b8f96bc2aadcde3e273ae7b0ccabf5f65b8c85387b234468acefab59ffa3272292d4f9ef66929b85dbc2625971dd0830ec91e524389092fc362b07be590b0ea9bb5a3478e7af3afce24a40efe6e37ce1149003af88dc4e4ffd987b086724bb376df567c7fcd4a977e68fa06a0e3fa759fe6f5dcff3b26835432f451d1b7b2a9688966aba4b37c90c746f335faa0531f1d8e1240afc2203533cbf2118380b929308943115060757c79dd8a127bd7bb0a800987f7a5340a3fb2bfdafbc325a9fd94f834dd10187a2d2170dd6604196907fc9b38048d520e0d7166af1f05802bb1d2b00430fb053e1b598b45c6b8bf86f451a304db97feda36d2902561d36374e5be4835c3ed15814a7faf21f1ea715ecaae1d0fc66e80072700dcd8c6b099b63ff1045422b083996fe559cf24f8a5165b56b04d424d137f8d3a05ae4dcc798346557bdffe503ccb25db2e48c643bcbeb455deced92a9855fa1d568bc500db61c303454f2a5a7f8936ae30606f80026f352c2d0206822088e21b2e75e7067d5538b5487c652a7b622a74c6edfac7110f3e658f124cf186ba68a309092e7d9c7c3255a845ef414970446f81389ed4befbaf85f537a510c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h39a1e0b1c469ca727f200178f686392b180ac595e2862350f8e8fbe60e05bc8879416b0762ac96292d71e556c6d7b5acaffc199a67fa77d5efc61ad8ad76c38410cad7bafbe3e840ba400ce20e3faaee6cf7467e54c0633dca5fd2d64008a7fdc1f006bbd8380cd7fc88672a13a69985390d8378c3992a977068ef4b10a4982f327c3fe5edf9b4067fcb5e65e28a7b114e22d985de52b38bcc48f6b30483cda2263bb1c543d1ed251c77da788d75ea1698d7610237d16f0a9e8f22c4791e9645a6f15bbacd8911289b49cd65546910bd2b3790ea64688a6267d2658783e1ccb13a947f63fe584dd29d517aab4ef98e0a983667794440d9c803bbac99844a60de706629ec58faa5cb654642759bc74dc9bb06cf9e4262ac28f6faeb5e644078f0bf79a995ea2bace4306d4701c87bfd8fe3b447488ba71e5e595d8bc9443b753120e72f1bec43cde11d5f80815ff0007a2688dfcb2066e6b093f348949f8a8dab5850b78f94be03d98cab9a7740b4245f2df44e84fbb2b1767f1cee9277f234a5b3efc89fbcc8fbab36ea0fe2e3358d59ab23773811b78a311f71df766b27b342ea43e2bb76ade0bcc4b73a36f723a7d559c067e896ddc0f4c923e90d6b505d2fb04f00c38477363f31e9ab861c47a454f4e112682e7bacd68c787b974ae7fc7a3f6d0818358a7d42b8ebbcf34b455b5e2c59f25e3b0fae2c82297e63d19f7e75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb29ee3cfbcadfffdf70b50e45e3937c725874963e2325c3fe5a155261c3f46ca2c742b7cbadd9b4a1110ee4697bbac78f80de46c8e097d6f2e95fd940aa00fe9f415287691f01c6d1e8b59fc648f925c43b2b276733623a959ee8306de67507ba85c4ba6e46ce5f74d84f1b8a74fcb13089138080bab0347a049119c06ca7476b712cb3ab8d93c980b2f99225f672409d5d6b9dd9d4dd2cecc3402f98f8db900faea758384357a80209d6064bc0c4dc6eae02f37e122a868bcde554cd1edce4ee38c06fa8bae39996575da186a89dd5209feed6acb626f7f60d289ca225c6ab62a5a47feef9e839e9f198ca3ab115000a67a1eca431809b0a744f3015347a705e1cf82fcee71c0d744618e285fa7eacb5aaf0234e9a5d84782a948044e618f13d65842fe06c1660a489e15315036b1b67bc54bf0e18d05cee26514230d2b7b141587abea0b115853a1f80e576c18dbef0322f732bdf2626cf480c458c65efffbd89b45f46cdcc97f2e57c310785a41a83fee506c3680b8107a844b6d682c97949e9885e36a8a5d326cd2f3acee84d14b776561dc76b02358934663e80749f792e5fb1550d30ef846f61c4832d67556294ee703daad6565692b8dae4253a9f71059d5a7fd09a227d2da24c04d11ff9f750040d59c0dd4a1dfa32cecfee2740a7e9486cf950104c74ff04af2359f48ce87613a2b98c6161e89567cbcbf10b9fbf4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6fa939aeee10fc3e8216bd252a10d62695bddff1a2a21724ef9cf50389235e997a66cdbf14bb6f53c64b6d7da81e8156a322049fb61b081aac4d12444e54411afbad7d075fd6992c714d78a0c3fceb97a1c1c2e4b3231adb3acb9fb23f199ac9b8424039550d029dffcb89132f41bfede82a40ba2833ef55e798264d56fc1322c2f6967151b467ed8bf9cc47d43b4b77b7d1f6e8df48e6411fe01db940c01bbb230cc7e57bf4080dfb1446a6bdcd49351c7178aa6940915933b55468394e2eb3cc2fd9d9c5e64fd7e76d1cb49aa7058d8c506560771b2dbaf81017185170a4dbe6506b9e98da32cc119966c8fbce74c229919ffbe513ebf25a69ec95d6459d889c74a99ac2f1f0dc5fa8f553911dc9295612ff0c76c6df7e2b2a5ace6fa1ac07c9943953e9423cbad3cc6b409979b9d078c3f520d46583a7e99d67f07944285327fb6b96f78af0dd4bb9a634ed251ae01c8529f6293ef7bafcc00611b41fcc2ac8099cd37c88528f14a11cbbf9f04a566a2887e5dc0f364be565abfd993a370053cb53ba981bec4d15c9a53b4ec7da4a418eedbe3f430ed18a3a878022de69455dbfbeaedee2c7accef102cedc85b607a69deb92251eeed4cb5d33aed4cf83bc944474838edbe58cb6d3e4939cc18580c0afe7fb837dd13dab659fed0f9c967f9570fd23e208e58dc58306f199110b1fde17d7234e3f9be6167eb29c06411018;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h43de6c6434647413932a720f3385d7f0be3dd2b5642cc03dde0d35568a664da673e4a08eebacb00bea27816959326bcc8198f5e7960bcb57a0bf5bba89827fc062c705356036039f34b859311469e868057f3f068c17437a745765726787bb2c7928059ca9c06910a26def4ee747aa8e7525ff9bb9c924a6efa8f2d56b0c1712eea1595b82f7a2f086f2c376d023290e7eef7f9b9fd0fcf3d9d17fcd746e46656b8ee5c6c8fb37d888beb2bde14756f378b2a21f98d262752e4f27e225d7a90be3bedeba51997b479704dafecb97c54d125ab97fe4258f091e4007fc12e90b4bc5392f72fc40a5add687d8508b0c10e9531012aac56b65bed48b697709636bad1d0e64f4702bd274de2d6e64f13e5f14d530c505862f6769f7568e4e518e4c609865b75dec068afb744e6ba673b999d4c458de8aff0dc739a528d5771054ff0e3db23e88c9cdc7393502d2c587dd97443ae5cbf85dda86bb19d818dfbd629b6c0b58022015c524606cab1b6e83dd910f61e16395e9543fea5b55c860f06446e467fd9e424310a97794c484c620fbd44b1b5251ecf89f97b5f927b76f22e2107622dda55fff92cd92808b8b0b491711fba2d0246a99cfbd7883ac4afba17e0f8d026770a80859fd60c3a93098adebfee273f5d42f7c75d967d3d7817b6023400f7291d333f4bb3f451c2dd0912ef4a69422290ccd3f8704e51d3c8d9543af7e4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf1678cf6c3302846504adaac5ee90cd3173aea96b0ee9fd2eb4524e4807014ea2cbb5669a07d33a7edb591e35130280558ae44ff1255352b5351a874230fa4bef04993192f84e21b46f11ec9957c2917b9dc073605c5e5416f8663ae0a2cdb400b76871ad289295b8964afffee3c63efccecfdb482671d182bbe91dc8050a2ec276eadd1b0e8e6d3395e3e0f59021458c3d8b7923cba62c50f0c93fe85e9044ba51649cdb890cb94a6ba5d49240c4905a98a3c6c4463e6396f813f1dd32f5d223079f3bd2c822102231f8ecac8aefd98ab95a82894ffbbe4107e2bcadbaac6220eb6516b2f90e2c024bfeef86e77e2df6d018c9ed89d907f0e5685e149a3c04dd9059454f9150c76370996f030f70f04f208f18c4a50f6b33d249c8ad3f623fa9a40c2e93584f40ad60bfd2f435407709d7d11d7db6e6e8a47929c7577c42e4584d3b84d66b3cf099a17d4704844b87e6d8065bca6073c44e309dfc66c423207417d3b8a02bfdd5e5117dcf29eb3e1a6a789c844857ca868bef2fa01fb896f491cfee4e3dd4691903e49ca1951da2736a4c5662186330a00d66bf30e4f1236f7312b8878fb7498c86a4c575e36cb19570491bf742e8dc3f9eec242853260e0b8644f03d6c66b31a2cf239d65b43709181a16cfd3cc847b071194e5f0630eeea957a9da0107f52570f15de6af3a1b045f20ee3fbe9b573f71c3c4b81db288b0de;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h82efe6702bd3b34c57ebf71114a27ffa956ea7c296e0ea121e0322e713b2ad1f68dadd13a6456462a59634bd6ba06d147d1b1fe49e36855c48b7b168e5d0c07d9778cac5d011f652b78876b7a5035d3e9abd82da3951f5d32d591b661ddd05f525286b48d46c97c3cb8eca3e2f4b5a455dfb056fd7d10d744407e9bdadb513bcfaee9186e0f3d76a4ca72babcf15fe1aae08a4496481fadb6f10228d8cde2d5cf5385d06237997e424483058737c248bc50f5d34133bc660cb3b54ae1a2582a4687ee59cce6ccbb028cf172364f663d9faf448d13a4aa59a2bceb15ef61334ca896bc4bfb3ff222591ebd494af8b1c2dac1afeae6bbcc4d9df3a4e6c15a0961a5d20d950da76712fd2ca31b87dd5689c9dcc32d396139dc92738ed16e0919b323b77001a0460ad6dd4ae9e5e578a86d22cf378da33e7a4ce9dc0b25531e0c52617b06250a2e172a4a92b6af665468a0e0b3f959a5afd1c6fd1db823d1f6978658f58b7eea7ddb45e09fcae7970242e395991993ecccf377037b94299a65cb077a485780be571d960e3208a7996671e48e27ee2fa6459441d7b0475bb9762cafef99bfca9deb12795a1ee683c93eae481228bf16a9babe7e43c592ac320332baae71af223912831639323b9d0e907943955ace0fcc6558fb650a01bd29792dbd45b632b4d4faa6360a37c103288b82348eb88a0d2d871afd8994b261041ad5bf4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5926e6bb340dead67174a1eeaf921d1b9e1483fd97efa546e2506984d56c88276fd10cd401f9cc2ceac5b7c6be1d18267850f0ad83ef23fccad62e3dd41895d74d7258fe3f1e63979be42cfad256c042d5b39fdf8ebe1fb626366aad365a19f7ef293401cef6e7e2b90bbbfcbf0eb23376d680192052f98f6ad8efb45b7fb0376a7b51a4915c09c6e243b3291a61deff7dc9ea1315644c0ee00087647a326195ea346d21e257d90a53fc1a92aa2dae27b9d69929ddc0a64a5cab26709bd1d39a68ce4c1bcd8b60aa2b6b541bd47dfe24683e1a87ed4e41334d029803e63e467451e845b1987ade7683dd829a2f5024c02eea7f241f17f81e7a1aea63e0747c2f8d01262a380ad271ab5bde684527176988a35520a694d4dc0fbb6d23531d58ddf2849fb66d2d11b7c4153b2589e6c1f8eafaadb0892f18bd93b7097e6ab2b91b0c672c7fa8c3e5d66b821db4caf1a89670108169fc364dc44213dc2048523e7d10ea87a52dd6d3dc33b59731d7563e91c4a45c3c31b5d8df84c37a7cc2fd1839cf8c5326102726504738e96511e4f1be4bdabcf46f25284be8e5aaf932b7a9093cfde9ba957ac79e8818014cbe8c1dca3fd7aec61bada91321869b235d5f977e4f26bc9060dd7e506dadc981f362696399b4986df628dfe65ea2d8174ec64adc422df5480eec985b3cb36796952c499f3e9cd85c060b93527a733cd5b3eb9218;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4521b51e2423702bb1f62378efb31a8d3c9ab2fc563659d26dee4a63c6d28cb103aa3dd5fb0f33a1fe10bc2f8b83f6654b6627ca19415df3db84543472407fc181b8abb7fd17feafa400ffabdeda9032259cf39e862b3a3613a5362f5dadad624af6624b63d4c3991143e386197bfcb3edb2ffd659a7a3055af1b017135b9bb6681866116ac7c0d64fb4e4b265a39de38c7d922d6d5a8a1b0c837fde324859132ccae619232f113b087e20b1a8082487610416bb0298f94231a87a8c0d5e75fba0c04ef01985f6a3e3c3786dac78b665b0f3bb4c46a4d354ec3a04588bc3baaaf6bf7154bc2cf1463004cfb53ed62b0d9e26722c4b158c0fa11f0cc55aa4e14c105d9bc3c2e68094a9a6ce1741acecd6f3208d095db769b7e1d4d28769512f2ec196ce624aa5f02dd00b08cb1e1c66c22e4c434dfd1e3a56bcbbd6a4f4ebb7b24766c9de6a17dbf3ae86761a3c94e209b79d5bf655c6ffd6acde3872b6082244f7e0d4180e16bbee80e57eaa4504243927a18562b17770fd49fc15f9dc67656918c95203d810ab5853a7f8e33e51336f30786338cfd3741bd829feb3f291a856cf3f8b4a601d5308a7e42fd0a55e03467ba38c1fbd53a94370a63d35454f04ca610ee25984150e639c0a6f70e8b8f4f5a27fff6f7ee1cb2c66b0854c58a3ffd08f3f2040c69387379feba8813d61134429b28d1da4beacad68a7ba3f42a71c9c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd9c03888367f8ce5be5bb392d5c3af211a1ed040d0b29fbf6b6ba98dd29afc2050de06e3bd232cb0603f5c9b470c702ed8a3f8dc11377460a7450e64c9822d42e84bb898696aa4df346a0a3cab21dc5cd3088b9a2245062ee071ee2477bc2d81f51b453b6de38425d1600712313575afbe0a0d4c42fe04ebbdb5888727a16555f708ae55d1e3943fb7875b9868bc0f22c9afe30400d889e0c2178709dacc4e065328df46f99312e8ee12e2a9fa375527bd84ca083409d99dcd4a6656758371867d1c9c3802312496a3743128bf6e147a332c58b9a5d18d68e0dd87538a7a3c9325f64098b41d1086cdf44ab65c229e1f5c0a00f8bfa3d4036f38b700ba9cacdb3324d788dfaa1edae2978160f02eb3fe069da7dd5b4b41632df4cafb8f7f80dc0be1b38cbbbedb8e9d149a79e59854e67ac9c4771f62d49f162f64d0650311896bfb7904d4787b75f6f0b7d7700aa9ae931147d69b68417e007f1bfcd3f2dddb8404134b390b87486866c65a350b12cf7185138e43759e3f52cefda6091a37d70eae8b3a032d92a27b7cfbef7306656984df8b8f93461af0f77c450e7eb32e3c48263cb8a4b14dd1d538f76b52dde64f432ec1f607cc793c2a5004b7c83b6d2f25ea4f21c9c156bb2c8f0fc09af2de75ca5bf9b05b02c712e40c7ec55f0beb48642ac215828447ed255beeaec554d0c03f6683ba4814c7fb5e1f559d9572785;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf03bc5e2b53db006c4f4482f3c43f87e69d595fef192bdc34be040fe5ec3dcbdd1cd2fbf0d33727015fe806de83ff872cc961f90b319cb2ef1e4ab3b8eb46fd2dd1b44c0d739307af085c70ed1f4c4345797b186871ccf3d967f0209dd9c0bcd347906ddae42b4dadf7b853fea47aecf21f703e73258a8c8a947f3858d7df0ad1cd47323eb6fafb8b94e406f8e299644a076ae081ba6c47f7e159ab18e02b28c94759381f0fc025e55dced9bd1d8bde7bde464897da3f325098f8c404736053c85801cfc73f5d6bb8fb6eea02219506843b3fb382e99d68d5dad7285ee67e3fc5393737c94463bf760f8b07e5676b033096b5bb063a63b77c34781e94fe866ce942f3eb8fba638ca31912feb81ac6ce98ebdd72be8cd64076d66ffac6fa8d65291b81ab9f6dcedf7a4ea88e71a23c16741668de9c0660436ef30bff6fc6baff60960041c4ca289fe3d7872357349ba2b9cb913017c4f251f230bc871f70107745a5c1d55952984330ee063c3270f0a0c531116b63d254d48f9e704a7a8acda33e8efba882fc0b0667ee12a57657b6f1b11ccb41b4a0ca09c31b142ecfe3f02c9eb2e7a388e4022c84dcc8c00f65c51a94113134b1abc0347d06042f95b063783154dcfb2bb036f825de0dbe174a4ed78fd9c8d445a69329cfc85d3f22e33ba40602717f9bfa212a981bf8164d96ea5861fc09e662add6a4b31d57dea3858b7ad;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4e4fc27d82678267dd9061c71cdae0a7cf25668cafd9ba7471f847f7e104d4e90f513a431ae7fd7fae66e7dc34f67ea518bff832ae78cadbaac03fd8f497125353575342b6563775668c5c8865d7e8f89d4960db76173b1f71e7823984b9bac5574ba6c0994ab33054e6c29359386ee51e7ecfc167c1a3f54df9c867ad7b264e8e3d21b5e35d4e53b43fc7e2e6c10d7086b35e9080e06e4a61f1d9bc8727b6a63102f69b6bf058d7810ea1badcebde45b58c337e8c0cbc44e26255d6768e89ba4e6c5e25ff133501c9769540979df3efb8d5928cfc282db18db19abb5a0047845c1e380614b8e287b9106b9e321929d1d6b541323d400594fe3fc0c06ff460cccad8786e5c9202e4a9661df9f9e0df91b67b527aa09e9ed1c46f75a97df14bab8dfb1256df4d2c16cc7d37a9905fc9434f7943ed9ae4367221cd96584e9811ca4b7fff49e47e4b6c48e84041b0cea9aa8f49c79b2d5a10d75d483abd5400cb24553523511ab494e16faf554e0eca222994f6bc5ec9d7fd79890271599eed43bdd133f7c97dffea2b05ca6cdcec1b58d410d3f69f8e2c16a764645aae6c6a29f31b08587fa317d99f5c7ea09c953f32e6a9f7f99331d6ee91b371217d64e6bf5c80d1dd4740aa7478c91b14af787bd90229bcda4ea899584f5e64f28dbf6aeeba2b77108264a333404bc1a9bc779e0dc0e49db77637af5aceede6da30134550ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7760404f7d63e7cf3b1bbae2cb0030bdeee34967a8bd4efe48a462a50feb9cc729c71e9b89666b7d713b9155ee1016704a496ef22b1438f92a20442c1b5bd407f7fad034d569f9a15321c9423594b08b577ab601eab5e32a05309a4e6865e45da1172630f6869476adc42cda02d8558d4d5e10975524bdf96e12c7d9b7e61a81e85187c749df345bf3f6c0dbdf7c819b20af8c549d5fcdee3e66b32573881881fda2961729ada9da1ffea19432400371c034ee7093134ce62be968c69f02e2a47b5042ae13ea8b9ecc04849a38680538d0b0614006308a6967a875940dd8732f332a109223177bc7f5887ac213e8d0e3ad50a5a46d7ff14332e9b2bf6fc3bcae3dc44ef5429daade2be7d7db0fb6877c29398ddd6eb129c2f6a26f1c491494b745836f0db031a0a8b891c038122760bdef4524edcca3f0964cd1c3abbac0eee2c44c2451c9a45c352d9d3b596340137feac8da6fd90e424711a3ddff24b0b6edda16c8abc0d1c918c644dc352e8c96089a2c5d0a5b67dbc7677412a76a653f23a2990506635eca1bc4b82e580f9afcd1251f2ab28c7e5eeb48c477706689db79489e7b78d6913e3f2dd15d788edbf5718b28bb5e15a4308b79ab6294f83c6898cb9617744dc9a4bc09258c2f4124a8be10d072bd4936964ecb7a43b77ddd187868148ae9b4512afc95bee361440edf11006ab8d974f67aa1715c49e4c5cf5811;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h34c129d9b45de72eeae6b6f1cee1b83500872541343532e669c7830f6e7f7208bc30e02145f2632382c2ffee532716cb23bc08bef499904973d557841d71d59ef5887ae3910460b4179bfe11533eb88afb185fb26d180aa98476026d698b7ec7723998433602572aa75eaedc2cb882ea9262608669f3abf2a2b1a0ee9ceebe62163c8630ce883452e6f7a93969c103385cc23eb9508778e2d3cfa275917d92cec3a1eec6ab4f95fb3f3958b2af84761c778ec9704211c1287886e24a2aec65106bae1a14d8270a526958d4dce1d2ab3aff6de362c0e96da6ec6935580ba6031d85b19994e1325b9379301ad163f49c9cd7d31e4934dec616d9ada10beaa5e9f1bb59cb6e6ec9f3c12b891d4aabbce94b94486c630a346506ad86dabd3398b1f6cdd9ddd3ecf8d3a534b234b0933b01f12d6a707d1fb5944d41b48473ec34cdba866832644df94a73b1f4b6926b10dbadf3aae0a8f16db3be21f27039d9a74aeb52cea959d072006297729e74d38d643e164b1ad455342a61bfa0432feb4363e69d9911b6faca4dfb114b4cfa879242df5444dadfe4bedcf0f7949ee0d8081faa84e7cfd00cf99a0f4d9f6fef98a24284b4edea0442b8843011bd4e770c27d8943d5a16c6c3c36caa7dd269db7f06323af47bde548836f64ad6bd5d0cae65ea7f73fd4040bef7d63be9966ddca4d905b658bb0704d7702a87e717d647006176ce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h697c9163efa8c8a61f2e8077da241dc65656dce285915ffcf46ef55b79d40c702a8805ed25cbf8c7493e814d782068559c2f80ea7edca98c331e4d2ad000e4fc7f5b9de3c57eefcc26bafd7f1a65d23a995bc82864c321bb6963c3110d5b4434e7ba165ee59e6299891bb4699d7031143a291cc2753c3a16255267930e64ab90fce714eeef3686de8b7beef028f8265cd1b09ed5d2b95fddb718bff10af92cc74c4fce601fe1c287bcb43d610e89343f4dded7009b945e942e0d0c731a39f46146c3c932c070e7707c0696eb61ac29527c0e8a273ac200cb95cd31f52f58b7d225be9aa6a11651c0815613243ddf9d35cb0315eacebae675f5c1f446b8a261c20aadb4b8be14d32b07373b38ced570acdd6a3232c6519b104d7f6cf28c2b7ed617d5b1a2049932bab016a30ee11a606e23337ed02eee69bca3f0ef1d0317bf0530bcc76b8deeafb738a00436a509dd28a7a8e3da12d6ca180dbe676677beff2fc2b693a833344dac2720d3da99290aa070c64c5e2733bd15ceef4b07310de0ae8bfa48604927755cb30c5fc391db90325c4d6be0c30e9301eb327b553a050807b650320c78aeea42a9bd28c5cce1b002dbf219db686e7ade830b40b8537b78290f90614584fbc127c68ca7b55fc5a3251e9d0e055fc9b2696994bc741e3614a1a057c74774707adacadd3a610fc8d1f586956bfb823f319f10061d02e422954d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h60437341f6bf6b847f4eae4c1e8ef58b42c6ec308a1c9c27ca406523ddc1bb4ee37fc46e05d14ae08dac39e4495e40ad945c4ebfab358a201f11f0cfc57f4fe1a95f3e8ec09d3b10b5e471ecfdb8521cee7757bfaf64955d39b17049f19eb75e646d325cc7ae012de0997cd3718ba53318c872b51fa2f5f96d96f69271e661ba51525c464831c38819115787719a38e4a2c290a609d484798ab6787851363b59bc63c25b3427be98142c31c438d46ce0d2c046fff5543658f6a7a72b3d528fadcbbf754fcfe229d3d5f6e897295c4228d35d79bda745c829e8d1d30cdabe282093194713920e09e8abe184eb1f447876210b292c774cf2affe2e1a36e08cb2497483066c50fad88c34183e0032b71b47016d0bbfd4ab18a9fbb3166b9f14b880314185b664c7a5497ce090d95cfec6310f198e08639f8d0e6a7102f7c8e20953915c9b282a96f60d42f53c7cd66908088a15f17e8b0aa8110c73c6cd6bd70da4d8392601c847cb71f5fdaaa5e8dea238010d45bb45bfeceda94ffcd6bcdc162d0b8a454ac31984c40c4c446eadcdafee373f58d887cbc818d477ce0f3a2ae5d6c1c0cd16b6cec7ea97b7c2b69e6d113c157ad9c9801007418ea34b11c51b7a9e800a025465e202d3230e289236f27778fef728dd1f42195f91aff86b3513ca4d94e39b58fb0c954bfca34b29bf5463052ce48d47b4a29592986f887afceea5c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hed6753cedb4e9b84720afead3bf964ebab1cff5ea04595c5867d769e02a8e1099bf55554f7a2e5028a8e49bc862d463a8614ab7bd397db023512d4e6f9c4475dab60bc49f70d0ba63e214e266807b7de579225d54bf54d1fc280b6984cf58415f21c951485a63dba5349c382a6426cc33ea7d30ca77a3c54743524a755c0e0bdc11c9b1b1c8bedbaf802ff80b7712f954b4cade674e65dc282d6726ba00b411671ae7854d0571fe643b14206829c2afc369aa867a41feeff3ee71fafe19b1c552fd08a79f8eb580eff43e63518cd9b1531b654ad5c9a1225d557785063407a6835f77bd04efa145cc25460125c3e773040c5489caa69066cb862d24c38e9df4cfc096c5cc987a0ba779b396c3b7445aecd0f1df26dfa33982881653fdd8001df6065bdc8a8f02b939ba5e8e73b144e68136f975af2b7d768ac8637b1e0fc14c6e04cc4782461d1850de4bc99ad6da8314d947da0c76edeaac19337ba0ba567123c15481098078d43a214f95150e2a023e8a96a8e385edfbbc4f9050eb21f61789bf832a9c30835196d6708176cd4c1d339def83116da622fa7a77dd651c93dedfed419defe3b16dd67e494403dc6da8ad3dbfc925da96a6c6e27e8a52fb0e2635cfa8cf5ea6a78476a3badbabc97a533eb55bc4356ee07a76e355323771f2c503a2202fb3e2ec21298a457bb155ad60c8447a698ccd9737c5a7c59b1beb5f57b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h98aaaa9ed54a37f887e9842e5e7b154115dbf7221b2d155d4fcd5e8cb5d9483ac8022027464f6cb512ea8c1ee2676efb53f392dd63532b26a749f1714b3ad375c731753b83b472ff85aebace1e1a0ca347f98e3a8d4b50b7b218a9bc8a4f92cac6b7fa8bc918891514b390ad7b3e120953c2ec3b06f5b6ea37860f7950c98c917df13f5afc53cbc74dfabe398734536dff9436787452a7292f94cdfdaafe4ce74bfe63683b241b56c93cec5d8e2150a06a012512dc006a8c751ab75386ee008918aaac02f81e8989116ebd5c5de1119adb0527a454155a4b873f98d259a348726889b5ce3fb49db78a364a520c0c7d06d4807aa438c74c690f1f349751471ea140267800286c704c9b0a54cbbe102f6efb045de0f3ee37ade4a26b222e9b56a20c0ccc42a8c2ec8d4f0d363f7d19e4ac9538ff629dfa56bad93a41a0be8754f4277f5b132fad22e139f64e3cb1c158c48c64171ab21d3f4cffa63524b068461bafee780c3bb53906fe93b9522064f41813b577ccff45c72022755c6f9bcff8e92f127303bb73be5208055ecc9200b03abd27633e210dccd49f251e2d14e7ea1293763d7952e9d3fd35080339ebbdee56ba2cf5cf7d2a24ed6b6683f557cfd07941230cb00088fd1425d1829895792dac2798c60424c0ad596598ece6bb7dc5216037cbef6fffe436ff620e72af0086adb2daa62a1023de8b93b8200e0b377dfd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1bef55a87c405bef54a9a0e6bc01041ac3edc62ec12344cbd2f681a38766a33129368873ca4e14c5d03fbb84b731b4ca26ed3ca003b83610d04eb02ad8230439904050c9a5378bcadcff6230f7eec9f903aa3ba906ab5165911b65ebb4a9dda33ba907246db364d7d69f809f034cf17b075f937e6473630c95fdb0648aa1bb173a63cb9ce08277528089f75b5fca91e73b4c71ac284070c6568137b2c44926f4bf2f6a342617e386577211dce2bc335f21aa016dad32382f0c7d66ad6a1daf4f706addb6b9875e7523f5ff41b5ec41167c0e53c08152e386a2c72e12edb3f171025c95c8e6405d9e186a3b6c4e487579569b49f8fe4dbf0d9d5c095c19d1c4ae8901a714bfeff3cd4227573be9065708c46e58440a757d513c598e7290b1bd963789b2b4421e8d61ff8446bcf4bc159c20ebc4775c4c8b0a78abbcbbcaa510ce8b08857fd1d80f7c1578a83f7e8d6b68d4d07d2465ac7f7a56862ac392d630a0a0d9e95bdb6392292a3777e5a019fbb86b8d1e2f2c1999ee12ff284896ffd190af6574b685acb6f146f3e222ca7aa348d6b5a97c1a5a038cf3905a7008d9386d5016e5560b00a08ea51efe5d2afe983c74d8675dfd1554f61e7530bc454213513920729521f34c916c0dc940bff768718af9327b791b6b047d6988a8869de4175c091753794c8d5cba66fc3351d65a27922a7d2d89511cefc68ea28a48d523c0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7c3f2d6e0b41633785ba486c39533b124b0810132bb5fe85023e8c084bbd622831bbccdb36de505068a04b13972e042ff82b845efb9230e83a894514314dc447d206e768d7c447fdd1037cce1afa0738ef6d77041ad9ce0fea7461151d34c5ff211fe3faf696959aecaadac63f87039bab81da95a166225249f62dc661b906cbb58e497be1a3855f4ab606b85877962dbb83583acdc6e54d23c2ae5fd83fa64e38721ce130d9845bf0276c9fc94b2541b530ef711677b22fac66a17446b979814b8506028b71ac49f9a46a16c910df81769344b110591d0a76efd6a5b1504837550e20fe9d3607aae6306917a6d619e51e6529691f665d3519436dda16fa5f2cfe6935052101b9cabcef39661e95a759ad259b579eddd7c614dbd7ba2ee1e2037ae4eb3360a68c521499a1d3a1ccfe4c4fac68a98b24b616fb17808cec73cfeb7415fb0166d751f45064eb159a1fa3d6d676767a5ceb1ddf1c138830ab05a2df07459b89219ff4402d9263b5f3df2fb9ae93500a77066c755891a3dafb69c343c07fdc7d6daf4bcd2ad731c4c047f479bee5b519e0805ab35ac61b0906bc5181c2bb52494c648dcfc5d6171086883e84fd311bbb45a277f233ee3a215c7ddbcd9af86516624934b051629d4b6e526a4190d92b86884983ddfa1573514bca72a79bf11d8fb2030d9dbf310051657632724250d6989012429a478f743bc3c6c4b0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hab674f79a16753d3bb000839aa82d353ba73f76f55b9a23be54ae181d7f30d9c15271cf1ea603bd3e5d70a37bc3f3bf2496151112da18554902fe058e64a82e59e8ccfd0f163c64aa35c1c42a3fc7fa1b96e4c4acb53bbd0a5a0221a0a4abbf3453db69a5f339b08d05c85a155c70d642e3c64c894ff3b439a862cf924bd01d51b30e5cc03657d01ecdb0d1e47b79e9c759f75b5d96eb0c39fbeab1aa9d3726601aad288a62090e29b89fb6e2d7c92c94409801ee480033a734de3a0250cceb7d409b20c713d36845693a36861b87d07aa85b0862982d67d93f91d44ff4492f369e5f482e3baadeb714d4040c95a47e1697e6a3dbe83656104a93b6736d9018bc260e82b0d7aa4b06f5b993deb9d8e26b925508a5fd1a725a889cec8fd4b0e646dc9b045023c90fffcc253773f971a9d0506f8437a046f816eafde44affb35bc0f953fb3e902a99f9267a8cb924af9e1ee31461910b65fa8dbd07103c607880fa6ef165ec8f4ec64c8e7f37dec1e4daf7e189ea37b2a08705a4d62e6b2081806fa7b92f18eae950297e91ec9f97b272d013ffab83acb6b14f8badd43eea406cb15be15b10c799a137588dc39af12e7b95fe8712b5a10ff176176c8e5e0a0592abdb756adcda5c9784f934cbb07d9f37f63fd346b0d5fa0a77986f54079b90880466330f0112b85e81696741fb891ce098c78b15c427b2148e27250744eccd829;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9f68e8a598ac6dab01d2886160ba6e50e45355a5873ffaf0837a4d375ce53e0d6d363718933411b27de020693d7440bc9e25a19f49b87c9f061140b6847dc99f91e3905ab815f4534ff54ba6d98fb937ecfb218bcd836fb6b12183f4a1b9df5a92954e195b6a9f2d0d7aabeac683d38a30cd56e8ecf6036b367c9f9f462e94896e25c7820e11407dbd6d9a5e5bbd33e9ba57bb8fe605f2a9190d215882e73aa11caec1dcd9a91fd35b73d6e3a24be07be48737284310f858e275a5547f08c1bb974402ea4945491ff4cee9a25e4e8eeb4ea6f1d31d15c7e59e35af29237abce2f283423b3bfcaa2844c6aa30ef780d8e06959bd3658cddfb22ed9dbb50520b8328b03c471c5e9bba7e76072e51624122e97c6ab74b8bb5c02055a64500e8b691687a22c2bdbe824e2f8edc017623c5cf2914dc35bc8b9a0bc8c6fb27ee19e8f4bbe5a121088ee5ae14e253cc35d3274f9e9e8a6acd15f8955da1242f69c9ddc35143f19989c78ffe47d6b82fe8f4316b3f21fe74dca95d86d22ffc00e36d6a194fcdd96898de276b2b28f15461f0dff4a45a1fb9a7f2bbf7130b0ab736397b1571f49c8be7b4271899fca17b97690102b497f63f69c14ff89ae02909e8fd7d3964d3a16f79f3c9e50d972971964da648a468299cd09e7891e36a2b7e6ec88caa33d5765fbf7293e211878948d3c9e30d72db379d724c25d3ffd20ef80d2e4552;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4580019303ff3de139a9ebc7fb25f25a77779ae7a1bdccd7b84409f6bc88e821999aa7c5d909589a92ebc11dc445cce1fa08455cc24b6d10296ede0bc67256383a679584d9c130c8b8b98faba5ab0255fb0b8bab0b5a7224e08b6b04af714b0d31e4a250848dfee799f377bd7b2cd005dbe3a1b92283443895bf41e15c55a6c69f7367942b74757d731a80fd22763d01c742ef45fba90649f153bc737d4a739c2baf32e0dc3265197dd447910b2768facf9b33c9c8328a66dd0166245e5191b8d6f3f60d39897ef7ac105726c1490c8d8a5aaa358ffd1dde4efabf9807887f24660b5807e3fa2440850fb3d4c5de3f983470559b692825a254a7f126c06d1bb2611b2e4c5b98396d067aa6047f3e2f1178dcc9374c5d95adf61923b7d7454da5552bc0801eaf216733e25bae552f3753d7f66ca40a0c87ea3ad74d415f12174473109daf508ce6058ecde47b9b8daa1e9cfd3ca705295b3b10e612539b36ab095558a531c1c886a79789cc190f4d8c262259622ae3d55531274bf6dca1bd53d392d85ecb4afdcab46f26c86d21162929c747ffa3478e7fc87b1804746b88e76d498b280665a3cfd7e803b44a4eb76c8581f1e17add3a2f044cc213e51c86a4dea6478afb69caba7227a23b11a68f284ff22c7781d3777daeaa4d65d18208ed009fd90f266ac5291aca6e68ecbbe9bfc278a8c60cfe23cd2b194ae22f6a9ff6c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb2673b7ab6015308f14fa092c6b76f224aa69b2b39a2344494ba827190257949d33f28010104e2aa27c5c09e62b62aa3363e8579256f45d245939c17da89dc1a74e96d85a8389d499e7f3944c9a68cfeb4f10095ba3cc2ff09e7b2db73e63e3e9b3fb892dc90dd67b962af24a8b5660593d03d3e698a3f30ef062b6589e042ee38432f66bf1b5d55b29d31d09f1fbfaa0ad1e5ac8401f3d565a0969228d5721fb9158aded7d77b341576ede56e02e5dc434ac120e16e1db295e1c4764c6d7f645cb224cf3c5ad29044f67c616cf33c6bb3089855a9abc1b11ad157e5bfef9e7713ff9d661296ee9c85056f66f7c0cdfdcd4cf1b80488cd256cd72e5ed296a591c6b3c1ca39646e60e35780c747d303a518f668ae364f46077027f2c0bac446561e7d6aa5029fc7fe1e1e89670bfd499ed72fa8b598c16945bbf5436c390833783dfe206acad7ecc58cb9ea096636f14749ba8029391edc76b5e63326c56f5aa923081880e5c161c7e5a14d6f250348a602bb20faec50df49f7617b63a92948785aa5eb88f33d4de939d0d7e2bace813357db287b78269f99ae570d03186fcffec972c6392dbe9b09359f01bc0781e1726506375aa607d7322ec6cd8320db0778a7d1bf3908fd03ea3e277fefce03da8ced02e64b6f4ce3b2486fa561c88fd150c9f5a0b8ec7df7d4f59a876147dda01850bea4548ac44ec74b0881d8de483560;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7750622eafe4f83d901bd34f5070de1407ef1027046ff55a3e808100df6de2fe2c6247a7d3ccf5a28bae072b71038221941139f31ec44863e28ffdf1278ca6e254010610712bdd5a642e88a051b360c2a4e34c47225257898151b75cdb0d9560ee7abb526c50c20accc1a3a7b2b0d6fab0812b2ebe2c6626d49578c04798bd17577cb555873e3dfea619837b9cc44767912ccfc0b4ad32cc14dae64e5389f3c7d5d9e3bec63b03c4f89492ae408bd8599e95474fd52e949cab2e8a6f7613b8c81d5f442f64fffb66080eb2959847200b8552dedb8ac4887174a1a309a8ef7798352d6a02152f450ab9d40c3b6c7a4f66ac70e7ed4f9958b3fd0b3657c2b5ee058568ec1181b4271d3700793e601efe39bbd9757dfc5faa45ef44f41b68de75b2b789362abc0a39a551318bdd4a44210d80222e75338d1c47cb328e667083be9eb90b724bc696129a4577b9878c05010347d2f67a1c151ca798dc1503aae3f1e232148d7ac0407dd6e2b1db28552d637fbcadf833538970655af7532493c306bc5d5b637f846b815b60f929aa4457c305cf6e8fc60bbc50eecabfe35e7424f5095c30446b5e7a87614d7fc919741cbbdba682a0a7ba38077165d278f83e65b045aa62510e084c301e49278590a33991207037a8cb45e44cd638d5dbb3be403de86c7ab1623460dd5f742dfc86084563700d806fe1f2656bda9443adb8fc74da20;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h40a703601e41a1ca93ae511a9de7b51bf439e0c0ef788fa248e2c4165e0f82405c1ee1fe00cf16a35960926f854cff8d079466280a28c8778dff5cb51b23f1771f60c1d4f281359447f654aacae4206863fff681b5c65a3d333e69855e1c8200d9e463f7edc57caf661fcf1e4015c719254cef4f6a012627cc3a82eae73f9c1acf78e3d751c7f7000ac09ab453db6305caf6e4883219aad03aab5432e9d50b59112fab04593a98c2516ca64f9918355b01e0f62f2d7a30b7dae4445fb69b44225b850db5e2c6dfffcebe3495d24510938eb55394c91080e7139ee8e571037fa1ff176e443ff55d82fbed2997e9775b4a77cf1aa5fbfba75648620c35902608aa134fbb9ffb22df8becce041a2156be03de397bff020adc041b2301bf76e4450544bbe4ae03fff8fb5dad848ab05fe0fcf867f6a2636e7b824345126a3e96aea41e1c3288dfd180c99f490577bf5d0845776aa9c8d31f2f9dd470722cde5be9192f43e1707cf7f26edd5ed72e046158e282842f8e1974b5ea5e8b7ab1b4d6e3833ff4a9fc07ad641a88654770d79c3ce970db76a9bf57742576bf13edf0a363949243f5b362b6fad9cda6aae79ba32a7eeed749eac79226a4dea67d7ed4de8d25707d374b428489adec349350efcd35e2a944c9ac193881f073df9688a975baf8de12777c64596ed5465097ac46ba583fae4a75b5a701d0f61c8618e809cf3821;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdbbac314c70ff109f6962edc8d79ae6d736087d84a7012c2ac2041fe1f975eee94b843d26845f5a9196a64ceaeac9f4f384e49f037a91750b9cf95f9d66dbec6522d24c198934d89756c8648c32b98a52d8c3b193d0506de6be6dee5a61ba54779d2049c3e14ea9db8a3291c744c3f2dd52b7e71f74eb87ca789c629bfada6824dfb4a9fea89f520f1b81a12db701b9e5fb665e2310dcb6cd7e9bfd81bec38c31915cb7f7a4e07655a9fcb6c15828581850a9d5dd9483565ed312a83e4482633dfde38692fbe3f282faeff0330cebf05cf30eaf34a8c34263b3de22397d0c0ad12b8f89b14fc30ac086a07deca87dfc90748463c64caed81f9d17d397775c54db60ead2bb4c1df784473dd9cf4849a52234e6d8164cf9b4b6fbb24a43207b0ab7f6fc6f9a5f01b3406494f339e60c8aabb0d4a86981b427a3af6c25d6c2805e71b532bfe70297e115042ed843f48886c6e99df43db56cd8d1aaf24cdc1cd202fbc649fdaa21f0600bbba85f0802212c358be56fd4be9d007b7f8f5b2611b3e04e07bf939113c5b698fc4da46c78af281c914e8c6ae2207b04b9839744be7a74c564b41a396f9fbd999b297fdbb8a9ebd9a9e032fe3ab4c6cc56f058217dcf35d1936a2fe8de0857399961733c8cfa06274bac77252deaa1191708282c979356e8cda26e94b38f1efa78b31306a8c967fb737b827df7b0aa4e1a60b1ac57b9a3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hebef50e0512d93b03fdb608e06e281abaa1f7e1966c87d8692a0a108f7ad0dbefcbe50f99fdbb6b6d6b272cd547ecc23a562b2253419c70778f7b6d39be86859c2a90bc16ab05e3da676a783a3cdc614b8471d857f3237a1c29fd81745b6339973ea1d27d72355feb11685cb455a5ff6258b178a89370293d856e47bee9619f0205470f91ff79441145bdc017c9c4821bdd3bdf8338d5a0e6dc57d08eb13cbbfc90d4fa35d239f913dd2cd89f4b57c253a44d337e63b48484d2dbf0c9fa2dd15382baf4e60fd2e71a100d5925d7d0d38f03166fac4846e735819b161c5a22e269d9e482eadce54f623b80f403a43c6e10c894aa766531a926db35a06ee276ea59decf97faf039da858e58a6ee62852d95a74f55f490504949b123bdcfee2c8d329b5aab10b1cf505fd77872dd7cec007460d0a7bb498f78989a784435dcf7349a114090e72b068f854724b680e69157a75da014061715762d536c151df2871be6b5cc228d2702c45aea5eb47ed9b214d54fe565ffb4bf157b67ee0c2ff8049f0a396b4b381e240c37459ccefeedf29fbc6151edbd70d289318050e43e7bbd4062fe73bcdb49bdaf6df4669f0ba3d0c2afa0d78611dbd97d8421cd01b27c7dc2363f196742039d1fb0939dd219ab835744473877957e3975f33d7867d11e4fb7222bbff02e77712ca4868cbeb9839c0e45536b8a782c58256a60afe4faff224ba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha249577d19fc6e8a1b6ea6364a9b36cef0bc2b7c2eb79d820d96157a97fedec4161e24afbdce9f01372d0a8b7738bcbfe03db1f3530e9b85ec56061abcc6c0d915db1c757a949376dc1dc9d7929604c4abfb1a050453e19d7c65d6a75176fe16c36fe24f173b9e5fa5d7cd2f76c7e3d2c85176e06d369dcc853dda6ba30ee55560a040fcf48701af3bb620ddad2bf1d87c7065da91949a08d89ae9151e59e013a75662b1fb45d7454496e06e3a42b196a81ad5cf29e7d611eaad199f2694c8551a4e190c463ef20581cb388f373cda4349a6a4572aed7cc514c9f925f502b769544dc5356739a2150ade27556a5cf8d7bc9682c607bbb7d4a00d488e7460df6c69f7ce8e1c116fab96aef0f47b8fc12bf193eb644c89eba69ce36b9e0d50396c52865657d44d5f0125fa2f64f2910c4f20b385b60577ee36063b67ebd3bd5a5dd7e9a4e9ce49d573fe6cadd76a8debbc721eae12207c77795ae01839c5166947ecdc68af28560111675dff369134bca90c9b327dcbf6ccf167cc5cc45e4ec77cc3ec9c4b7123fc50a29e00e76f35ee1d09c1acb0936b638179283a9de695314a6c1759e97443addc490a4227c02e54b4dd0e31482bc3e109dbac8b57603006b31a30dcf875ac5390afcd1bf46b7bf7913fde1eeafaee42cfc35fe408bce0f6501dc9e0b2083fe71ee5f13c0e9ac08f271f86788e29e14b32f5d5238bcc371363;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha6a199faa1c49319925a4fcd0cf7d461d30f8e7d6de0219a6f8b3dfd0ebc251401b5f82c7aae8866caa129798d2df8bf86a35618e073613c2dc3f406288674629c0609ba763adeb487622d3f847267cead65a9a56364d2f9bbeb6b5522349a9a4808d82b3c6566278eab2e1dd8b4136ca65739fcf7720a33dae53c3174bfb5587a8ecfb796d28dd57bb7475937b44c7938d2fde841b211ce7a254e23d91d8f8b3511a07ec4a6e71d5ceb68318a6170c91c508e415e73fb709bdd6c56a439dfbf001bd30cd14418b300e668bb57898d33e1151e12e2ed26e72d0d359fdaa92d985d72466e2d4658311d2b068c81afc0948f54f43e0f64a7613b91ccbe39cfc067843b38e81df5cc1b88a6f737b15a5ddb0d2fa3ec34421ffdf9771f3f8757d76fe69b0e7e3fb7d3bee5c4f58201f73ecc6eb62dfce6e7b216733e56c3f59c37913c2861d81e62e8da5a3d05322517e1ff0609f359d4519ba1df297acaf487c5bb35b83f2f40756b43781441fde1ab62db7f59e590d9888a326cb6e62dca512d3f00927b3b20a1ca62defd1b7330af103ed6cc96c2ff0fc53ad17a2f3b00555f1e5299005a48d4c88eb4bc8707e2b642a1d78415246613335fba4e65318bdb1422c4f223cafddb07bfee9464fff83afd41a06fe1ea7b57d3cc27323efd996ed258f84a362e0713a6629bb7e8dce0bff4a4b237d6799e40ce35cac2dc46bb6c7701;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h293d98487b6378d3ff542afc1084af2164da3770b0af7780460b48765c7dce47e0bb6682ea11bd95cc52b2ddf8c8dacaec7ad331218ceb981d3eaf5d5d851f9c510db565feb5333520c1e48e4f4ece880f885c781ac056275f6f363644748d881adeb3457527decdac36be63982cd56ee0db38618740c7b53315baf9fd56d29602feed911ae1fcaaa0c65eba321f0c993cbd82ce35a16302e58e322379cdc665e2ab38ce90f45863f331e5ab448faa0a38dfc29659508fa03177c676531e52c1b389ca820dd8c45ed8cf704e825f62ba299f7fdc517af1f467c08589548f8ea8c5eeabd562db8e66bc0bac62acb2de25f86e72d0fab0dc9cde22824d4f9ef5689f4e871dff069464d5b6bb6278bacde1a66c5df36b1d67d6ab3ef0645db9b73e85ec83fb07d074a4887a0b15b3e8a967b3450b7bbd20d86ef2fc36f4cf20cbd9dc92f2a92fbf6309b95bc67ac3ced65a12507d8973533ce3b148f08677ac325948270563f942e441205b1603e21a669e9a0ae7043e3838ea34640d464491fa6f88417c597d3d478d9506774eea771e3701dd1d5b7fe1f0fde227574582aead65b7a3eaa0f34f416126189674bb6455fd0cc37ef69bdc66c55b2a53b1e5ab2de6faeee8f2192492efa51c93decbb43bf86d0fe821cffd9e18bfc694faba5fb99f33cf9d1b1bb7ae51793848b93b4fafba25697ec01c891eeb1018e59973a4a5f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h73b272533c67b3df556a7134233f09e106ca9498b492748b104dc293418b5e7affa8e03ba6cc13cfa9240aafac50ddf127f08d1fe6be0f07a8829cc515b14f56dc7ed1bdd6b30b4a41efea2193fd9d97eb2ef8cc3e675abb7fae6590a297fda328b240044e97b6db5d69d2479571c5c0ebf558f1a851b83c279a50ec4a25ca3758ff3221647041365c5a064b88c0308f2abad2915d63fbce69711f0e32c02bd555499cbe79b4629e239e7be1d4cd0cee9ec90235a5e65a37206ac38c400c3cdb86c730c00381e1685ce4b988063a569f33e2a8f491971e2d76fc7cc4b39e456e8b27f1bb75562cb10932cdf4770498d79f6878c41e3623d5b7bbf74bac551066fbdb846422d77797c51f4d7b6af571138499560afd95e450e1b525a4b7c0bbf361530a9edb3d0b589aa4a6e8d28ddd54318bcd063a426454e64653e95b9b0e8d0f9ac959f20341dc54c744f0a510aac06ba0e7e462137f5decae8c105c62a8fe5d2230cc8ab2b69a9f6f91e2ccac48b046df36e04f4db0baa4cb506e5a92324806cfc409ca6c185d3bea8edd6165a43564bf440a800a581aac9ea67d34e83d1da20c3d9d6ae3754b78cc34d689651dd27c2741e2bf4678b49bba7daa49bccb6a69a31557e680939cedb3b00d36eb6005ef2e1567688f40caf4608757a05d1c2b91c9d466df28cb47ca11e404f7c97a83f4325eea391c88716ebfbc8ee5a78c0f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2bb563851b8ebbadbbcf27325350f4d4ebce19c3186402c55c4b8e289a68e70dc5afdea027c48ec21cbd0e41bcd4dac1dee5363c231ed8dcaa644abc7ffd7e9b20a9b087ed779698df1524fba6b6ecf6ac271c62a80b3f9d76960b8601e1d5cfb9b06493170cc88699afefad942194a01636592a79296f3808ff625e370f4513b720e8081cc2b3d30a09c1ccafb64e63386d51af931e4be56467e584c3985e6cc6a9eab3ac81ea05710af7f98be1813763f28ed5d21d6eaa27eaa13f439ca634b5635a7513121cb7dcf97d91e7e3df018796653700beed7ad9387eed241d7d9f7890b84d0b9896796a46000da7f4c78e41df194818932e8c26e53fd79d1d95163f9ac96bccc6625a292128a4ce82394ab901dc3c2a892ba71d549cdbed625b52e54dd7a87e33d1955a7e97b288398532da09299fbf243e3f32f9c404647ddf1dc04ade11a105504f3e3318d628a002ee1b2029944ae6a20d04f8ff76f6b29cd89d00400bfb8d013164ba95feb0c901bc28ae5e92914c2e13cec82068ab8c51662e5e97e9a17bd00b4504163081a0b9129fb2a306490b7c31dc5b115a25f5c52c6df5bd47bd33d5dafdb4ff3e09592a1fd7801192a5e928160cb05161f96172824adafe410b14ed35f332c3828b6d734c039659bd7475382ef20d496973a7bd93d2c6c479fe0cd1c3454c8a9b0dd940032b129e1935f02d87a67c6214c13cf0cd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hba848e1bc63959861ea89aaf5d21c2b4c84868484ae3cb4f3df3a383f63dc5237f662508bcea8bd3d53a49b861241f1cbcb0314786a3c44a4897ca9526ae1453d382f873c6e2c6dd4a962b95a8243f2d30e3f3d3d462f86b45f22d1d9bc4cd0596302a601d802ff2df4a53d0bce5ff7a66f331b1dc06e81e05b8f8b9166431005e86a786bbf3da68745d1ea8936155624184ebf552ccddd2a8f9aaf2f341ce1cee961e6af1f90b7172ff1624d478dced742515ff02720ffb219f0f092f1314791c9e2793723a517d9c462e0d4be947836cb03e03070692412c65f395caf6c1ac95eb41dedf09625cbc9dc355c743eec4abbced5bfa0fca6f4254877fa91168409c587530d16eb86e8348d6cea997e865c0b771abf771cf96c735bfad410e62171bb2bb9769c364175d855d1e74b8a287a457f03512e7db7f72fe8137c76b8452cd7af6fc5aee55b5835791b8784cc443172bca2faea4a8d8ce70af662fa664a8c5f82f95d6b156db68524691727786fc6fda22d66ed416cdd63b345838ee6e408c6326838b4acdf666ad88245421ee33a90e0039010425732cb29ec68b90170fc206c98841e948e612d500ef12a41fd7d8536f1911c3b6c5fbc0dab28eff012f212f26eb5b3b335edbc759d67ed57dd8d065b809ede44b5760ecff92500ac223d860d00141a70d1a14fe535c825133b6a2fc2a6db9344d1d147443c631fba859;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5a05151ed07abbcb09bae6d595b7b8fd2ca0412f8ff635a42f1782e9bf4e119251a17d73b2b315c9b7747b761c8c2907512644b34714145a7c0a9a27419459cbf8f5eed822df9c6f7394bd3b40cf401878505f7c38969bb368f617be94190367fee54bf9d0b8790af432a9dec0137052174ae75b3665cd57f02bb94d67825012a7018863e8e8b6677b461e8a361dcfca7af27f9554aca4fbfbc8832b95f3c78d0f2be005ac0f5349757eaf9610fdb4fe91d52b7b8aeeda137825f9a2614531146ca52f1c50a0ae2471fefd1a839b5b318adada36c992bcc46905add06e336d0a36d0f5de8f197280407027f586c500510f1e6c129051daac4e1f3f69b5a115d824f00a8ba6d1cd76ad9775adde0f8729265db0f2752bc2d238f6ccb41c475e2c17c86a1d57993e7a27bc2012bb5474bbf062660f05ba020e8ae0662b02aed1a3ffcb509ace71e79bc2248fce63db8d2cc13b54617185e3133238bbe38cf21a464f5ff6455ffd525cb3bcda92f3ed91e643a0a29338ea12915fc5091e2d774ca167e857664859d06e46649e5a4de074e06fdf29b1a2473398e74b52929b1133d90f3ccfb508acdaf55a221318100ed49e6c2bd0297e1c4f7d858384d72c74d79b5d21a3df098fdc9de8c92e823cd1b8dd86090996f85a04baec601eaef6ecefabf94e4ed2f24de3e503938deb60d656fccc726e9f1f1102b917ebda6bfc5a6414;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6aab0f1c22a4259c9945df0baf4f458f4b50b1098cff98a51d528e4c221d1adb520ea40535577886fed453ba7d09db495398461b518ee4779a2c5c6b18e607c9385bf271e1fb788d8316c6e7436885983ddac79c1b7ba168e7d53564eae8dec239423ce14487face0dcf01455f4453e40d1b6dab56d84f2c55d35af3a87cc0597fbf14afa1fb6c3772226f254a3efcc5371ca833d36e5ef769e60c3ab17a91d619297f8c51142ef90c7780d9388a55cdf87118e363da3eb91da5ab970ef6454214e3e2279025c2f0f58347ca37ab5aa37def4ea52aee696c61693dcf6b01410a213e49d8e39e4c07449ff3e62297b32fe049214aac9782e5bce5675eca3b2008d85f12c2ff231add9b5238ccb4bcd837300330f57086785806607e23dce70cb300c9f924c9d7e75b6cce40fa389d00969163c6c3517a17e2907cec95b301fdcd08e7f43c1adaf858f8bad44240f33e603d1ffdd1eadc30eba6d8b94c19fbebebdaec12880dac0bfa38ed8e20059ff548875c7d12cb806490815762b0f43a4344582406a5746130b06de796046ee3e436c8a7f1a6329b4070f01afd33b4a98cecb6abb64d82279ae3c9233bc532d48af633ef91dbc7bf4829b2164bad5359daf0a8bcbcef5660cb80b22a8f4a52fcc0cde9194277c2c49f050230837e2883121b3e99b0aebe678d2ae25187208f0a970929184b77e58dcf6173f14fed06029f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4cd4857f35665d913a67b1fb979db1fa023c7bcc3875955e62931519d1d724fd0c1aa85ce8709b45f2326c0ef7e3beb41a4fbb7efd2c00373d2035195d6077f44377f584f0bd0a8fc2eb1a6561dbdf24598eb28711494655e88649de6a5c4a16a524642f72bd1d2b1582a1b0e137c44119804f8ea1cacfb7e33e89dc9e3b4e121520835543bf2c43c40e3123bce63995ccc723f294c24d9399f1d56b28b0cc9729cb85e7431d95b860cbecbbf92a24d20bfa3b4067f4b6e6f2d1432f994efb6116f5562f502dd2d4762c1270ba2eb398b3fd8b60948968d6a9565961d2a02ce01fdcc96df2906a95cb167243e72248877f7340972b748e8a6f6ec463e4564de37432e62fafbb90aeb7e314f9b14e4b5eb8fee8fcdf2162126e4000ae2f01a85b673f7847f839dc0436afac4d276564d40185f36379477cdad7968dfac377764e2bf29f13890f6c5cea35cfd22931570316ff3b78b4ff9688ce83422c7029315d9e81893b1409f1645241dba430045502392b3c5adf1e6b175435d4a74b2affb28bdadd5223934d8262f47d9ec8da6495ea4dda96b36b8b346931a1047f94eea4a758e1600060c433c494eb3c9dc95d87fd100e6941e51af68abef72788b0f5584776ec3c7163a59148700cfe8c930b0943244f0b64983aeb5ce41224f549c05a2f93efd5fa535ed1b3c9069f702e0cdf22596fe083df7a01e5c0995ec8aa46f5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hae2cb49e59176e5c90adaa0189a67fcd62992e6d45a3f2a801b10b73633837608deb9b601069bac0b02200f4ba291b7ecd824e3aea8a0a0edd8d44929ac655dda6cfaaf986c121e9c63d532b7ee8d154eadfcd6adaef959bd4adde7605af969194a9884014ab4187f5403e6d0a969dee275db52fae58c07642c18c6dabc22ed7741ed902432a12e1685907fde2aaf9447029fd7e3c2f12052580862edf3daf62be3ddae79a79dfc1bd2ed9a40ba27ce6813036864a43ce8f7bcd656a39d867399ae75ebc24ea94cfde44f112e07480e87911c37adb4eb10e00ceac80af82fef05cbfc817462b8e777f9f48713192aef76d975a55b9a48378a6a45f3d9d8f7d222928a68893f82d15c02c8c334c0ee113c58e0689f910f95911c12440ff27ab1a8196b3480c98e93a49606b4f15a4165c59b566576d9ab5ccb5ca47671ea8752222921dcf6775cda551e771b9cfc5e32814c89554b02398c277cd55f203860968ec76c2dd8393a70c93ad3d5df4092e760a138fde8393b33568a8c85c7d6a622d12e5e31a27a38a79145086ee3e6f21fb71494621d8bb86b85f780701e602a973b4403fee8f52694051a7b130e7bd23dbea3aa18b11a43c35a6124caa4ce347a4b0f7e40836e45701d792f1fec4d4c0ee6af1807bbadab7ac9e2b8af86bf6377cf7071b0a4feaf992d4e173678c19dafe32762d5f3f74565b8f5fa2053983f600;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8f8b002257619f2790d8fac2c7fb5ee5611d3e22352bbb092e7b95c4dc879f0d19751e52ec4d7e462f57d0764dc34ce2348cd6897d1940cb095f4b00818403e64eaf3f92c93af8e70d66dc2ca9c43fb579839cbd774bf9976939c5a1680bddc3608bf9be8978af94b8a66cfc4685ebbb2b93113ed82d82f064d43d63addcabace9f32108184c5429d18968d85c0fb1c6e0fcdb842890743e88361495f6beab5a94c82415a1de9fc3fbaf79bb20815e1c660e23dfde20693f3dc7c65c3bf468324b81736ff8a609bd4867ed8b82524e7c322f212df301c5cd4281f9ae893cc6d9ed2280ce3d6f0c9c9865f1c5d2e2b7716d4c5c9594a64ff7a6627c33119844ae5814c2f44e0bac0748ea7ca58a129bde9de9a83c2fa81346966b8d24d5f0355c34cdcc765bdd74159f2829df78cbb5ac11f11da9b0a073a14c56af6761f671b335644e2a0ca86ce4cfd6e36ba7f943038301ce25b8e5b25b4a69de7a1e01eb11a5f20d919a6f438a57681cef14773cf38071948f38236c2c550007531cce6de162bd9f492e2db66a72cf29b7278c4aed4cb5f913e348f2eac02e5c663fc4ff4b34bbd0ae6468701419da5b326bd8656c3a6c7f6db1fb0a852a057d7022b3abba69fa9f004229ffa6f1f4229eff59b9fee2c332b3cb813abce3c2f29c4e7a64c812dd673088f06b2ff0d95ffb7e7d77aa24d9b2af9bafd93aa4f12a2d92363e10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hadeb9d039b6f68bb13ab93cfce0d9dd77d723f7d9743a176964513aeded967c44d1e1d0e559521eb05c6da7c2860609141adad80f22afca9b52725fee173108bc8987d4deb90d7c1b3b83bc51ef43c7780fb614f2827305ba267f57d846bd0b8c20240de5b23e95ac51eb8e64de0e50bc28a7b597146daeb1639cde5649bafbe3749dd23101d6bb30c6dc94fa468544b2c731e1de16687bdbb63237b62c2a0afc5c1ee242c83f58dad82fe81a62553db4322914234aeb53d0e589a67ebd90542c2b7eeebdfce73fa5eb1ab257da8f4ea9a8d284511539168434a307b6eafd88935e94b952df49c8e5f3ea3f52975a629ff789f3b7c736660c40783b1097ba04c8c19f62b27bfc1f08490964b89b67b8eb14586544688c533b54d77d218cc523bec39597214281a88d910cd4af78ae44c02ca060ee596d77858ed07e1a91a0a670d2da7ba8912eaf58af234b04fc128def050b1aa9e3fb950747cc5f490667781b05c22d866e6ecc8dfadf218e29cba764383d95a58bddb9dff29838865431768df3d710eaed0be74668fa3270a7710f9623c02b37254dfdb32897afb8738f8b97b1d2c0418f132b7beff529ba306111c7d4dc9f78d56858a4957a2232f13c8bcba1e85b8957cd5820d5a03872a0da5b121e675336f4204d3e1df5d6091f84d15989167b04fa42c29f833e6cb79ff2bdcf6da9cbb2910867068faa2f818ab0573;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h50b6a3b03eb4e59b62804eea7fd9779efb7e87eabdf824b180f31336cc2d75285264ad3aa825c7f6f66c4dc5e8177d53fd9b47e05946a2fc38a9de6b058e9d256af8e0b910fe56dae1e7971ccb54046471fd271aa604b0c4177370e16c5bfc6953cf4b07485321b37ddac140c9e280e4a1294b21c3dc3bf1fe10b4726780126446c553c31c4ca370fbffe56be141279fd89baaca5e3b224ad8678b66744df92c29298e108ed55261085239e00b9bd168aee62bc8de239bab01592103b54b76fc1044f7d3f48e0f8910101e5b9106dc92ab13b53b4e82a7760511741c60e435ac3f5d2b8b286c7a6b299ee86556bca7c2037509ab2f5183c5ad55bc5e6efe3838f34b58070b927daaad41f5c9ad5c08194d9719cd35818646b409b38fc2e210523d8ea64c65fcecefa4a33a1a4decacb43ec151de6e54a606f9cd442400de66afc341f6d5342531e6e300472ffe4ce6cdd79ef86b433e5c729a04033b8b76dc2d1728216ddd77d1d913ffd2e3e782dbaf5c2709a48c93c6cb291ee33cd1004f91f0ba01bfb35428a2831f4e74d8ef38541b4d5fb751593a8611e55963acc331ef4afdead1dc201d36badf2a058d09d45474667e1179fa2aa6fc72c93cd3698e68030b56257ccccc196a10009e02e2a96837ae4fd2db02ef4cea841d9754a404f500ef80d6e863525f2301c0e433c965120b07cc5057568854c50aaac47c382a9d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd3fa5431b5fdf43525dd745c26310003ca626052784bdb63942960710b67e441992bb55436b14ad1492796fc61de08d7e3781411583c8308abc791ca53a5b72ef55c7d5ee6fb54c7985fd68ae997d07e6ffd63f9907a49b996a6d80e686ad6b4eb4e1ca89c458d4b2f3dae05e66e01b426d72794248275fe851ea535e57f7625a472c82ab01cacce4d1035e0314db99d8e8098b740091647b7f05c4753ee055df10d350a3cb857ae6f187c057dee7d1950b466375a443501ac5890469f60f47bc8ba9c6d3bda4d53f1a35d4428b0950588e5b264a7eed5c4222cc8a7713cfcf67de2697795df0760cb185aa83ad3845b07f52564916e532169648bcd05ae044328602d271565cc614eccb11885beef9877401857e1f4820c0b34f5d0973877e4b6670b98e68fda1daf720521c38f1e8c076434ac08f1a9a5af983edef9f0b8bafc8920bdace3d94025088cba2830180f462fc810e8c83ec447c894185529c4b76a639948c38871ac9fbaef1b7c654179a0dc5747122cd73bad0f200ccb8806e65f211ff1eaafb814f860222e4001103e7815ca2abfca5050330bab8a785dde43d11b6a252a0b772aed34b94ff680bb760db116270b38d9b7664944f2af854bd0f8aa33f43ecfd6ee8f3d4908183972feb2438d2bc365ff3f4f9392b9bc6e5e92cc21a91b52733a59df50e799c77c5d500a35b60ce58807371b75d165458d20ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h98f33f794d8cb919c03f80a577f027e9db2b0e4f88760bb53f2097649e7d053d8a6d621190fd1a1e832dae3d3662622f4a4484572285ba9caafbaac96d0fb5f4f305ea092714599d0cf0b22b1e22a9b007585aa07d92113a3091f4ed4cf767bc6a1cdc3a35d4b8273b7f868947c0180cae125955728508cb779dba7e59d618342e220b4d2ddf43580f3a593d5d08d81088a8bb89e377fc0dd7618c3553c8983eb6aadccb5bb02a75cf27ff91cd3a43618f13f478173a2ea4e771b7b4750bc6028a69963a7ccba85658b35043039a373d0704b09305e8d6d81545e88ecd6fcffa12445ee16498234dc6cfe35c4860cf82ded1857b961f0d73aaa0df78c437f364ca4d80ea74c34774df9b772460af2ffeae2b3d77d1b4624596d11ff81c6a0c17b3757f107ac66cb2acdbf7a7512f3486ccd6ddf8eaf728fc2672b5c18f934fd7dca12210f136965bad922836d44b44f1a4e6f51744e2d1d4fa8e8885fbd289340c79d637dda6fe7f00d5abd126a54338dbfaec841b856838a0a7813f970e6dbd7d013f3697c2820cc36ed0729e247040e7f67fe169be006b02aa9cb8cde7a8290ee03f49f4d9c7dc656fc922a92310db6995c549570f4d37aabdbace28561372e869765bc94ae2822d379113cc3760cf6ca9043421ef068d758f7fbe5313adf42854b719b997a3ebb6eba68d4f1089dae2fbb12bd3f42ec9676ea47e62ae5f5e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h677dd6cdb870b5074e0fd905b1d7dc74402ba26a9196a0f1234ece0140ef1adcd49f25b347840e7b0172d8e14859bc6e7beb31ca04f9c3dd9a55cd6548ebfad805d963ee03e83f73d8ad3d973e9ca154cf24da74a5cfaf16f926665e07f5d627a261b1cf12768481c5237d0f865a7729bed46c28fb23dd60d1029552d47b0168e3648274600bbb13b1152986c0a2df5c34e957f50fbf25becaf9f30d0a29d272a95c619679cf29b2a03e450451c65acd6a5eb7b6420623039ca9e09b727096231054ea60266fbcc2331c56de6c076a8ff06cd15ea1e370c7807ee811dafdd60932c0d581a593ef050954740db6cafb70757ca566943d25607a9514e6f1240a83d8cee4f000850e4a378dacc5f650bd7ea2964de3d96af741a6356745eeb5153ee004ac85160a1fdf111e00977bc43f0b3dad8a3c6ecf91ab61d26a7674cd8e55bf57948d04bdb6e8b0298ab4bd5924256544e8b479acccf2bb6c5a8063fc7e4f0164a16ab53fe33008a91e507f9d5277ddcb57a6847f8b4cd951e3d7c67de7e6a458dbb634b59f63c7bb4980bce971854a36c7066bf9edbe5dd0573d5fea9e1c93dd2286a495270fbd17947577a6d7ca12a04f099332006f8d2986d9321fa3aa61df9f0603a772aecdb4961b8ea043c6b8fb0b1a0f0d735c80e67e968a6dc29174ef0913d57c2fa1087c895add78c693c465a5cc1cb9c44a4805a9669775f01f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h465cdd391182b14a7b668995fc8ac16f005ec2f1979e5f098986f1ade4e7e519669e43c19d1001e8211e5f613011e0840d955327b837ee523e8de2b1c8ceacd89f22fbd6f8e540819f953e7bc304df3b15f495433974aaf6093ba50af9fbe891e3fe67c7c9667e99cda8c3a6eeaeb226a8a487c366643d7af23eadb10f8eaee827b1680c6cc9abaf5bac9c09e5cbaa051e167eea3199c56689f226b61f012b78fd891db3385258fc62aac6e9757af588a434d283190182f9bff8a90254c0acc8c6b0df8e6de5bc7269299991fa264581a60d386a37c0b7ce8845e4e94bd2d33de2825c4ce84e90344fd3941354eb80cfb4984b388c6220254319f1092c0d7eeb62b99cda76d6dce81a31ba6fe121fafb6225e1ecf759948c410532e99f073bfb30c8744d521f36a1f7207f5d9ae288c83ff39f51a08c1982b54496d66442d290214698f659fd9362feb153cc69d45e4a6e209896c65af5a52fef0e31433275df3e298c438ea69b5bbc7a6fe2cdbea8428956ae1cf8a485e568300129aa6de1994176f43e4db3336c41a0f6a4cc7def39247b76227c32cb1d63e9f0f528ef1b7dee0f74f773542d7de84c7c7e005ddc365c61cf93baab774891d935c419ec49611853c8689fdaf509d85a4cd8d127b3c9fd87a9ba95a3bdc5d931dd476f18940b728f7f8169837dbeb46c93cc5308ad5db85b1b85030c4ce8822bf4cb76e9ffa6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h99f47d91300df91d39926c9757f6140d9762ecb18f54c05d7834f72b26ca8b8dd5f86763409e40e02c9c34943aa2fb624c85a9f7d9ef8e0f2f2f95bfdd0f333f8aa5008585957dbaf8e9caa6d0ba68d85962837fa25d88993e999990cf37d1fd5c63d417586900a20f0b02d79eca4b805de8f76e897cf86d5c36774fa68522a891ab9bf205b126cbfa4b9d9aac6c46d9d275005e2c11f2dd3f9101a93ae36b79e0dfc7591fb4f5810c715e7cc43512e924f75099eba283c63dc619009476933da3687ae8ced9561160cf48048e1f722a524829d15d013c799c69b68020dce781b79d8b22e9dd706195d85e579401ccd90533f27279371ae5001e914a7e048b473619023fe7b2659537c8082c8fbbd4a73aea9e1d215af745b451bdd30dd203de9a91c6b2c36f3928079a42b8051af47a0b18c259a32c068cac3100f1c849aaccf1c3b5abd92bdf5b35aca8d44219b27a87c9a2802e2f7f63ce5347ec4dae963b8b760cbd9db5a7618c1806b7ab32df067ebf08d08a401822bf287dac15302203bac3e2d17d97e8193e84c38293e3ce7f14d9de0afdacdc5593119d819425e2f2319dda409172378268cf678c72c10dd76d9d2ea2abc1697fbda59c1e1b1107314a25197020e2b2d2aeff6ad17d1af12daba9879ae19a1b5507d405c1d5b16f872f7f0483f37a193c071400ec0086f92b2873c44c2a20ea0d80b6a686992e0734;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h461fcebdaf812de2266e06d6953c22283eb1d5e410b339e9593a619f172bcfba8f5b28e054c6dbfbc95017cebb3bf8048ebd53371f8eff07239e10383c93ff6507ab8cc2b54cc878ff6d9c7e86b80db4cb0a17b1413e653d9ca39ba3aaa414b21823391946b5689284d7f6d5ffd22bd64bd94858b1247dd0d2ef335ce978ff0807b2adca272bee559a538572e9a68ab69950c66748d4f745b311b465e7bec7f73a97cead3ce3561a65919ad5da71ea5ad53702393932b4b28fa0f6b783ef1bddb9c2d34f361d2e8cf3633ae462517ce7f0eae7a092d7c61f506176c0c90f69c0632808386feac8df4fcc6131e92c7f10bf96688dcc6b6fcd0239d83ec3025694c05b196d49be1599b8704c4c48a35874ed066874eb8c5641c194d85c56734f4a2257eb515e0c80220096c3e9ded36e3c28fd198e3c5417e4c74986a8a0509911d16215b75c277ec8d1ec4a4ab4bcfffd9ac438783da6603d7930957de4ffc06ea153ca00f5ca6ac68536ddd43fc298cd9efdcfc39d1e3a6acfeeec50fecc1c7475f225e09dc9ab0fbd448db1322c8f599597b1e831ad88f1b8cf35915a358365f54c0759dadb5da2d2be9a2461c733b83b04d2e350e908280ea2671ee43c7b1a88740c58b529f6a1aacbf048e528ed4d58d08221e222856c605b74867bc18618161f69535a3209c3ad04c1b056b4a63c6809638f8dcb9c23d2925e82e1cad748;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hae9d65e82413b3c78a4da8851d55a57427e654993878724d4915455f0d70f1c3adb099a642b8729efced44ce714e86eee08ae85388d521c024ae7025a390f11e6d3d925823f5a0da6ede24d2e361929aaba3345d1083f1135aede0f17f1b129c5481303ebc52d2e335e72c0741efabdd4247b718d70b3ce86be6a9e976d2a947d35ba3dbec988f950a6cbbca6b03d30f56fb91765799ab7583331c35cc3b27067a2ba7022c583fd81ca2623460e02d323bd334223294b52f0d6e64bb0823e30d9cdfe7c7c2aa14f977ba6f6dd7a77f363bafabfa92a484dac450ce9d5f9ddcafe9ed5132411ba528240a20478c89b2ff807dc8c80f88d9fcc86dbc3a902288e4e90e42056fae2c41113575c80bf1f823bcf8a899cd78c8a6bc5ee00e6e5557be126463d8f067c9b46d1be81661781165378c6bb19b20d55458017e1f312bf7e23966248418a814ee8906456325e458e45fd49deb96d8a391dfa50765625babbd4b104b2ae11caeff953049678ef150affd1257f172c4da2818b0465cd2dfa39d9a1f5ef4ab1f6421ef5cd8c1118cc45491b3c77c8d6d6315a627bdf9c252774c55ba67e43735414c116ff568ead9b4f05a23caaac9f39a812c5d026da446c03398b3d24374c09c59e19739b40c88acb6fb2c2ef13d1fde3e2ef5c41c2527b72902fb179de85df83511980332ee95b7db4f4829ee6c09450ee23730316f51a761;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h12471e259d372c5f7b66eda9d17a4687844383c899b078cc5bd930a263576412938c5a9a8adbacf3857d0ae083a641a64f165682e9bf241202c3f6c56e35bd4b4a80480d956916d53507de23a65b7e5174ae24c3eb87eda8a8fe9c3e2dd007951e082712fba3aade376c0eb3c638473bf9102bc1d0d8f00a083d436734ef6090713f890388056d1edbd56d90bdbab1984572da315c7b69269e4147138fde1e6916aa69512fc077db17eac4e139766fa982c7b47066fb02a7948a2a717d351117651bffdfe7471837055b49f98cbc8fa2f5c30f8c8c7ff4a2efaebc6e5575aefb317f381eddc2733a7e2803010a5f2a663fb031fa62ae30ffc83731f8e153e116ea0382a1f5da8b2aeb50a89af9811d96b04d80e4a556d7c2c3281c61a487bd769ea7ceba5ca3e905ae6700fe3ea8721eb9b0c0b0a20ce0ddc288cadf53524e9213edc7cc7b55ca6951261c70bac2c4ae99fc666c941808a8e2c004e35f19c0945cdc69d279261bcbb5c0e867161ca41548540ce04c93cba01a393236bfecb418394aefd3c922c5ba7e60d331e9bfbccebe612dd875467b7ff931c99f0808e680a0c05e49f9781e90cf2317e5f53d9eab56ee93e4b0333d8d8934c36e4764b22e5faac0d5880080a75489898812212d12f8120d86907ce7078e4afa9bd4920f491222792224ebe695aae72c2d641f4a5c600c5a29d9705372436e0f4df72f699b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7f59220cee58769564672e17327e1b838c94094c2eabe3ddcafcf47ab84922a2a54442897d58e343366823d5d84bfdc05501949f695c6b0e82ef9df5930d3bf951a7618f0daed9d9a51b6bc682efa8365a97779a08b6d65192fb54ebc84a06a7d55c2b62b0a5af11b71b5a0096468c8f2be0ef6a91fbf7bfd03db4205c9f266afc1e23d2c132b24a0a7865e258fa53728957a8e618dd0428f00ee5e9f334afb74a381cd7ed44098a09b5be465f5930f9cc6a8990ffaa6411aaf5ce0f7b786101ad7c6b7185cf772bd730077e2a0733d1c8b0c0bb4764bbde357c74e832329537229b7fe87b21658c57bed59a1766339f86e2af9a341a756c6df99cc5f780896ac40618a3bfa2aa562ec54ef4fdb6a0405a04ffd67e7b876b36ab074f1b927dac1b9dc0c921c9bfcf2beb6df380191817236421a65ef72ff61ffef3c7c031c93fd115d08ac41194353600ff14eea3b614bf30dcd01473ef3dee64c5bb64fb98c6a006ba0d7d2528451ab292ba1d1581a5ea4fe6fb4f35f6171d1aee847d12e1324e7523a9b9b0275fad76b375d8b768901f898d1d361e45dc5bbe085acdaa7009b0abc7b667b90867dc9ce4dbcc9cc5ae71555187ff0d1d1b0616786b7e312ed33106151e5aefc2cc612e28d950d384b5b58a63a4858fbf45142f03c6b71d269a8b2a9289ae8d4aa96ae198e3602bf4f06fb20393926c69671a6d2835795d248f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h36bf29d398a81e238950c241dd7f94a163d3bcbcf041710a5e70046787017603537da350dd131e0d5ccd425eca04b3c4260fcbebea6dbe99f2d93a84c9a6126d4b6598b727aa1c139206d22b12bf8004c21c0df9239177cac9ae3bd3f3b6310d01eb96a89c034ccb05e8f65d76a64058a202e76ebf553854aad25f8837f404ba59924b9dd93770cd54b36aa51ead23ff60f2585c17cabc2026cb4edb1e849964baa3892910d8bc2d4f807b4c5412a93a200a4595b18769af3e183f15a8e1882e2d2988ccaf563c0febe0e9effec1b7747c74398835e82db94ea51f958d4ef4e6bf3775fd7f38450c92b9c16ac86e315946d2469cb3a38e57e76804e9add8012cea4687b56c000ce9a9238e49a0f4315ccccc1a9ea239ad2b74de134b6b48f0657ea143f015d27adf03a1e060427605fa0d61cdc0f86458d0aebefe64b8a92d9c02abc13074c6bf9a40790dbbf6065f6543d7cd3c111e81ffc7a3d7730097ae58e044a43075ac024f1338b76ab268c26de7597996d848b6106eeb7215d1ac8363450c662dd88041b6c4d3789c706b106c10a475752b64c376c345982349819fdcd0f68df83cf42e8b8dc03a5908ef9a4cf409f9ebf2f52e69c413475663b0ae40700225f5ae4d362ecde9a85cfb7babaa12e3d5ce7d0cadbc5e197bc7237b15b928687c50e48272b4c09569c3e204fd89191d97c68e3611dfcf893aaeafd8b85;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfb1b471d1ff05e76cd3b9de32da440d45ee649a6c3d15234fd052b0596b6029d7da9aa7d15ab9a2dd8c22d94d5a4179394ca1b114270a944a5bce27875a8aa41bbf0dc0f21f9cc50f06784136f2d05408e5c2d55faa07c8b1980f2422351f719f084e7f5923670a2f82c764fa34b52c90b9488c0b7b7330a841d8775c87f4e5b4e726fb257e953db8c1248140497738dbf98841037b032870fd51cb3f726ab6827636f455330309cc7b949ecd88ead3b315e757dcd3a457ec8bcb73cacc8ca08b3818e95c9ec401ede97f5a602dbbf88c0c13f5c5cdbe3022504abfcf46ef0f5d57698168d2d26d657078d875213bcb5383873039d53053aee75686569c8cf491433b3b143b6e942059a6faf1bbbba9ccd427614cdafed329d90be56bd4e6f4ede76788c1bea299129446d1963563586b9d13f3326a163f53a1aea8016c69c628410f84a5c5bf9cd2b7f61c27587bef4a879d2464ae5c9f6c42db421bf60b86d6d98792812438c1af3ebf5a562dfc8ffb7536e84bbba09d043625cea4dda0b73a8bdec95d18092684075c9bd4efa988897f726f2e83b66b0de67769567497386ecc795c8b3fca529668a447a9fda1b0634ce3cced70264605928de7794b173b34ef8361fcb0aa52141fdac65ef7c01276c56c72fab9b9f7db6a91b1ef3823d7bc443b4f6e040f87d403abb17d8b486c4aa6b6dc92664333b29c845ccb2a42f5b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'haf35182315a9971c09b6c4a79f4fde0ccef886f8c8941502370e0cd63861950fcf53c1a05942013a71aa4833db7bd9081a6c6932e1f609953d814813efdda62e61c47fd4bfb45a3d1cea21ff6daf5680edb0154e4b0fde2e3ff345dc8e1439533ca6398b45227085ecb57625b1ce5ef5a3b88fe9246c387e2bf48308b139e7f1492428be4517f0d90d15a601c6846a1baa29edeb9abc9f4b93cdfd652570f420cb56d8428c040f225abd934c47c5172e1dc6cc4d90556c845543df5ea0ccdeb41dfd72ff9ed19e087e5d8c153b455ef33c883553a2280ab60fb7f07c0122b6091ee37e1410560059cd7b624b948d5ee158bf6e9e0a493de8e89814dbeec5d74087fc6ec88d35c89a86b9fe485685150106f9a99bba23eeded1c7abfe4f26e2f03b4994ad4b5cf057a31b22908792c3666b91d5b756175df3a4ddddcf72c8fcf2248e6dcc4cd203ec4c710b97e10b95a824409f852dd1d1b32df62bcfa58023e46d8d1facf2bd586eac5dda33d293271ef0ef3ca578ff77ad24952446e928c3eaacc1e0bdc71c5732c208a63c7cb4328198a54d9c529eb5afc15f90dc4a9c189ee34a37ff751fa06fbe847fea46403d8ffbe8956bb90bcb8c40d74e49246bba54fa21cc3fe4e1538b92a114123f95c9b13b290aa0f00d812c038bed37cb73a3b31100d7c9e6387915084a46f87a59da660251e5c24e2fc6625368f10b6c04078c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfad49de5a914f8d1a7fa153ae669ea78640797d190ff4d02ae2f6129d802d4d51e491ce08f98332223f4d13175d7dbd756883c20d58d0b6ee84a7541d7bf11cf5b21e27b83be322a15107dcfaf0d251e5d749c925f18e7477e2a3054cfd3d81cd08d202b16d3e468eafc2db824c8e90bb3889c6e352badda0c96ec4b25e886de64ad7b3fe3f3c33c350c8b0f061bdee07ae50e26cdd30b6198d9a2f23a0602d3728a62fd74c7b3cd553e46b21d9358fd89faa65226fbcd226e69b9b52619487deae8971a723d922cb0c05a24395cc8c9b79adb2be3e9e7901a281a3a89f7aceb843bbd3f4ee10cd2b49d076b6409b68b0ea0a03f4629d38968fd0df5453f69716613c1dd00df7852371dd11896b8c7e127e1da913a18f840b32a58e384211e61245884a4eb7a8c7b6cae8c807c5f5164744faa6ae4d8260c2acf0225df95f3b3c0749ec686360e5cb0a0757a1dc710d535d534603147f09bca1eddaf3451f6ce6c02d525570646d6ecaf1d242a4ab68ecdbcf3a629827d08d1065c5b212ea8017ea0e57bf37f0612bcd1f8e95ba384fbdbe155000d6125436f858894f1bd9b85ac8961cfbaf8087f08ab2146537f0361b5ba5c6cbaa078e3d1a8904b5def6fed5ba7912c0f2b51f6298fa3c215aadbffe0729d16c452f75756d7270ad8c2824af77a3e9b5217b402f60ca5badc5a3f45ce947ab0a5bd1aa1e8000b6ea5ea773a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcc1d13ebdff635192e5ffdf6b7d242b124a834d0047e292c37cc542f0560fd1404bcd67666aa6c895bbbf9e1c756048ddf85d7cd911fe7a2e4a6e79ac380531015d5ece0ac5322e8c1ad75f91c4e5e460c6699961e2dfb160b051a827867f1e4ff9368450bd25d115151685547e3aca5b2b9e23302a20aac2e2ac6d29377a1d2e2863d29951b0e60b6049837a8a3693e9b2da0f97051308fb0e1692ed2e221cc6857a9d8c2fd1e2825077bdd9f2e406bdab58ee3f553008a92b52a26a0c95dfa4b767f3fbdcba9f9d87eda413d6dfd9fe08d20bb58743cc1aa2c769689e9a50764ccc31f550f61e3f9264154b37eba5b039f1105c60c8823d212f987459787daf8e81fed066564329a9f95189ebe4677e8e16bf5cd743360d7a58e896b771a1778f8c0db35279211a4464668ab994974bb70c19862677f5558347daa618cf9f074edd967f3ddbef2a813e622059b408fe411cfdc0b51ac9ef20e8178cf533d86c393d21d10d6612cf54aa3caeabfbe3a62a8045ebb2f8fbf099a6d43fbf1083a3e4afe74c5fcaffc784f94245bcc88dc77731ae3c3ef79e50f0f2cf12c4d32161aff69dc14c54cd818433de7e1be6d46c2555baec543b150a8ee627025a8fe5f27f562e3d897b49e27e54332353d44aaa979a5ce5d7d7153830f5d95eff0e30c2c22feb04ab5d16f93cb31090384341e33ceade624ee6a2f3f29ed10c080f008;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h12d8723eb30c0d4d8523ec3c9d72a4d5d87178d5d30d9d099014ae581036434f3926e4d5604c2370d9a92e7185452eaaa34fbab7600e998ab458fdbce6445dee9922a7e121e55045f2b3bdb7e630c46241be117fb2d0297c24d53e85fa84c40e63ecc20cc536db74353d9082163962a4124edf66e6465a6271174d1727e3af680230c94dc8b2936fc7de2126f0eb6134586d34182b24c9b9f0246f9e80d56ccd54e1b770be09ebf1845bde964906d8128d7c4daaffd3d9ac7ab49bc512f58c8ed1840e50c4ab6c7b1d74b902ad41d02d63d8fdd14b5977c33005360e0d0a14646879c659917d1903d448c6f689fcc910879477e35ea5f94f6c03ee842ade31eec10d8154a114de1583f74b75853907745a03de9c4341fa0c613cd7fbf3bfebb51c8380f6476a169ec47477c5c0a49479df1cb7912e0bbb20a98c5f346143b3ddb9f3653db65a0ca9231b9f53d5efeede8088d589c950847196cf3ddc7a96b1ebfd18dd95ffcb3df613aeba74c47bd5570d2c34ec35ba01f8fad38dbd464e610420b828672b013df79010d6b5e5a204570b16c484926e2a92b9c1050d9725c74055750680e019f90a472be91b76cb0e55f960654d9fcf68160923707c4a8374dcf055dacb0839fe3c7d19fb609a1fd55ffb497ee9e990934f2920a09c2328c4091a10d00bf023dd46b04d855565471521ebd79e4debc27c8940509d4dd5f88745;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9d5a33b843af55d5f3913409c815931577467a2e837750f6c775861ef2cbb46730fe4badc585e5cad7a13d1c84de2f048831c3cc8baf347540972778b201b0ee34750c9bcb5a80c4e37145c978d9f62a764f88676f786aa7b3b2711944c9b0f00f674c6e436f1d9f506430b711a1e08a3d18913252094f087f89745d00c75787c24ac61f5ce82cfd50717477a513fbe6afa58206ef5a897ffe43646dae4cf6c6acfb6f533fd7170fa19c5dcd7a739b95968035a3cc972dac414b54d32da4ef4ac8e0ae03aecb2a9236bd07360bc7c2b4464fd34474c1519ed79e1ecb259b03c11ee736ecf4bfb12b99f5713217279115958e17bcd6dd275de34a1af2a1e67de82d826cbc20419717ee9be0f31bfe942e0cd46eb261341bec8cc8218fe6714c03bbaf825e12c2ad55490c5018901d77d7bab9a18397949ae4ddad577efc8defe48d8150efdc950e032bad1a7238d876bdc2162761e1237dabfbaa39776d60163486e07f73897e2c4b239999b2d9923cfab900937e13d9384dc76de806f4831d4840deaf17902c526db3821d699aee780daefaeb251a6305704b1811c80e7f7f92c38145f29e5027de2500b81e1c697db79dc71f5d365a4051daeb39e7ee670104b765e54ede103ee9bcbc4db9081b8f3daf3363b20b6c57b01e12ebf29f4f3607ce44b6bcf569b3a42f9e1b82c115bb9d0b28d48775a11e7a780183a9c32d19e1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c6e92122e6e39796e964feccf5eb1795e71ee5afb17b4dd0c52b7fb808c615f08921374159bc133ff786bfea64dba45388190332537468917d123f0a1327afcbe96fe6cc5535556a4082d4f20a242f3b30c55013c29de1714cb59e5ec5cc287e435444d280c36ebf7a7f6657a04ec984211fd29c6b18e0f023c50353deb7ee90621f1552c7fbd7c823e061c47ef673742f5aaff2144ed790969a46555a650cffdac64d5a9c0b3eca46a383a69fcfbeaaa9a57894953820c5603ec825bca7f4fc7c532895764905e0adc07846640eb634a15e3993f21ed14b814e9bfa28de99cc31e3b1a2374bc4b153263f2742576aeb1bf34744ad967d5962fbc015b0d7e62a14e3c73d23b7d4bda1545449d0b705b4fdbf817b3d1a5791c147025ba0ec7ebdd078df3aded2cb4b56c94a302a14b7957d74e1d0f907633c8aaf1a33fd650872224216f33eb6aa7a808ecc3b341cc9017ce27698d46d2ea61ce066063128ddfe78a3b650639b928b6a84fdfaba93dfaa7e7ddbbd347dbb168812cec09111a8125b30e2f091cfaa09662795d3362273714edb37360d203c2ee77f069837fd9c938bf2fccff81f385dbe19aba029505da2407e2e699434bcc8bdd58b05e5ee87757e360123bc6413a3678561109853453f9104f4b9c6ab56bdb6628a869bbe1eb307a7b8b0b21e559e185c22fce6979286e0283b370a14aae95b757798167bccc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h68bf3c7942e045ba74682b11361ead0a6e47c53186e15de327a20d6ede6efe854d9b2a989eee319e789798012fa36dad93ae651312d9336b78f842a506952a6f6b3f3327b9f9cdc15e189d620bb5041ea473e461790f9aca8bd1a2f1e9f51e0e98e9f7edc8ae16bd79a00a6c0c70416e224d76259eac56b51aaba7d76ef448211c818cb880b08af555d9c271f7c4bfb1815e91e823aebefa7bc7becec944abc133bbc6384f23b6e6b0ff0813ae39f161a9c6c34617ed839ed67e8d34a1aa2e01e7106611d00f2ff6c996ffcd7a6aaa1d9305d88ae34da25f2a775c422f223aab077cb5c2db71e9c8e40a9365c0ab59da032f4fd641aa8e73a21fc262aca3be416c4e2a6c0abf86f83460865c8d83c36fedc6a9103e4426365937e47f64d65f529d2fea926828da486d99db117c0638b0718005e7afba8b36a12cac1c85a6305a35d75295e34517c53e6af1c6ab036a29a89304a163cc6488ad7e79c71eda7761af9e079baddec5a84e3c0f2bf20d6d08750fb177e2fd8b73e2ca5e400fa41a7b54669c7843a06b88206cf1d46a23cea9fe95f62bab03a44317b71482e599838e6a1f9144b17aa923e08cd4494dbeb2b607e832a3c019ac3962dc7860f61c166b0802f9f7d636d3837b3138da524ca49491ef6c6e980fb02439df8cfcb8c50e052058e83451afa18c179fa33385662cef958a8a0598a25aeb108de2ef4944d0fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha65820dc7d9fe459229cbf63f68f95062b6e212ae27a50228b4b5be1d110f496e1b2eaa2b818956fb47fc32e29145fdd08500cbc2dce202bd3f79d846d3d46436fbb22083d1352a50b791f66ada35c7f9198a273f44727f139cc16339ec3811676df51f7a312a336b32e4bd638a46834185431885592a4f9d3e03d0155ec881e9c4232105baefc28479baf251ffa71492a3991ed9963c5bdf3aaad962b318a161cc8cab70ef0a09372783ed9b749acd9449eb829e53655223897c676ad791563d54f02c08c36e5b872cb99cc52871ba40e3d249c8a5e730efe0c32921811f5d3e9e24b151b87c56cd552e2013a70fd9a65031311d96eaad046374e59359ca61e0761b597b81f8ef8046cd057cbe4be847e0aaf992278ed67b576fd5d5370cf7ae7ac5e5b22a12ed50238426b64c85002f7aec9c4e732209216e8e5eb2d41feacbab079a1005c74385b919815b1f2b76617a7369a2c2f13e940d831acd53f3424a735711d9d84456134dc869250d79fe3655e21cf040052a11f646f5b27c5c43313492abce4c3f55c69bd647374c0aee804ce5990b2db3971d84295762cca5a4abdcb4b96cf7cc7c0c5a8aa91f755eca2e29eb48d0474adab9e49ac08b2ec3dc035ccbe71803c2292603f55a9e86f164111aeaba5e73b939895f6c3d690c9057bba14b3be12b61b91f35ce31267f1396ff95609ed40031b4f4f9c455d8fd5d16b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5b36309ce422b019d428995408691ecd070fe43ad7ee199340d2274116b6e2b689c94b49d826605d673a97c08d96f5f99c965bacd9deeb23d901167df10e68b770941da6484704084bd53e697d37cdc73956d9b3806d7e744f860871ab098ab65438f10ea27f590ae0681dbbb9a27a83f22b9cba051dd2d68452a22c9d7948aa144b15f72e69c5215a18c2dcd631b269dbbd67d811ebd96f928785eb53411b12fd7b2200bcf701f47e6d46adaf5f78a01f10c7eae4b221e7dd251f6a5b1139a0701d6a9b0a43af99e354a5a5af814232d6b9079512cc789fca2754a9e7bb7a905ce46fc39da14a52854ea8093b9e5a9c3850c3a3aba95c50430d6ac90e9967faf7e3129c5de711f08d7b4aa08bd75b3c2ebc7ea85c4f68873da8a6cd80b456b97af899a1f583403bfb674500c5d2b536b74e04ef238fd755ce144ef192783b60ad2dffca4431796d2cbb98b0ed03cfc2f25a4fcc3b2965267ed0218740a20dde207289f86282ebcda10cd8ecf2728b81e5be77fffcdf825ec65e1634348ad9a3789c4378454af6e3b887ec0ccecb96869291fde2f0d543f7754699b5aa06dce7ef85bda960c1ac9f55ce9d864ffb47f5c6f02bb10e4611e33fc339cac99769d844451fc0960741ad1ab935d5d914ceef8c67cfbfca0d133c1f425b194be81d338e5bdcebff633e6d57e423e8dbe590e70b2311c0bcd6c9bdaaff199f9deb525f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h641435834d4a7b36befe47b048a899de05ee2d78cc48347f9da68362ba20bf1a86d8dbd0ad7ca0284e450dbefbdec3420185899022c58bd69124a99f6244a86fd74e0756d1373d52f9ed0c39d7208135a4afa689de004209a86e64ce2e480aaee42ab5b32a2a674b000dbe459d699faa5bc9489a257b49bd754075e00bf891104d10372d330c98ff7f56d82408aa1328b75076058ae10af85c805455c682c27eac70b58e63a7827bd78729fd75d375380ba1e040a8338e0afec0b3a27fae2723bd19607e8db2663c215048c20fda4e821fa56b403b20e163ff86022ee80ee7b68f876e4d0160cd7acbe8bde60af12a844c053f21ff08a9a1fe5baf384a267adaa5a41d28e9c9397be323723a365aa7a9029ce4606a0114ce8d1d09de5c6782de3f97b8e618710f290a7e88788267d7d32b3ba222b24bf71ff114593cd9b35bfeeea659fa1dee4fc285abd44e5fdd82c7bbdddd822107d502499a5222076b768045626c6998f1d64d3d87dcdba8675f474ead1256383e8ca89f1cbc273a1c2382a8f522135d1a6c23d4bfe68447110fc3057dad8ea024c7351c1591ca740c2a0601f83f10d3e52f1204bbfbc62a884ff2f75c512953b7a28d0b045ac22b7b6ef6f8b7cd7047a2219830c5fd7fb5aee07833e834b9341bba26c4c78750a116db7a7c369c6fb880f9b8d98bba043f3893c4a7cad1744105debb2cf01462615d8151;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h563a69101ad7e9ee98baff55b480fda1961485430036b2ad93d4d005064024815852e4fcca0545b0aaea2f11582fed4eb0b0bd2d61a8cd3fa2a982178975cf930f1a06c5b05b20355d66e6b7a0a5c1ebaabc98fdd9e405b92598a6b43421669066fa10eb1c217bc5140133bdb0da4d87b757e78c92b648491788c602e0fd01a44e9046c0a028fab83349fd30dc1cc409b98b9197e4a738ba42a7bbb795f0cfe2d2e8aa8870d3ce9baf87771b23a12b438b955baaa8fb901248d3723d574b42703f318b3150ea70c5395c085f5f13369c0704480fe73ee3a27a6a2140fb06cf873759e8d473b256ceeea2729b38c1db65fee35effd1c1ddfd20a3138f19f77296a23948e4024561cc2071888d285e10bb56fcd8f30dbd4a017da3392afe919681b5987865e171c99cefa9b299822fa71adcc5f950139e616410c34a9e8ecaa772762825407f07961b7230906fb515a7c456825588dc68dc6e26cc56e1e3342351103fcb4eb1d2cd8d28b42705f5dc879b4836feb432f5ab1dbf31313876152eb18ee277218433b6e1e2fbe552717f2d56b85a5c0f0a1cbb67d37254a1632dc457b19a04853d9bc1093be9e8e57000dd3fcdea900d0371a1be009ddc2473c58ffcfadf2617a1d5d1ee457bd18695cb347688d17290cf7c86e11a45e7fdf08fd02ccca0819a6475a57d1b6d4ef8982eebcabcfb45bb1b9f9db741b88e3187520998;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb634651a7f4db50608a8dea15bf9db1a72580896fa3c2e5b61a13485a9672b655a187234cb0cd59bc10f86d6e9c535cf3fe9331d09b9b33e2e9c84d02068cf234278918687dc472fc00394c35649723805e23cdb9bf6ca116a8c67428261b90a402870e146a3ab5e4b66b6ddceaa79a741d70e12aeec48a827997bb3b724ad90b1d915e37877e8db5474aa908b10123861ae489ff570dc7eda71b87d84425570dd14c28ea9c661afc932d0d70bde5a09066bf74531151b65c0158fb6dff5252d2d30d773ba382c033e6bd8daa01772da303750d90df455d1d5cd6e63c1b035c18a77746e82e4b509c2ad8546f6919785722209b6758d67f134e78bedb31149c108f77ec0a73479a225f2e2d185203a3d1b356f035783db0820c7a91c96f37b97b15137832346e86526a78acbf8908495d119f76166d53c48def51096985b27448f78c5bf162105780a2f6e31766819bef5ca659460acc10ea24a7a7ed16b0a4005b7ed52d4fe2ed0887471245c4b2a894e7f835c1f31344571dd0a1b36cb0309d6d3343016b9c7032a6679f09b7939f9b938240110b06bd3cd6dabdc2e4de891d36406f1d5683c60135c9ff2fa29920903f80208c2018608b9d40536e5c5268f49f9f891aca7876f85838ef2df4f92bd2ea17f5cf654947564e0dfcf694086a43d07004376e431ea2fd8f065636b84c4ec5a7bf2fa521a13d17ff180979fb2a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c5bdaba508df20b5f48dd6d2e0a26a97086b171c64941b886fea881c3ff09f1329cc357984e800a5c9bc8cf57129d68f20a406538d0467d6872e820da41a59e88838e74fd5653bf2c4a2ca2263ca4b6c49c24029824fbc6d4696e3dcf4b7ad77118187e3e389bcb9f432e8caf5fc3474783d12f0fcc1511d1c7a3356c0c4269f4d9dc7c9283665e880d089f3575ec37e6ecf6ae2ec6c58e826ee0f9d1f6e56c551855e2ba612031ae4163d6fcbece17254cc026e71969a8788845cc674d25a96bde9553a5ae1b823e3d6d8abdf080a05c327c70cfca7e9bb21fd8d6b368956710b16209f996eb0a4ab4c66d33e8bb5806c678eb63dbfab2d982287976917097cf45c180df9566422b2f398b1cdbb7346602c8fab693e1ad2e24eb57156ef573ccccabeae65783adb3742d760691c12ef7ebe51ea08ee401023b16da926300e3d6ee4faef08ad760e20ca8b32e790cd5ac822ba7039216c22fc71150399326d96722bf05e8f0dd38f6a74178625c8225f65d695382cfea0ebb9ad09c8ceb38670f685ab53503e549f3f7a0cf33354de7c2ed3dbd5c0eb6bfee5f0d3dfbff782b6b20e57947b6919310b7b38c14207f981a8e176d6c137896157619f565fa10b4c16ab512ce1bda47b69b4a2230b22d94b12f06b7b3fb30843edb9a9deced0b4c648c979d73c81c366541872dc72dd31892a25e72ba579194fc5987506331139a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h56f28f417e3dd86131462932ef3ff3150eae1f460501e7fe91ed05c45b484e54dc0d291d7ce791badd303677d4df1d980157ef3237949eab6eeeacec3dc8049e9c03c38543468f888d0a38ded63c778c0540610349ea16120ef2328f081d36dffeccaacca1ab9a7b0cb9a85d2a1204adf195467602b6fef772c6e3959e0d331d586383ae5e38eeabe8515ace5e950286b48c6e62f181d0a1df66c39c7dd831c94f6fe92ae40ea1d4759f3a9af23a3aedf0584675b2cc4658444d1d4880bb3f9303ac77ebd97724dc05ca1b7fb44655cc013d1091bec444e194449329a8b3690a02907e107bd65fa809c9934a93f96011631e8796addc651505f5e697d1d43cf602581c2fb677a2270532ec3b7e14031306c88d04ac03c70683f3cf386d5d2d5b7ca4144b8233137042c18ad5e811192d51aede6b568fb89e472de267c81493b074752d7aa74bd3cbeb6fde5e9759e812733eb07181cad4cadc357199134d8332c5e17dee71f1652af1ffe87e011a3af286e487b8e6ef69c87c351c368cf5edff5261198c367340b099d57b018bbc5f13c482669c2d1b39d1cb6e12531185b4a41e330e26532146b23e524be4dd8a71e79adadbb61cc52b0161cbbb989cba9943f61a86d0e875904b3302d635e55c7143f20e1f55d8d25b57fea29a827e24fdb6247f4f0e167cd78de4e461a365e7a26ad28c24b9121a5577be5472ff8ff0afa6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e6391f13cae8cf7ac02e5847095a23f13ee1f74079d2f015f51cf376c2d34a3a7b569a54dbd3f9bf41e971fb44620eeb4b7ec5d778a9c6873edb2b0180ae1cea7c87d4e306a8047de3d1342368adf84d6a9cb3361126ef8e26fd7af5d970ba0f50d817ef5f9e1fdf888a1c2113d6468ed2c0e5cf7b6420eec0a4a184740ac81c13f29abde442de433a84383685e8a52f830e2c922f526de71cf95308fcf3a8108264e2b8b7cf8b1fbc4404fe5b04c34da7f1628701fd65018a425702c850f5f85c338627cd400efd09b159fbb7a1bc4f6bc60e461c38866fbded3a5113e5bd3e49295b3a09b7362edfff5655fca80b96484384b8ae82ae756d72b0e8df833eeb575a1f58ac686ddb4e203fd09068290d55a9fc739a84747392f632b0152faa3ad1cdd7992f46ea6628685a8e68b4197be34acee57bc5222e0eb457765ca48aa4e2882bdf5b0da31ee9a0464759d94706f2286f2cf5a83653b77eec5f7d487ff57b46826e046d9d3fb00bf48c25570b0c70ec67770d1a942601bc8aece76727ececc25389ceb4e1c586657956b108c85bd21381bc98ddcc72ec976ce511f76140cc2aa11176b41e47788fe71d3d3fb269c039a4b315e647617207fa271e9782a85759e98afa415614339d0e2838655db5dbaa4a905becc669c9d41048fa48769044239b2f18fdb7897d52ba654540c62001a9df63af469cec3d03a6b0a9b47af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he800fd6d990fa8f46b8b66d04dd59cc8fe287bd076a53e89910a39593a669011d29ab658d7a8acc6b3ff34c25ee23063674a0c06a18b26038c1668b566f404c4920fb91a20ea10f4e1dc241ffdea8c35d0fc5078d18718ea827358a141f90c71ee265d45af8b4cc0e068720b6c1719aa37480e5292afbca584398641118f2d933a7d2d65fd172ba27b5d6e92c291f6372039f52bd2c272be174ff2834c5dd2a58ef148d2c1550e3037bf3cb67d3df0f86b84a7de5b104ab9bb4fb3903de2b0297efe9f77c8efd2265c3fe9ad541b18fcad3c6627b646d133e1edc9212e6c0acaa4864a7cf015e5c95cc8355948a996ae0094574f852241892e0c3f93307b83ca2859fd61c9da561e3e9d5040908787b2573ce81f7e18d62366052c6afc1cbc7ca4b36a180b82380c6e5c123e6263a0b7c2bba58e906c721d0980cb5c2f9bf2f49460f2e144f2601d935b5ba1dababff747539e0a3f30862bbde47a1a2d291350d1d911b77be5f5f7e7ef1773d7d97fa671eb57d7013090354eeb475384d125594f6a713aba16d9c4b50181ae3dd7ca37729800e070dfa60a853e97e5c2dabc8ab088b15b8c8efa78b058a17b1961f8a24d770a5767df9b3317d3560b316335bc50cf4f0af02fd9d3e01822dba05db301ad4a37b343731eb8c494b0aeb4f7d68e2ab063357b9581b2516818110dc0383bdafa63cf9a41914381b759819d8aa952;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf37d04d3f5ccc236da91fa6ee5fe32a6df38ec83a4784f8e6cbc646b6ebca44c22b78c397a8f587d87e07db12df2af9af4c8dd785b72fe3db72807f5f1da095b87bc53c98aec31f714fed4e288a1d2cc248714d950a593457c4097593156a7208d6c91c29b99733b0e788642ed3ab72a519728c04869f7a7f078cb9d92b924426c542cb64807f3a41502d1c78f837f9d322f01c0d94282f4b8f643b7f418515de792c806b13ee0fa5a0635b3e4a0e381d82e4c33a0bb18bba1ef027db2f9992641c8a1c572472fad9d6e0dddfac6e412845f3b0ee1973adecb1d8993fa194d988cc7c0fe50ed6932f7cebbf5340d3deafabdedc3b0b291fc26aec163ac2a84127175c604340f93fe036016f3e82dea9b97250463192ae6cd309bb6149b7511fa69bcdd057c23077f5d499043d6f8e9297581c348ddcf4223f78d90e8ed98ee4047b8a026322d9cd78f2215da77806f3946fc6668c965c7822b660994e0f425740763d36fb3b5254d3605379731f979de0bc7319bfa3445d29efc2013606adeda0b1e4794db1a45bc947536c717cc43fdcd10bf7eff0217b157773755432f5ffa9f333b6b246c42190423c2f8dbdaf58a47cc14f697b9a22be49396b449cf2ca13dadb40a8e696cb784f8db273de8145ddfe1860b9943719bb316f755a87be0495d100ff043167db3e8a2e3ef7d8bc8446e3fbbb29128b981b932c674f9aee936;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf8cd6bc97f3ff7a4a7a26ccb9e5fff1a150054a9639ed974d3db171510c1a624bf349a20c5cefa2c32b90f6fbe20e6d540c618a87883c16a8719d8a3654a30dfae1275af407339c3e3dfc67dbacc79f7bb4ce2ce1a841f6d38bd14c52eda72ca7e05e397745086ad3870c07e00f87a0594ad45fa09c21c3da4a96cd4c63498badd0997d5af1f1ef860a40884a1425297fd10f5e10c4be2af2df0f62093c72cec840a0c1dc5cf55835472320872b0920d6f757e1ec85b4b3d7b749b32a12606945e67fe5a6c63a4fc3e03eb91a6b5760b303e0a0628dce6a68eac731b8768536016218047361b3566046710e8be42a3a2975465286ba4db1fdd8fc07176053164df3a4297bc4908b1db2891f8ad9cc92e16b0d29746343ad28b4aac15a31404993d5d5b54caf4647bc880194c6825d6c5c6214a9a68f511b92f0e23075b11f213723c1a32fc6afa31766d10211ccc87851bda8c4edc6211fb271e61c4f186e9281caf07b8cb30e829ff6a06a69234ce8682a826e66300656a7a99086d40d4145fea9da6bd2719ae38d2bdbe78a28dafd80965bdf7a083793e52ebc8f4a29b90f496ef963d611cd65c5fadeb713fe35618b68957e1eb487092e5910ddfeb236d14dbcce51945a3f8841db4d3b692bfcb996beaad658f7400314e79df7573d9313f4d99a169afc6f0b391e1cd5d379d71c367cf287a3fe7fe1f4892f23982c2e9f1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'haff0c6cf3dcf314d15c4bc47860b080434b54d0cd6843d06c0e5a8303eb58ff8949ef6c579c1a4b89156dfee59b4777146577ff9cf6021e3dff41ab3a50098c3480bcf82b6ae436d33573b966d95df28bac809a287f695ea15a4aa81ae8f96427423a5e28c65e5a437d1d322d3cb1b5c593f09c276f312c933e4c052a33964c6d2cbae21d8b662e9b7f47dbecc05e964fbef1a2a1daf0886f865ae49ce22e85739f4e6e95c69cf689e50cd5bfe76b4e7dc26111ce68941482c687120c490fe8b3e9e738c62dc56d14fbdc9e7da9bca173e320cd135b42a1bcbe9b404ede5ba68aa7a843e5f63bd2322dd11169c16766492f5e839f5e23e8406a6bd6974edc0eda805be26217e371a08c37ab2f700bda732cdfe89c3f3cac9dbf1bc0813b96da0188669397003b00532f99c938c0abf70849f0896433c47973151b93343f31aaef67b9b4590ba7299501f177bacf12d1097a90b228dc814957a1699740c209052aa1f9640fb03173c40ce967958bf01133b4195148f8ee4a19b841599c7bd2f61b77922fa7e8880230fe70f878ccb6356b9ecfcedc2ece69d007bbc57b0fd5bc52d5caf5c48ac53ddaf72b4eedde1ced9adcb0f3429943f646e7613fb2a88abb9885bfeb2b02ff75938cfea86bfdc929c2d8708f3168fe471106ad2f5e863be79c4602680831d8d71ba14c17053136ecc1cea0aa56eccc7f8e3a9916ff34570fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcf666b5a5bd7a72b0d42fe0fa4231e7857e6892463c8751b1fcd5931a7ec8354f22d773f0d0f6ae41b55b669bc7fd842e6560727492ab811d3bfc2418f5df0b5c4e430e138479361d299cc9e4bb218bc0e1e7fda4fad416a7defab5bb1b8f9e70c323a1fd5036f7c80ca469704711af45138651a409c00b4ac221c6d6a51f3d44acec553de285c3d55a6c7fe6cce7cd4136de7468e05784c6721c1482300f159db39914a786a2db0c583e76d29fc272a5c3b22ce3e36c6e9ab2a3f6ab2c015d6001aa0ef2ea7f85440fb1029edbf4819e45ba45f5102fdda9d85faa4dec80fbcf7ffd56dc53ec6a92bd31287a9038e7f45dd5198f9ef12b62d0ae063c1b08e4cb7b0278b166b4ccb7993dd182ec383e192071afbd07b7359a343cd4771b3441274af525ec4c02db37388175791e2a6f336d32cf9902e842fa99dc74ff81141c863afaaa14e6aaa4a34f34576c78a6a3123a75395f571d4631b71ed8e44b1bd9585dcca9bf8cd1553118b452d7d8ccdbd0cb028ad685c946928a08853a178ebbb1c4eb60678e04c407a38fad81edb9707fd90e41d92e3b5ce5eb77a4056a8dafecc9df0c355e705ffcfe92429f94bbb9d726f1af7d045b69de86c191d5826c2006159c656f978ecaf0406fb162b1c1101778be225fd204ee67e277e79e97adad123831f15599811aa0e19e3bd33d3876cea8bd66242d43643f912fd2eba4d2440;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h812b449fba2e080bf4875b828afc4422afdcd598cf12dff49e65d6f49d2ea0589bf4f231bf4453c2ef7e9d375f807e5e02d2d5387a686afeb6f0a425cfaf5f3408e359614481b64a284aac19160c1f9fd912f7deb93f6fd9b7b7ad2a9959617d2705ff2cb93a1c6ea96ffa4944e20cb8c79db22fc2bb0d819c7ca49308e6faff1baf48b9ba5408e7b23610fa98645e7d32f2b8ff9033b9fbfd55de23a6b30755f4f6782a51ac13c7a3b1b1fe93c266373ec6d6f5a9b15d7189ab140218b7bdaedf7b7d82c121248d7b55e5de07f346b4e4598caa5c8e85044b195251880fbcab4673dc2e936f1d0bdcb110b9237023e32efa5904459ef161d1ab1859021ec52bf2fda2eaca518e5a4a091ed86e4d79178b5d8c5142a1cb087ec0b9b86ef3f264c61b85bb60e65b71eafff56503fe2d9f94316aef74fac6fde35f8fb05634110b6b98e3b373077630c30a0cdd64231b32f94e6352733ad197b615fbb4ce6504a617129ad8d08131ccfa787b9609b044791256f1de6edf9c7da0c4344f368aaf8a9b3fd0c8239a66807113a6b0bda508909853e04cb0ea161a44f151720579c4267024c201c4114538c3955f3813f9c4684f6378223c02bb347564e8fec40f43bd97ed4a232e841d5e63ab3c338bb2d9c5bbc23a939e90e0dc55dd463e7d18bad7bbf826b23646204659846661eafd88376805cdf98555ed53a31b3b2751cf8980;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1ce6c6fef5567749461182a5629c82b433571560cc414978ec058464a95081d86a3f2682490763e3471c40b16b79e7f2b9a7676f4b6c66c73e6ea1b2d8a56e442be39e013fea23056732c1136a2c73db9bf1ef5817a8b7e93aff7460c0e6b677d18856d6ba89f81d7fdd49b814a6727b435e72792bf34a0c1e686b58054e5dab0d5b14cb62400bbdaa44e23a5f38cc7c55abbe7db6adc4c7d8a93ff98248f2bd113f933d7b0abe05847fca6018d4ac7283a87b7aada2f10821648073a453491a78b9b6e6d7cbb8e731af0db82563e771f79f12e40ea6f023b7f2a35e7a60265e298020a1534e10b302264e68ce76bbaa593a2200ed2d55a1348c71e638edb0d0e5277b9cb4e30872c37dabb883d41043ca599efc47d90bde223e30a30dc378d419d73994fdf5813e99d9c5164151872b031089268c6db1bb7a8f0f39f00cbfe23265dccc72416222601d4d44b31de585c94fce14b1b722d823e3a0ca18c07029f67b4dc613df8fd808fd09d47a3349259be6ebcc50b308718f5c40be074f68c4841c7c9ffb75b57768337559d4dfe41d2a78724d04ff369e6a95e1994ab3800a266c966d551185c15a109c804a2bca13b07de864c8239842a96f3437a6ae3900b717c1d80bd0f875ec07509001716e7c98f4aed804b879d860dae19be3cb7d278ab5bcfe4e1b3af5c20b3a5c4ece512284c79dd60cd6d836fa5cee7aea934491;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he75f1b1aa03e2ed00ad60a147a3abd60639ed301b83c78844658bcd7c15da5b906012b29867708087b871049c56ac434d2f2d0d1fbc7d31f31d7bbd136a24555f2859cbe05e7a15f23c9c6bf2239036f4712efb6ce2988c1bbfc9c2dc725b5d59edaf34e7e5b9abfe6b3de654908a7f557478f94f42e1fa998fc839ab21a0ab8c4a9b567618cff5c1a50c797a63de928b1c1fc8d7a1bc896f13a16cd7713139d47b4c42e4bb7ec5645f909dabd0b8995dccb2d19d1f0ca7bc6c1a0f56cae22e8476b46a7ebcc8581b059c60f22c90d6dad0fde7bd80e20168876bb5b15ab28760165095d2d742303ff497cdd60b71c153eb791a7b73fa412e719db71f83c5610d34b82be36ff60384ae737bafa05effee8f36ecc43a940b262a710e8edfbf33f36874fc5f4e2a6528fafca3e32cf92bd7be88f047243a1d4a725178845f16a73e923fb9b626c46963e5af7a45056ca7d14c0120f88fffe35ad634be04538e9c891e71b56b89ea45fbf97f6108b1266fd64fdc63124086d7432a8ceb334357ec42c028ac77bf7a68f2478870ff27208e53e7aa708904b0e286054928560dd8bc027a829b16b3c3fe75e9eeefd81ed434635d525965190b3b0570163cf8378185fc2469ddb19f2a84c4204e920389eddec3b8df05fff67754d69a40c70769bb1266db85d6e9c17635873a1b94e1e04fff195bb86b2dc92da115786fa16f5e6dbbb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h79c955a85fba3fa3aed6d4392d3fc72ff421f60ee492bc76ea870c458f4d80d723e5e47704d450f943a107b7537e6aef918144e7808f0d84bf82c1816e288dbabb6a2e3f1c0f967d3d5c1668d04aaf366d859f418b8ef58f8d9c04617f5719293c29b11258cdbfb6f4f1e438514c3b67c04e5452cd951008bb3e9043ce144e4fe247006a811e0e47ed416fe0e360666999232cdbc6ea86e8885a6d3d46f1e2ca3f5edb4471e7d37f1bb3e957d2e7d429ebdf5879063671655b56cd36515a6afa09638be67f9217760d813a1dc4860426958e0e6faa42300cfa522155b2dbd0b2683b2a9c340966a4326ad30056694c106097743972efc5ecb54b72e56fd03657422b76b3ff608bf403eddc4202a2da0a810ac7dfc509efb8dee9c648e4f22a257686b2e8df2abe1625d86886792251a177dba53924d19fb7eba1dd0111661bb535739d2c80930c64d4e7dcbe41e6d3d67cdd298a7965939b5dfc903d30643428653639e1f5a4d47a6810bc808da02140f3458c870e2dbf0ee7b42f57b303b20b3f46a7b3a038b40a8be0fc36d777f3e3dd7acb5a7b4fee3981484a56cfdb5d10cf6427a99fa35766cedaeefb01009852cc1d8ae49622579d492ec6dc522abab4e721b8a2710cd8d40d5babd4a3c5c94fc4da07adb8adc6f9ae12ec6193ef3d7992b4974266949bb26fe5e59dfac5839e04855fff10e66cf7e25d206b84de8fb7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7ce4d97bbd06986d5b9bf421e96752a4aaa7eb97f101d11b0542dcf55e58571f1fdfbd6078aac00a47c9bf5c34b4f0a523878eca49e106fdc60c303a6bea812473d138b80bdf611eddc420cc222e9558811745135158ceb57fffebcff3bda3a646b6c210916fb94cbee6fa4dd9f78ce05c904adddc79c279ef4b373ee3a0aef9af687f33cb16342c8ca63d62c0fdfc4935d0e2a71d24d162f8fd1e7142897cf69737ea268a16ef8a6440b60b8575605b5f806e5d8399265c3df19da2493134e7b98be8c70156b80ea4baa468b4cb10b78909c322cd389bd6f4e5e7e032059ee82325d097fe7696055a6e446dbdc2c2c58917a614e2b94e115be215c4e985b88d617ba8ffbc32a680365a24c6d35b268f598334da782249cab4d6a519cbf4d9d63fd07e7f2f0b9f1fa326603719cbf84bb039470f757f0d1067b37013d1ae385d35d4f342e2ce7347200ab7e1f03dcdec5ea5783c6a0011f05145d3b8d28b0f3ae4c53c0168ce7adbd25af620f5e0154880debe0eff77acb0e5f3b6745de053f7051d7486f3dc0758db2a133df4516eece0a732d3e6d5a6d644cfc1bb034b2229b92cd1dcc43eb44be862ec4b0950919f420e2c77efcb487bb7ed092dc2ecad976ba50866813fd22c9e1cede021d2cfd1d13e5c2f04e51314248ba39a3a6140e51d2265cfa0fb74cbf0ebab28597608ae92007759196c571c530615c98d6e5613;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h31d9f55fecd9e47f00edf962e88beacfcc59ff9ed78a113cac738f93b7b149715cfdf849d99977f3518d7d94a59aa0ea573ac7586620a7a405b451c5bc29b373f9b7417be00d8e0146d0620ef56ed0040fb0eab5aca443fc901fa2ea9dcf5b888d4cc0d8ee464cab290498027f5eeba4013fa7b58b42b617ea13f5387169f2e8cfb6671544df78e2b6633e95c4b61cf4c83093b4803b00fd5ff58938c69ec293b872e8fa6e2d86fb2319af0e47ce743e5987ce9ed5f4f898f789c07174c0bfd367b6e7d6acc745477b4ade8f4732eef8c95745cbb702fe3005337e951e6f22b81b613425e04df42a176c720f19bce79afe8f6643ca2b954a2f5771a1fc55131d963629452a541317c0de446270beea519d3fb07d365af013ed6f7ea36d6f37882c220cce12342afac402322eeed9cbf7fe8ff9ca25ed5b1a9bed479d228b5e3dedaba4d7082bd1d4e5c03bf2d1fa2006b331fcdf378f28aa110dbe61b0b99d90cbc89133cc1ed98a6b4008522088d7e6c19f0be8ea715a720e98ffc43db28fbbe79c61f74c3058769c59c01d3c68bb6e4c1048cb953f8288291a99cdbb39dee962d629d4ff514fb55539a055c6e23567994b88da81aa59f514c31689fd322faa4a3588b7b8f9cda803fa5ad61fcb1050f4c1331d1d8a015ffda1460edade211150d8059163dd4a197ca72c5ab8a82763ec93e9e167046653b0c1d983f850dcb5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5ae7e10cc2309a0cd0504ee8287b4bb281b00a58b4c5f119297c85937fdabd757ae25275d66a69a2d887027eab8557cadf9ec250eb7f85a8536fd334101655d361f7075e7687ba5509418cee65dae93c21484ab0b35844e82536f53b2fd437c91fd72d9b49d7896c30518bfe372433cab130a1217226aacfc36e18c278f404bffd5b1f1be850f6f8f9b3b68bea688aef54ec2da58746cd7b2d5330ca8b2858a9670da2b7431b3262e7074f039d7b527414460ee2179a19d1e331979b537d4e940184e6d551a739ac6c49751d04f8d4117afcfd2aed7878707046730c86b7cbb11034ac6e013d403e1d025994e5e09b71724ff120ec85e903b0acd782dcaa9f65dd502958e34e0de6ad7eca7093470c29f0721d22f25eb096b79c2ed9ac0ee8a773cbdc03fc0919a8dcf2c5bdea24cad9eaf8e53e550f8aac26ccb58bc1838d90a5a546ad5649e2b1d4e970d598743bcdd37f46c30aca87f4a627d1ddbaffec9493ef521755bdebf19084200bbb733ad6533749b6a101ee09bad4df5a9f5bfe40c8fc575248aeb55912f7ac2283db50770fdf48318c73cc910b4106fe1ccdd937bc2d57be32123583841444ddd2d50dc991571c93562fd2be6b4806859ab9465411fff87cd87a3d733fd31cf2da2e28c809bcb93439a1027e2babf8a6aa71dd158492faee528f0fc6dbccdf5b5c833a5a8cfe093f79d69ee1f439c18800d70a37;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h84f44b443f7b5d529f6ac05a9b29d992d7bed57b0026cad91c14ebfb3175104e6d019dc94031526fe690fa756333ef8325de7773ee2bcf2a3a78626abf62148549957587a2fecede1250e486210a6704b30472d4596ca0ae8d075e63a0a521da74d8143d39878a2529508d4bf3383e374703cad40654feda0e322a9ac39cf5d869786b7b63209f210466dcc3eaae95540f2eb47aba7b5e24a5bd5ec521febf007396202c4d5025f15b78aa065d5aefac1e7bb6454e4d381427436f96fe0aaba24afab46f7ed7f13826cc85c9e8311ce84103e835203560c123a22e39f4c9613bef0e28fb2c29a697735ce7ad8fff77738a3b1cfe6d10a962d744ff62ea2bc9a2d3051884354e5877310a6e47b3c63dcb08ee1d4363c22b83e243a8cba73d61e80d2aac45a7b6b5f31cf04fac7525812a15ce1289f929884bc9a8f418d77ccbdae0ab05f131b7d8c8c05cc7d01481a52cf6946cfabb4effaa7d743bc62048dcb62521f8bb688f07fc219b1d68b954aea61841f5c8738a818c4db14cdb5347cc7e5ce0c982956c9e50160aa4c7f72491ec3ed56e194ce042c83e5f6e2abfa5ded4cd4ce8e9875365e70d74016661e606cd8b724eb073452e7ee92803f3196cbe5da163bdd271879d0a0f1e8e6e9b5aa7cb1be2a0b49f77be25a0d17636a22852b808877f1ff5a83fedb9e01d98e09c79a65a55c969de726484c96ae03e872a6712;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h567311b9d8c6ec3b283cc58f41a5c0981edf293e28eb2cc70bea65dae63b2ab71037c1b813fed27c3e4d7943b1563a753e25cf9c62645b0a4745dbd0a323c76f8cc516925b60fe452ae44ea2e7808905844b64fe1f109dbfbf84bad656ee30645a1886cd9c640d673f7faeb4fd087abe60d1e7ee7c380aa7f182207db5f3d181a0c720844a65688677ab7baaeb86465d795e2d5b512e462e918029e8465e75b1b90003a2114af60670aaaa5b6011bc269aaf406f4cf038e1ec90b2416e09bb9b58fe3a856928f593e7f1847ebd21797fe6a05f4f6c8f1de5d090adeb7947c40f02b455ec19e959ac87bfcc921b7de4eb22e9e632c7aa729af31523f431b11ba2d514cb10a05131e96590532d5e2e4ea1a530d7a7c292f10be94709015af256ef500f1193a607f5771f02f926f9aca66e2e89a516907f9385966dffd979f11f5e37c31688eb507396d39cc114faa02c54249deebad3d6067a890679b12a649898f282a281e136c55b7cffac17d6bb9ecd511e53b430d5146ff60bbfe62946d8a3fc2d7562b88675b2894cfae504d7a548bab1d142001f66106be03e98c1cf9f18f8d441cf8ffa786de91d2ce531f4eec5a187996b0eeb27261d2000e11443d4e20510ec0ed0bfb7dfbaf72f576483b97c7289b07dc29523f4ef4ebd49950427d0af20b94dbea27d63224bdcb095470bd1709fbb01a200d63cb1014284ae451a4e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf0dc346ac2fdcc22cc05ccc836cffda5bb55a620f491784361c3816d6b2bcfe5b41f56f78c9aa3364903d8e8d8266065688bb901185dfb2c73929de60a5357bcd5b91d4e8d8c35552939376436c7f6e8704bb961458ba9cd10a4c374d30f5ceece3be699381389ef6eaa84e1f05423bae7d92b5df742f24b65979b07f9d0184d8ec7831d44bc08fa43b7f707e50060fb87126847d493da265c853600a07e9619ad9ec27273cfd7cff99a31b769d6e3ff1c9ff2468ba8fbf57f0b7cd2a70f60e5ac1878ee7f246413912bab59feb130e399ae59153f1b62793fd28b4dcaac28df05e123fc5a7ed28ee29691df422f64cdbcf917916754003958c5bf3fe3645d7740913493e8597b0a094b27d737441d06c3c9c0fccfeb76deb10ec376dbe709f0d3b2853651bfa1499ae56358b3ddf76d61cbb428ceeb9f986069d4f2f9f35bf7aa06df32c831feca3ed0e39a819aa710e15cde4cf836c22545ecc5230e8e213823bf4e6e713d8c07e416536777e34079fa2131e77a0cdc29e85704aa88ffb2f6aa279f3dc5b6170ce0cfbb908aeb9f2fccdaa085fa10af2c2c038db1514b82934f95e16d41914123e419c844ef9a5338ad44a0a8cff2206b26af8aff125ac521615a5b81a77a83e128f5cabc13aae55a407ad6ef8ff3240e2a13d373b531bc54278a257b9f35f9ac95208f01efbcca9a5ca351acf85e527101f0b6dd0af73597;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14d364cb02218f2ae9d0fa4143b0ffb617955b0d31f3b16db97c97b0e1b21f42f4af046fb600f02251e42ae70ac76e21062a52c39737f77733ddae66fe608b5c59ebf5981ad65a075100ebf8f84880ea89f218fa2e2bb3dafa6b7cc252ac54debe3e496d2f35dd3830b89f51c4fd57ecbb38a1375b2e98f2f9185a9fdc4be30cd852e0a148b121b5badb249a465f3fd69a36319d7ba05eac8214a0339bf46afc962682688f9cb5d9593da6575389ec2e70d0f79e3b70234b8ec3f0fa2ecfa3413bec62f54a0a92f73a16e24088650a01308928f905e537b2c947f8cc39756d1ea8251d3c0bdab1c831137a319c47b22b1ee05e83ec70a3d8daefb839f74bd002787ae8e8d63ca78fdefcace43e66f57a77704c937b319c961500ebe869f4a68bf4387bc41ce43ba56b3daa353073398e6e9cdd7c1503f2b27dd26f34dec318d6282d2ad388fa58c771c5be0c999582d34782b56e4989c805f9a01c35d25a09163fd8d42f809d43cb9b5aebe5a4f9ceeb2fadeb58dd744774c39a4b641d69da6c68f4f7d38adb321298b2c65b90686a5e09d78fcf860eaf6fe9ab887d36c6d0f1c35050dd5f2880fcbe5d15cefd415e8f67c512a69748194fd7cd467cd284e5e723fc12b116802cd62c2abf93083c18947cd8c8a53a8b5d417d849ea2e87119fa478b038830b92febd7240cb5cc26f3b72a953ef67bcde42e187cb8ea4a031787;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6efb14ce07ab91dc8996ebc68e9223ce7a7021f2991ab7b5e593a4809ccfa5e691cbed1fe04c537488baf2ce6291b45f0ea492c3d4e0ed53e2a36ee6d0a4866ab4a75d8c3f65d4e2da04fb4992e1be169b11d2b72ed3d5357f12ab6fa3098f0a40cfd52f3605ddea4a0f23fd630912417078d57a6372b3c6de04707c41e2412dfc7de610695510bde97fedfe5caa2a4909300ac8538264303fa95742a2a6cb0a86645db1805c890923ec812663ff31f9fe92a221246d12e8e8b9c4bd86dc026952b02c60f7f5fab9724dda8ad6ba50b2f0b2e889c361d569d37701c637d1a813dc8d07726ffb96c9e963fd688fa7b08f7e6eb20ab2354ca1b0d97ca2c25a48652e1a50a74db3d3a134fa2abcfac9505a50034abb3fdd482b5f4e2ce31282aa607f36f2a8e03037c7f5a9ba31b5aeb9431c8fba1a6bc4a78d3785a9d3d5dd05bcb06d85778a73ecade956f51f1777f789fabb4b1e548a6676a34bbb6bffe31aff37707df5c1eb1660992446244b4e7f0914c10e1f96c349c148c105deba95c2497a146ba2f997db5117a37cd70709b3f916ba0233790b409f3bf698ad5d485541d6e1601beed5f9c572e96bce24982fa78d655b6d1e32b0f6ff66cfdbd3a4477bde94e88f0b3b8313b96127a7b3e5b9ed5b1f56b9d5982d622e59855b6bcfce78d3f62c7fb7fa949122bdc2f8c3b36f3732cd4ba18f1c67543476027b22525e83;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb94cd7dc75a64267d3d1c2c199302f9d88056b6001b80f6c03d9a5c5c40db0cddcac335c6fbc13064e548d1c32b76e6ce9f191de228acf0784e3c536a3b5cc1595b9167b273d3aca63438ed35b2f43685b64e71ae6e0d6dd6a07473545869c4e23d0ba40ab3e612a16899faf34596f079409f1f6b67e99c25f8b0c881d8f99e6d54b1b79a22918f8555c090eb6ffca2710a846e283f81ab19081225df8c8208fd1caae5c895881d3e59d9bae58fdd13e2652bbbc17278963a65c1970b7186936ab4a3b88854e79166938cca516c38040eeb885f5db57f0b649b0e35e404e7d256058e319684af613991d2366af76691e7479a585aa565f162fb7525d162f72ca03e19387a7a7ac0bd352c874e52f37815b1e565a86199b40f8585dd31f67565e75e4df711f19364c53f64e02745ea2dd5a558675a3c812f775379b2ce2fa245333452b32d5970dc56cf7a8c7fb72324bceed8757226ee82cab2ede6f74523eae2eaef18cc1874532f6531697ef24f66f20d0d5b9a89eed628d08889fc1167adeacb2d7baa3710511fb7b11055ddf65db303b30ed097138e24729f14eaa6c3c5347ab51ee55d33375d7126c94cc28073857fe74c35a437ec9589d16a0f16362662178f5411e496d4ba17c3594e1bcaeae8211f9afa511e1cb51c4d238ad4559118601c1115619370fa62746286d629a1c10553cdbca80a5380d93c95177435814;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h78065d4648834bf2cf142b35b910f12e2fb3f0c2fa6fae5843675a571d2c4458f2256df68e4c11e4b1a752c89e9d5f5e9eee9a6e963f0fd7a68a65318a44e23176bae1c68bcfd7d13d1bb263fcb59d12870c0b30f08373f4c347c5f491c609237f5c7d8e31b27b1039949d1832e67223300e0ac5925af863fcd3aaced7be555a45e4cb4e4c48fad3760a04661080ccfd6f30ae69d6642c02d7ef05279aef76d86fb405e0b9e8816dd7c4448029024ee280cbb5025ce0859bddf0a143ec4c0dbaa6f7df873f32c9078e204b991033e4c225d798ae227308c2244cdc32e6dfe33e5686289d1b0efabfa1f26f2f43f31d292b803ae921002a3b17afad7a6c0a24269ad8076ada60ffc240aa2d792af0994dc26d2414f3925ef683ab1331f99ec3a2b45249ddb75df890a4358d1e8161f9a182485275a16246c524d534e451df7b3f2fd42961c7027718c17aa726e9bb3d2315164e6c7d63ced360c130d60f1009ed1cc798714ec44cad3b1e3ad0d7ba5b9bbd770b46f36402091b177e76750c0c50ce98d460cb2d8c7f86d69da3d9d3755794bf41702c49353bf672e1ad4beccee24648173d27676a451b38ba95028dfce9697e708f721f69a5344a01abf4eb581db593c9fb42213456b9d61bfcbe95c4782b7f181f316f37894a86b701ebd07f497091b828863c2a1895dcae5f6875a8f7d65e78b3a3e886ee248974e1e87beef9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3efefeaf294cec7ffb0807ea1613fd30cd6ef5008b8b7280e31e5863a19306b1c1d8fa8f9a30be4df57f799a5bc5d3668e186c6c787e7ccf9cb78977f5267ceb44c1eabc49f4a0ed0d0f7c0a8e44cb39407b3e4c8387352e8ab16b2e8d89591d8a76298f3d3fc33d34aa01a5fe13497f2b056fba1fdb61f4bbcfdbda01c4b20eb70eea9087d55dc44c55a9b10bbf091ee6cf8a19887fba06069cfef1d0e5ca2e6212d23f5f5d648dd357f9bed87192942bffdaa72a21e2cc60fa6ea022b8b9b52ac72bcaaf727d6da2f7d4ae416ea0114e6ab9fb24fe8831a5b4cd41f6feca94e95edb5b381e2d9d4f6f99be23de95d1494b31740dc75924ae02f11ff1562b4de111b4a57042c7fd711690c1d2d0b84a35f9cb5f2e1750fe43ddeb7d4969c6eaa95ac4b58de38e01b5eebe5cc84fc3646f3d670779a4cf9233bd3f21d73b22c3ea0c10c80cd0564e26b29f2b13611aadafa6b31be10969fb1b02abda340301ec7937b8521b14eb175c5a1f6e0ef64e014264407f1b4e191f2e76fd6cea4a7ef537685f8158bcc2f238f900d9efe3cb09dc7d41421990e051cb191a3f4e6272b6695f61bd401d3996ea83aeed994dec5a05975fe6ec7216bc5a16fe8f052585b052503e485529a4502e23a3fe71dd6c5c173a11a819d5b6093695de549a792d92c6830e77a81ea98ce5169be93a591c88fcf017110f32dae8dbfdb7e4fa269303;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd43bd55bc5c3e3e440486fe114e69cef185c4bdc34423120861fd661fdae732d5e7198e266e9f761ce2445ddeb9975a9e56d93512ec3285a3afe23e4eac698182943014a7fa231631912f0389f1951fe71ac81480157966139deb48a65b9428c18a294fc2434f96fa9456322c552e598d132e4d97f6b22507cab27636e65f41d631426226c44aa638cb8d12de42c0d2d9384c0948b1ffe7f374cbd20d5c8696266b41b7d8038305d4b1307a2a99c05e8575c64168ef4c42e49e9d476d16ea5d13438d55f81de3ed18098fb92a7ad31b2176d353de7ee66151d5b61b8b73581535ff0816c4e7f404ef0d4a112e2871bfb02be2faf63fa0d539ab71a0ac9839cf16d545cbdee21ef2040422e4db1f227f7168afb3851d875cb9e467e6467b8907f2b73e1ccbad631eb74e2a770795d6f645699054895e01e8f4128412659fc8826039832cff7963ac674025d66bc5806aa7ce2891da16fb6548fa88eec852239d0ee0431866c25c58caa1831f3a94273c65c2c1e9916b96a39108c13eb3f8d3b1b9b50e4d20faf07e8599a9a982f107a7567fbdbf53409d42ebed0c64aae1a7fa7bd7e663233370e3fa833b9c43b690697ddd62f7287467ca1d756cae977774f353d1b762038df614f95a507198e948a801fda38e50d67751c1570db4f358d772d4c7a1de1373e650bd924c86d5ab24b10bbb44ce45e12b67de9899f52ea3b39fc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h12f4ca44f64d5d69a5805ca80de88561a147860503da84d1260e5013a5ee1d25557b8d533657b06c7c3de82ee54a497f404e0a9a5b39b71f87a27017d0a76d639df163c4729ba4e9a5d70558dfac3fe086de9c8444117074347b8b2f5f80f9af6537ef38984cd772f992ef2b38b0b65b8c914ee5e44ec5906513e4c00d87a7cbbf5bb51e57f273983b2832bc83556b007f46a94704f5edc45ae1174d61f2a8b111c664b4a3102bdc128b017780e4da69efed61b54f68d6249178f79476ec61ff3186ada01c3ba12b869c670cbab9cb68c1af9bfdab44862fb6141ccd2b54ee111d82bef81d4e7e64101bed55515b4bcf1c48b110050403d7daffcbcf153729cf3e5fb116338b685721b10d62da4e61b514d5f97fe76707d36c3351910afa163ab249254e40e34254508a2559de13d9320265d2684be040325107b61a498c57deb8a38d911aa53c377d59b76cb0df86ba90381529af2153b59e9956b5933d83cbeb41df4ba478ca74ac6f4f77045545facfa97ef0e8493d35591b9089e94d10cda78a27862d3a31fe4e9872681f2e8315d571314e1bf3d401aaf916f54759e3f4c26c90598578200fa9668b734841eec31b2605b0f5218abe52738c8e4e73f6fbb9f594be3b2ecee366e84de0e85a5d87e17eb1cc0ad41f5de9f5ffd2ebf758a6c7e9d4986402abc794798f73d6431fd78aa45bbff5c0c5db653cc07ebd154648;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf319ec01d3f8f200a938d615665248fa8328ee595a23c4053e030869c710594a97a62dd1fa4e6dad8e3894e595f768e6b9d9e0824ef4545a5812f32bc82d624f3e29d5305a7700be597825eb6ce865eeb08ebdeca233e8e61427697a27c8db528ddd4b756883e3012a279be739e0396292223614c6602214d8e9fe8b7d5f90ddbb9ceffdf6e96118de177d88308db5ff6ee07c1cb0407a8c642335436b3259b525e1cb67c86738fea0b87dedef1bff1a74951303fa02fe0f9d27be84939aa8ef89ac57b7c76f92a569d088e37da3d3bf60d1e14d27776d5c8aee924b1669fa4c9ad0a9211bb82e708f7d46a15a995c98dfe740c4da96e77de48632223db3b924c0c8c9fb22bf523906f22648a4c109a362716c92e1f7826a49c047dfc0cbd66b67f91ca53446a38fcd16de00c5249e8fa7755c0c215ea721bf163a277901592b45b9909d597c89a2acea9f312f440b4d24b5a9b88486a486333ef057508e0d05c8fb98bc720a519412923cc3ce6e0e3ed13d3dfe97744f769427cd00da6496daeec28e0670ca38a1d125feb9fd233e97583c7314dce19e9ad2bef34d7370ce3bdf18f116575ba712f4d0fe7449c2b3e235a4cfe887f3dd17736cc33205e095d1fa7a8fdda93685f03e7a8ad36de021c95a72a230e4c233eaa3dde1c22185f0aafc2c5ad0c175f2f6787019bbd72e65b7726546a44d11d4dd36cc28d931e6b66;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha02a108a1975eaca98b68ec44dd22b70ca30678604fe086bc2087b532aab24be4234296b4e388797e268f6d0fd36be030634a99dc88429d4829b8ad014adf88b4c11f88e0d9bc8c0cf22303ed0ac8a1ef1e415d31e03ce2d25960ef9ee17c8f04e968a027dfc0722597508131fc4bb3991dd1e3aeae7227be23db4453caa3f1d63cf8a3d3e49380ca315b293eaa37ba982d11dfe832e368a5747ec7386d2d3d7176785c6c56b22ded8e42e32a88ab91223366e1105065c2636db8fc4e9d65cbbab499762cd6354a77b066da75e2a214797a1cada0514522d7b171536398792571e9df65b91c1b68b11982541457871aabcb0510e744fa3dc51b1d1354ad9f3c462cc8029fe2cad8ed27b4f066fed433c4865a359323d36af32a3b4066829de5006d8201895e5510dbe33260aee285b30ea568fbad0cddb600cc6fb081f80e7744083deeb173875c48a121a2bd4af72df5f84ad5af4743e989a36d23b2e4318e88cba7314433e03e61714a91026a61d5fdc5ab72b1b4400595db7f20b22a719ec65b0450930c630ba8971326179789859bccdf878e3bd70f2b1c120d5bd481311b71435a84f37b58bed64cfcd66c15bd7403523778d2e07221a244e411f9106bff859ce1533b098ca21f95c2bcf27c6e3b7563a111ec8f75273cb7e11daeba5a982b7b2de77e3ed74303cf5f4a5cda4c4eaa6a5e7340010ff7486656d4d316084;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3c0ff597e6e817080a9fa6dedf6ab74ef419bad0e3f8c91cbe335ff5cd887ec05f62418df2b07ec296fab579751a47712d13c661e68a4781dc998f865728b8d3219c2d980cbd5a47d5e456281c78f726944a92373b6027ec069083f4418f2ca5a16eb29979fe7fea19f2ef1771af138ceadf15c153aa85c8ca4c00fa281374a5eb309c89c11469e77bb1fa7f98ab6bb687948fe992948c863e1eec02f4deb7788490a629ce7b3bf487fb6776460c863f79871221b83ffd2c52d94491b088ed3887dc5da55cbff772dacaf055c6d8cba670e4bc5b10ec2977fd024990d7043a31b62b8a906bf5747815ee8039ad23c03d28138acca0748e9ea12c1c922b6e1b6a9626577018dbd1d8e3017eb4345fd52d165e07b14a2d380a73816cbf6ad5e10e99cd4a0772cb1982d23e1d3115cafeaee0ec92c43917b81622dddf3f5e8ec41f8ef837930512d9402690bba01aceb3fb39580ec44d7ece1139ece67201222fac5b9a6f48b0ecbf699422ee66a0b0d788bc3d23a8a60da8f25ddc959b68a0df9b1af09231c18de24500e6568e9bb87d95b19a2e71edc3b80f8c4f456bd4f3377177945abff65dc3d4a29a000881ac70b8d03d2cb2c9d67f6700c12c857ecd90e7e984b764f11f0305489c36678eff6af4c2a1d65fd65eb16bc24e78cb261fd0a7353ae260fc95783b4cfb3d21ffb3a7a83cc7adad1658b40fc00df2b814146eee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc07bd81c55da1919843a3a300e79f2cfaa1fd16345a617316cd8f53e3e785d33527ac14c5148c90b1e9ee513e30f2a87333af565ee2aed975c1ddeda81f9d197ba02eefe405f1e7bf00fc5111b095da591bd8bbea0c06009d29d835ab811c07266b334528432e0c9126b2ce54091f7c904d2611a62ca7121c19f4496a878642f6df6c912feb4408bd75be09ccd16ee462238fe0a9f3f39d95925a721f0ba42e8d51b609da3aa7109337fb332ed3cce084f5a3ee37be3db13734b3402bb32dac08520f1f6a59fa069c2f3e38d27cde886221cefdc587b1db08b034e24c147942f5ce26ad0d8a6378ce4f605195b40fdfbcedb25e33592a2bac030da2186e3c928c75857a9d6637019cbd7bfff0cb21e129a1ec5319b4fef4d924e7f3e2ead22309e7c80e026b0fc8b1b915b7523db40018d0f2457033dc2718c2735dc9f06767f44ed0e151faf003f865be81be13e3d6b5689ecb983ba3926d36da395688e182d7b66c86f9be352a028ab0a97c0e85cdee8ad724ac8bfc099c3194f0dc635c5b60ed3c39d35697eec630008568a1232a66aa8717931dd6e8112499b063ea877546790417b8a8473072f8d877c0279368c116246cee4b9e5cd34bdbf851d1e0c668e9e2cef20263b0b47bbc21cdc2a7099307be0bc61e753b8285c0a1e60a7e02a28e6b4fdcf4fffbff4a619a1e0ef61911957dd584a25449bf12e5b9fd0a93fc1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h135f9d6007415a605cdf8fabb005ccfcd984c853a12268483e12bbbad9b7b702992dae8c76c67ad1daf2bef9fe8b0a30e102dcef595a1a48026a0f26fc0da617f4c22f4a6cda99b1cc4d230ca8afa531570d40fa071503717ead2e9b06cc52e8834946902879eae23013aef5826cbfcfe85a896f74fd7029323eed99d054764f745027cf9d2fd5ca581c1b96d3c7f333507e033231035a5208d1e0df5d2d95a2c4d6beabfabb8a58f896934de862bab7016d1a06bc4e0255c1ebc38e3aff352412f7d8c2e1d82535464b75aeadd9027be735ffe85b46b77dd829633bba09637922736ba9625e2c870b56e436fdf238aca0052cb156c9fb77d501d399772a0c50e50af11fc7bc75a7f001e0c10a9927d6980faa7723f771986b3108b30e07c4d506f037f4b2b82408405aa07fac356935caa86b81428c36f85c92550e68ee02c0bdb83431537c53044ca8ab8f54be8005a0472eb9aab32599dbf6390efd64f690c448ee264f0fa7d04272b6d8f861b5883ea1db13cea33011d739dd0059670c63dadb4bfe026df14d39056c057ee26d605c244435600962a3b66b5eb4c4923038308cd785e32b38404a6316875f6204560665aa8bfb91ec46f3e60ecf7b2511ff99ebda786d405368b11264600cad5707248c3a0c97daa8a7c0fc8479ba57e6518ad2d84557a9dfc2274eab0a66c6ca51f0ffbb19beeb4a97b4dcd79ab11097f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2f6f31017b357ad96b833f89eaa3b5ae1cb0f1a7867a870e18f9ab4c6fd9e6e19ae77afb2aedddb26d9f84d4e566dd3f2b4c81990524db5f4e98a67d032f39d3c72da0707d199a77a0ddac19c377862503c14b30f2cc157d177f616b096d634d8261849a6bfe54e31199c528c7506ff684fc4c539c736fbe92c5d933b5bb3f077b3646fe8c3405d2dccd84587aa1292b99f17a1961a13f4e3a9bed1723f3cc5a20f33bd425abff1df54e3f52a8dba6c12edcc3299c9aa96ccd8c6ae945db4b711d9973d3dbebc75c51126d890d2236429a415d5172d39df737c42c21da84b2afb6ea03484e46af4d69acd549f7bb610822f5691c293e8e493e6edbaccc2a6d5e7a9575f0d950c8c765a9c8cd269514e4170c4eb9cbcb1daab3f9397e32217db4e9f7c8c9bd50e88a5db9c63a5140a206b283c934a66058f1cacb7cc63f31ea8a2eee4b3a63db0ab7efd2a832c9a533a10711b8789832551e7694e3cc975420f511707667ec1e149b507409aeb36c58944a2fca0a90a050d62e6563b3d427007ff9c8708bd3fe6fd50b23acedd618dbc1b050b489def27ef80206cb4730eec81913c2411851ce3e5fcbccefb5e1a9f3de1b5179eb88653105f0d55113f39f72c59e0246047c122b88c8310b99e2bf31b6d30d5d0c3bd5854014705e63139015007444ff73cd3e93ebc9d9d137d92a2b83fb9f8dd52a579d7978d4dbc80e72c358;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h19d313044264609df3cd9a6d34e93b43280c705ad0eaf40077dbc1de7ae7ad3a067e7c6297fbf7e3fbf1c6d215371781d721a3945e50a29d9803860e1801ce0457be65f229f735409e08ae8c1566ec95e139e066f0d23883b135ca01345b9812b003cb872928a47b17f7d3d4d5203fa9f911c6cf0275344328fc68bbb0c4fb83f1819e87b543868b2eb2987785a9eff9dc9a87e11af2a98a22c51b834386ea66025df01088ab11a03648ad2ae249855b3af8a7499501e92849cb9fd45e7e401c04e5f1047d761d62cc75155bfd156d3fff9bb6ffd2d64affc7e14791e12215bab2c494e42d5f5daac3ac177127c5d8239c35cba5e059105d7d7c38d8634aea58b932bb5cb2bd722f6fdef24077ac9f140aa760dd7601c299d9102356aa15187eeeb04a211626fa13a255f9ca2dc07a4dc886dffc5263c48dc5fcaa72b038c95fff12eaf4e4990a37ab03925ceeda63d4e12449f1c4e5b55855ca9288aa60bfba5b2c2f6b8260c38a6c99b7583e8011bd0fba9cd05783eb06770c01d1c583ea0f4f58865b84a543e610fb5d20ca3ced40a7d0dd0af1b99fb462ac25d8f85a1a6feec849f8c09a1f95b509f0e80ad12fe8ce5a5ab25727a85b85d23e00e213ef0bd5449da462811db4b8731d190ba7864fb82cc1f790abf9717831d0b8b2f40d6cbd41bff3f7b688a604983bd76cde5a7e683f55b7529dccd658d994f9c5f88558;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha4cce52a8d79e30af5b63b9be4784309529ab8b4c7e215af6cf41682deed2dd16c607983c4dc52b51839f63b52f275cffd828bac4df9a31eb5da9d5143c0f85c0c3ca2b2f3e619672046ab438641d786902334ba326a8f57a12d17dfe4c32f28ca4977ac203ea422d8f89603b969008ec0946520f5b6936e35e076d9e9ed80e68ffe3b69af1a755a47d466d82d949486a955fe800cf854ade2cd6b46876924f7f6c9ab2e21b961979afa056f1e6fa8eaa0fe01d28341903a2cfa998782f820458f1b491dac2a38b172bbda5503655222c84959d7ed32db39a4b87703de31ae3d3b059bf24b282b64c5f4d8e7487a55ce7e92034be373c7c9233861dced75ddf2d18cf4afd9bbfd1f1ac2434be1fda78cce6c43e176d224111b0ff03c0f32b4045b4eaac2ce91b00f2def8e518ff7ad5cec00f35a583ecbd585e6e9ae0c96deacdfb28088f5f2872c765c93d7a5e34b31a7a3a14939bd109287361bd0a49686c129e9a79202434b6b7ae9b4642f20b8926ea8b876ff127a5adb622b7fc0896fd1ba60f847e2cb85945803e845adc1b4f4cf697bf555b198648770b0b289375faa582538365743970801d0a53320955cf6ed64ed876328d0e11c85d23a03938551ea774931ace9b1f1dbc2b6ebdcd50811b5488060518f2f415a57157bb4efc746b0dfd1d906741f8f54365342054fa7b5ecdd113a7012d3665b4178f03ee2f1f6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heb6c07306777fbcb5c24e56fa8dff58595a81e0323923c39cf68da6f35eb7760e94da18e5b8c48cedfd77b465a3714fc184442ebe7e4a994cdc3bff0051c4ffd072dd134cf6cc72300207d4208353cc1d855b321bf33d1336040c953a81caf2ff454b92dcc8102d82dc849cf06e9f4283398feac839027a15468f590e0b36d0c94283f8afc6203483a87a4b4bd7d810a05be182968421b72c3a3468b56c348aeae9a7d3af4434d5aaad5d66a4787e0dd6961c01deb84b40a680d57245cccbcf0384542214add2f86c5eaa7e1b6d937070142367c8db8003cf5630d27b369fdcb01b673bf8fca006b0b41127c4e35ee91c575830c2cf96b6464bb9d29c24d2630d815bc9b62f186f47dceb54c943558133a2104502f757132e72894c0f62e688cab6e6ce800e8db1391a8e5c5d31b13b71944429a15dad18eb6c1e6f5167a9bf9b78610022674a47aee93e58fbdabf6dd9714c61909cd0dd958dc4d60c79a963108ab7a111e51a7733dfeeb799fca6bea840193f1289360f846c4aa6944427d0b0496229767c0b7f8449f73c03f9e18f0f141d7d835ad1b82ea53711e4c603ea1f148d53b80b1ed01e2da6a70c509691f4563eb3452d2fa1636cf25ea7557a5b828c399e5d96202ac917b8d97103f47cd88f598598fdd7948cf482187a1df9a5e6418f2a40276e8925a9f7395c6fba70ab3eb8050c46a064330e769afcda0a661;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha865b85c9195296ef6414962167fb7b9c8792980559933bba972777d462f5d18074c7a568fd3b9ecde8101d2bc3ab3f784ab5abad3de0104c7a576d2af0fea7b5d953934d184451737b9965711dd6e09b5779458edcddb29a8e2c26b96ca21f6af2cb8364d9b22aeb0eb89fcd174bad08db8a0ec6184c1204df2b0e56c941b72b8f21bff1b0b6d1b02c5a488468a8774820ad5520b583f22d128e6277d9b5a6a5324a7059d9607ff8acb729cff9951f8455a4310e1c1d69cb710776b9796ff0078b5f8e7ab6341f30a0cdd595164ab04bd3dbcc04a032a4d4a4acc39362ec9980ea3b2a8a1e5be84c7ed568cf40a721ced078512606fca704f0d85948cc417ab3b222c0852f2ed3557a783318778de763359215f8295cd184b36c2bedca78d6aa85d1404fa24a8e5051c0efa0e4705d9a1b11bf22d9df3a7313ab096fb9637494f1fa278981d7c95c275bc3210a01e41467276a3ccd534dda20cbfba227912ed82182033e46f8c3e98b4cdc735b49a4e2bb7bbf1e456d5baf114a36c3759d657a4fc7f21e72729ecd8b65f3923f0b5cc5f80d7ca0da82634c60fa0d3bd89bbf207877b041550b4cf6fde14c3554a27781d0fe5e41a2119079b328f958a6975be7b46ba77e90b9e4c3c46ba0e89a96c38fae2ff85d914982fdcac4600afca26bd28e9a8ce483353bcaf8ddf46d9bfe597ea1a1d61f0d30fefcc2a90151b545e5a;
        #1
        $finish();
    end
endmodule
